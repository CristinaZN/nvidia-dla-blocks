module NV_NVDLA_CSC_WL_dec( // @[:@3.2]
  input        reset, // @[:@5.4]
  input        io_nvdla_core_clk, // @[:@6.4]
  input        io_input_valid, // @[:@6.4]
  input        io_input_bits_mask_0, // @[:@6.4]
  input        io_input_bits_mask_1, // @[:@6.4]
  input        io_input_bits_mask_2, // @[:@6.4]
  input        io_input_bits_mask_3, // @[:@6.4]
  input        io_input_bits_mask_4, // @[:@6.4]
  input        io_input_bits_mask_5, // @[:@6.4]
  input        io_input_bits_mask_6, // @[:@6.4]
  input        io_input_bits_mask_7, // @[:@6.4]
  input        io_input_bits_mask_8, // @[:@6.4]
  input        io_input_bits_mask_9, // @[:@6.4]
  input        io_input_bits_mask_10, // @[:@6.4]
  input        io_input_bits_mask_11, // @[:@6.4]
  input        io_input_bits_mask_12, // @[:@6.4]
  input        io_input_bits_mask_13, // @[:@6.4]
  input        io_input_bits_mask_14, // @[:@6.4]
  input        io_input_bits_mask_15, // @[:@6.4]
  input        io_input_bits_mask_16, // @[:@6.4]
  input        io_input_bits_mask_17, // @[:@6.4]
  input        io_input_bits_mask_18, // @[:@6.4]
  input        io_input_bits_mask_19, // @[:@6.4]
  input        io_input_bits_mask_20, // @[:@6.4]
  input        io_input_bits_mask_21, // @[:@6.4]
  input        io_input_bits_mask_22, // @[:@6.4]
  input        io_input_bits_mask_23, // @[:@6.4]
  input        io_input_bits_mask_24, // @[:@6.4]
  input        io_input_bits_mask_25, // @[:@6.4]
  input        io_input_bits_mask_26, // @[:@6.4]
  input        io_input_bits_mask_27, // @[:@6.4]
  input        io_input_bits_mask_28, // @[:@6.4]
  input        io_input_bits_mask_29, // @[:@6.4]
  input        io_input_bits_mask_30, // @[:@6.4]
  input        io_input_bits_mask_31, // @[:@6.4]
  input        io_input_bits_mask_32, // @[:@6.4]
  input        io_input_bits_mask_33, // @[:@6.4]
  input        io_input_bits_mask_34, // @[:@6.4]
  input        io_input_bits_mask_35, // @[:@6.4]
  input        io_input_bits_mask_36, // @[:@6.4]
  input        io_input_bits_mask_37, // @[:@6.4]
  input        io_input_bits_mask_38, // @[:@6.4]
  input        io_input_bits_mask_39, // @[:@6.4]
  input        io_input_bits_mask_40, // @[:@6.4]
  input        io_input_bits_mask_41, // @[:@6.4]
  input        io_input_bits_mask_42, // @[:@6.4]
  input        io_input_bits_mask_43, // @[:@6.4]
  input        io_input_bits_mask_44, // @[:@6.4]
  input        io_input_bits_mask_45, // @[:@6.4]
  input        io_input_bits_mask_46, // @[:@6.4]
  input        io_input_bits_mask_47, // @[:@6.4]
  input        io_input_bits_mask_48, // @[:@6.4]
  input        io_input_bits_mask_49, // @[:@6.4]
  input        io_input_bits_mask_50, // @[:@6.4]
  input        io_input_bits_mask_51, // @[:@6.4]
  input        io_input_bits_mask_52, // @[:@6.4]
  input        io_input_bits_mask_53, // @[:@6.4]
  input        io_input_bits_mask_54, // @[:@6.4]
  input        io_input_bits_mask_55, // @[:@6.4]
  input        io_input_bits_mask_56, // @[:@6.4]
  input        io_input_bits_mask_57, // @[:@6.4]
  input        io_input_bits_mask_58, // @[:@6.4]
  input        io_input_bits_mask_59, // @[:@6.4]
  input        io_input_bits_mask_60, // @[:@6.4]
  input        io_input_bits_mask_61, // @[:@6.4]
  input        io_input_bits_mask_62, // @[:@6.4]
  input        io_input_bits_mask_63, // @[:@6.4]
  input  [7:0] io_input_bits_data_0, // @[:@6.4]
  input  [7:0] io_input_bits_data_1, // @[:@6.4]
  input  [7:0] io_input_bits_data_2, // @[:@6.4]
  input  [7:0] io_input_bits_data_3, // @[:@6.4]
  input  [7:0] io_input_bits_data_4, // @[:@6.4]
  input  [7:0] io_input_bits_data_5, // @[:@6.4]
  input  [7:0] io_input_bits_data_6, // @[:@6.4]
  input  [7:0] io_input_bits_data_7, // @[:@6.4]
  input  [7:0] io_input_bits_data_8, // @[:@6.4]
  input  [7:0] io_input_bits_data_9, // @[:@6.4]
  input  [7:0] io_input_bits_data_10, // @[:@6.4]
  input  [7:0] io_input_bits_data_11, // @[:@6.4]
  input  [7:0] io_input_bits_data_12, // @[:@6.4]
  input  [7:0] io_input_bits_data_13, // @[:@6.4]
  input  [7:0] io_input_bits_data_14, // @[:@6.4]
  input  [7:0] io_input_bits_data_15, // @[:@6.4]
  input  [7:0] io_input_bits_data_16, // @[:@6.4]
  input  [7:0] io_input_bits_data_17, // @[:@6.4]
  input  [7:0] io_input_bits_data_18, // @[:@6.4]
  input  [7:0] io_input_bits_data_19, // @[:@6.4]
  input  [7:0] io_input_bits_data_20, // @[:@6.4]
  input  [7:0] io_input_bits_data_21, // @[:@6.4]
  input  [7:0] io_input_bits_data_22, // @[:@6.4]
  input  [7:0] io_input_bits_data_23, // @[:@6.4]
  input  [7:0] io_input_bits_data_24, // @[:@6.4]
  input  [7:0] io_input_bits_data_25, // @[:@6.4]
  input  [7:0] io_input_bits_data_26, // @[:@6.4]
  input  [7:0] io_input_bits_data_27, // @[:@6.4]
  input  [7:0] io_input_bits_data_28, // @[:@6.4]
  input  [7:0] io_input_bits_data_29, // @[:@6.4]
  input  [7:0] io_input_bits_data_30, // @[:@6.4]
  input  [7:0] io_input_bits_data_31, // @[:@6.4]
  input  [7:0] io_input_bits_data_32, // @[:@6.4]
  input  [7:0] io_input_bits_data_33, // @[:@6.4]
  input  [7:0] io_input_bits_data_34, // @[:@6.4]
  input  [7:0] io_input_bits_data_35, // @[:@6.4]
  input  [7:0] io_input_bits_data_36, // @[:@6.4]
  input  [7:0] io_input_bits_data_37, // @[:@6.4]
  input  [7:0] io_input_bits_data_38, // @[:@6.4]
  input  [7:0] io_input_bits_data_39, // @[:@6.4]
  input  [7:0] io_input_bits_data_40, // @[:@6.4]
  input  [7:0] io_input_bits_data_41, // @[:@6.4]
  input  [7:0] io_input_bits_data_42, // @[:@6.4]
  input  [7:0] io_input_bits_data_43, // @[:@6.4]
  input  [7:0] io_input_bits_data_44, // @[:@6.4]
  input  [7:0] io_input_bits_data_45, // @[:@6.4]
  input  [7:0] io_input_bits_data_46, // @[:@6.4]
  input  [7:0] io_input_bits_data_47, // @[:@6.4]
  input  [7:0] io_input_bits_data_48, // @[:@6.4]
  input  [7:0] io_input_bits_data_49, // @[:@6.4]
  input  [7:0] io_input_bits_data_50, // @[:@6.4]
  input  [7:0] io_input_bits_data_51, // @[:@6.4]
  input  [7:0] io_input_bits_data_52, // @[:@6.4]
  input  [7:0] io_input_bits_data_53, // @[:@6.4]
  input  [7:0] io_input_bits_data_54, // @[:@6.4]
  input  [7:0] io_input_bits_data_55, // @[:@6.4]
  input  [7:0] io_input_bits_data_56, // @[:@6.4]
  input  [7:0] io_input_bits_data_57, // @[:@6.4]
  input  [7:0] io_input_bits_data_58, // @[:@6.4]
  input  [7:0] io_input_bits_data_59, // @[:@6.4]
  input  [7:0] io_input_bits_data_60, // @[:@6.4]
  input  [7:0] io_input_bits_data_61, // @[:@6.4]
  input  [7:0] io_input_bits_data_62, // @[:@6.4]
  input  [7:0] io_input_bits_data_63, // @[:@6.4]
  input        io_input_bits_sel_0, // @[:@6.4]
  input        io_input_bits_sel_1, // @[:@6.4]
  input        io_input_bits_sel_2, // @[:@6.4]
  input        io_input_bits_sel_3, // @[:@6.4]
  input        io_input_bits_sel_4, // @[:@6.4]
  input        io_input_bits_sel_5, // @[:@6.4]
  input        io_input_bits_sel_6, // @[:@6.4]
  input        io_input_bits_sel_7, // @[:@6.4]
  input        io_input_bits_sel_8, // @[:@6.4]
  input        io_input_bits_sel_9, // @[:@6.4]
  input        io_input_bits_sel_10, // @[:@6.4]
  input        io_input_bits_sel_11, // @[:@6.4]
  input        io_input_bits_sel_12, // @[:@6.4]
  input        io_input_bits_sel_13, // @[:@6.4]
  input        io_input_bits_sel_14, // @[:@6.4]
  input        io_input_bits_sel_15, // @[:@6.4]
  input        io_input_bits_sel_16, // @[:@6.4]
  input        io_input_bits_sel_17, // @[:@6.4]
  input        io_input_bits_sel_18, // @[:@6.4]
  input        io_input_bits_sel_19, // @[:@6.4]
  input        io_input_bits_sel_20, // @[:@6.4]
  input        io_input_bits_sel_21, // @[:@6.4]
  input        io_input_bits_sel_22, // @[:@6.4]
  input        io_input_bits_sel_23, // @[:@6.4]
  input        io_input_bits_sel_24, // @[:@6.4]
  input        io_input_bits_sel_25, // @[:@6.4]
  input        io_input_bits_sel_26, // @[:@6.4]
  input        io_input_bits_sel_27, // @[:@6.4]
  input        io_input_bits_sel_28, // @[:@6.4]
  input        io_input_bits_sel_29, // @[:@6.4]
  input        io_input_bits_sel_30, // @[:@6.4]
  input        io_input_bits_sel_31, // @[:@6.4]
  input  [9:0] io_input_mask_en, // @[:@6.4]
  output       io_output_valid, // @[:@6.4]
  output       io_output_bits_mask_0, // @[:@6.4]
  output       io_output_bits_mask_1, // @[:@6.4]
  output       io_output_bits_mask_2, // @[:@6.4]
  output       io_output_bits_mask_3, // @[:@6.4]
  output       io_output_bits_mask_4, // @[:@6.4]
  output       io_output_bits_mask_5, // @[:@6.4]
  output       io_output_bits_mask_6, // @[:@6.4]
  output       io_output_bits_mask_7, // @[:@6.4]
  output       io_output_bits_mask_8, // @[:@6.4]
  output       io_output_bits_mask_9, // @[:@6.4]
  output       io_output_bits_mask_10, // @[:@6.4]
  output       io_output_bits_mask_11, // @[:@6.4]
  output       io_output_bits_mask_12, // @[:@6.4]
  output       io_output_bits_mask_13, // @[:@6.4]
  output       io_output_bits_mask_14, // @[:@6.4]
  output       io_output_bits_mask_15, // @[:@6.4]
  output       io_output_bits_mask_16, // @[:@6.4]
  output       io_output_bits_mask_17, // @[:@6.4]
  output       io_output_bits_mask_18, // @[:@6.4]
  output       io_output_bits_mask_19, // @[:@6.4]
  output       io_output_bits_mask_20, // @[:@6.4]
  output       io_output_bits_mask_21, // @[:@6.4]
  output       io_output_bits_mask_22, // @[:@6.4]
  output       io_output_bits_mask_23, // @[:@6.4]
  output       io_output_bits_mask_24, // @[:@6.4]
  output       io_output_bits_mask_25, // @[:@6.4]
  output       io_output_bits_mask_26, // @[:@6.4]
  output       io_output_bits_mask_27, // @[:@6.4]
  output       io_output_bits_mask_28, // @[:@6.4]
  output       io_output_bits_mask_29, // @[:@6.4]
  output       io_output_bits_mask_30, // @[:@6.4]
  output       io_output_bits_mask_31, // @[:@6.4]
  output       io_output_bits_mask_32, // @[:@6.4]
  output       io_output_bits_mask_33, // @[:@6.4]
  output       io_output_bits_mask_34, // @[:@6.4]
  output       io_output_bits_mask_35, // @[:@6.4]
  output       io_output_bits_mask_36, // @[:@6.4]
  output       io_output_bits_mask_37, // @[:@6.4]
  output       io_output_bits_mask_38, // @[:@6.4]
  output       io_output_bits_mask_39, // @[:@6.4]
  output       io_output_bits_mask_40, // @[:@6.4]
  output       io_output_bits_mask_41, // @[:@6.4]
  output       io_output_bits_mask_42, // @[:@6.4]
  output       io_output_bits_mask_43, // @[:@6.4]
  output       io_output_bits_mask_44, // @[:@6.4]
  output       io_output_bits_mask_45, // @[:@6.4]
  output       io_output_bits_mask_46, // @[:@6.4]
  output       io_output_bits_mask_47, // @[:@6.4]
  output       io_output_bits_mask_48, // @[:@6.4]
  output       io_output_bits_mask_49, // @[:@6.4]
  output       io_output_bits_mask_50, // @[:@6.4]
  output       io_output_bits_mask_51, // @[:@6.4]
  output       io_output_bits_mask_52, // @[:@6.4]
  output       io_output_bits_mask_53, // @[:@6.4]
  output       io_output_bits_mask_54, // @[:@6.4]
  output       io_output_bits_mask_55, // @[:@6.4]
  output       io_output_bits_mask_56, // @[:@6.4]
  output       io_output_bits_mask_57, // @[:@6.4]
  output       io_output_bits_mask_58, // @[:@6.4]
  output       io_output_bits_mask_59, // @[:@6.4]
  output       io_output_bits_mask_60, // @[:@6.4]
  output       io_output_bits_mask_61, // @[:@6.4]
  output       io_output_bits_mask_62, // @[:@6.4]
  output       io_output_bits_mask_63, // @[:@6.4]
  output [7:0] io_output_bits_data_0, // @[:@6.4]
  output [7:0] io_output_bits_data_1, // @[:@6.4]
  output [7:0] io_output_bits_data_2, // @[:@6.4]
  output [7:0] io_output_bits_data_3, // @[:@6.4]
  output [7:0] io_output_bits_data_4, // @[:@6.4]
  output [7:0] io_output_bits_data_5, // @[:@6.4]
  output [7:0] io_output_bits_data_6, // @[:@6.4]
  output [7:0] io_output_bits_data_7, // @[:@6.4]
  output [7:0] io_output_bits_data_8, // @[:@6.4]
  output [7:0] io_output_bits_data_9, // @[:@6.4]
  output [7:0] io_output_bits_data_10, // @[:@6.4]
  output [7:0] io_output_bits_data_11, // @[:@6.4]
  output [7:0] io_output_bits_data_12, // @[:@6.4]
  output [7:0] io_output_bits_data_13, // @[:@6.4]
  output [7:0] io_output_bits_data_14, // @[:@6.4]
  output [7:0] io_output_bits_data_15, // @[:@6.4]
  output [7:0] io_output_bits_data_16, // @[:@6.4]
  output [7:0] io_output_bits_data_17, // @[:@6.4]
  output [7:0] io_output_bits_data_18, // @[:@6.4]
  output [7:0] io_output_bits_data_19, // @[:@6.4]
  output [7:0] io_output_bits_data_20, // @[:@6.4]
  output [7:0] io_output_bits_data_21, // @[:@6.4]
  output [7:0] io_output_bits_data_22, // @[:@6.4]
  output [7:0] io_output_bits_data_23, // @[:@6.4]
  output [7:0] io_output_bits_data_24, // @[:@6.4]
  output [7:0] io_output_bits_data_25, // @[:@6.4]
  output [7:0] io_output_bits_data_26, // @[:@6.4]
  output [7:0] io_output_bits_data_27, // @[:@6.4]
  output [7:0] io_output_bits_data_28, // @[:@6.4]
  output [7:0] io_output_bits_data_29, // @[:@6.4]
  output [7:0] io_output_bits_data_30, // @[:@6.4]
  output [7:0] io_output_bits_data_31, // @[:@6.4]
  output [7:0] io_output_bits_data_32, // @[:@6.4]
  output [7:0] io_output_bits_data_33, // @[:@6.4]
  output [7:0] io_output_bits_data_34, // @[:@6.4]
  output [7:0] io_output_bits_data_35, // @[:@6.4]
  output [7:0] io_output_bits_data_36, // @[:@6.4]
  output [7:0] io_output_bits_data_37, // @[:@6.4]
  output [7:0] io_output_bits_data_38, // @[:@6.4]
  output [7:0] io_output_bits_data_39, // @[:@6.4]
  output [7:0] io_output_bits_data_40, // @[:@6.4]
  output [7:0] io_output_bits_data_41, // @[:@6.4]
  output [7:0] io_output_bits_data_42, // @[:@6.4]
  output [7:0] io_output_bits_data_43, // @[:@6.4]
  output [7:0] io_output_bits_data_44, // @[:@6.4]
  output [7:0] io_output_bits_data_45, // @[:@6.4]
  output [7:0] io_output_bits_data_46, // @[:@6.4]
  output [7:0] io_output_bits_data_47, // @[:@6.4]
  output [7:0] io_output_bits_data_48, // @[:@6.4]
  output [7:0] io_output_bits_data_49, // @[:@6.4]
  output [7:0] io_output_bits_data_50, // @[:@6.4]
  output [7:0] io_output_bits_data_51, // @[:@6.4]
  output [7:0] io_output_bits_data_52, // @[:@6.4]
  output [7:0] io_output_bits_data_53, // @[:@6.4]
  output [7:0] io_output_bits_data_54, // @[:@6.4]
  output [7:0] io_output_bits_data_55, // @[:@6.4]
  output [7:0] io_output_bits_data_56, // @[:@6.4]
  output [7:0] io_output_bits_data_57, // @[:@6.4]
  output [7:0] io_output_bits_data_58, // @[:@6.4]
  output [7:0] io_output_bits_data_59, // @[:@6.4]
  output [7:0] io_output_bits_data_60, // @[:@6.4]
  output [7:0] io_output_bits_data_61, // @[:@6.4]
  output [7:0] io_output_bits_data_62, // @[:@6.4]
  output [7:0] io_output_bits_data_63, // @[:@6.4]
  output       io_output_bits_sel_0, // @[:@6.4]
  output       io_output_bits_sel_1, // @[:@6.4]
  output       io_output_bits_sel_2, // @[:@6.4]
  output       io_output_bits_sel_3, // @[:@6.4]
  output       io_output_bits_sel_4, // @[:@6.4]
  output       io_output_bits_sel_5, // @[:@6.4]
  output       io_output_bits_sel_6, // @[:@6.4]
  output       io_output_bits_sel_7, // @[:@6.4]
  output       io_output_bits_sel_8, // @[:@6.4]
  output       io_output_bits_sel_9, // @[:@6.4]
  output       io_output_bits_sel_10, // @[:@6.4]
  output       io_output_bits_sel_11, // @[:@6.4]
  output       io_output_bits_sel_12, // @[:@6.4]
  output       io_output_bits_sel_13, // @[:@6.4]
  output       io_output_bits_sel_14, // @[:@6.4]
  output       io_output_bits_sel_15, // @[:@6.4]
  output       io_output_bits_sel_16, // @[:@6.4]
  output       io_output_bits_sel_17, // @[:@6.4]
  output       io_output_bits_sel_18, // @[:@6.4]
  output       io_output_bits_sel_19, // @[:@6.4]
  output       io_output_bits_sel_20, // @[:@6.4]
  output       io_output_bits_sel_21, // @[:@6.4]
  output       io_output_bits_sel_22, // @[:@6.4]
  output       io_output_bits_sel_23, // @[:@6.4]
  output       io_output_bits_sel_24, // @[:@6.4]
  output       io_output_bits_sel_25, // @[:@6.4]
  output       io_output_bits_sel_26, // @[:@6.4]
  output       io_output_bits_sel_27, // @[:@6.4]
  output       io_output_bits_sel_28, // @[:@6.4]
  output       io_output_bits_sel_29, // @[:@6.4]
  output       io_output_bits_sel_30, // @[:@6.4]
  output       io_output_bits_sel_31 // @[:@6.4]
);
  wire  _T_1771; // @[NV_NVDLA_CSC_WL_dec.scala 56:48:@8.4]
  wire  _T_1906_0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_1; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_2; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_3; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_4; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_5; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_6; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_7; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_8; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_9; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_10; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_11; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_12; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_13; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_14; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_15; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_16; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_17; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_18; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_19; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_20; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_21; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_22; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_23; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_24; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_25; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_26; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_27; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_28; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_29; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_30; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_31; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_32; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_33; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_34; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_35; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_36; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_37; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_38; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_39; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_40; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_41; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_42; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_43; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_44; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_45; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_46; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_47; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_48; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_49; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_50; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_51; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_52; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_53; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_54; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_55; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_56; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_57; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_58; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_59; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_60; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_61; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_62; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire  _T_1906_63; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  wire [7:0] _T_2174; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@82.4]
  wire [15:0] _T_2182; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@90.4]
  wire [7:0] _T_2189; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@97.4]
  wire [31:0] _T_2198; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@106.4]
  wire [7:0] _T_2205; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@113.4]
  wire [15:0] _T_2213; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@121.4]
  wire [7:0] _T_2220; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@128.4]
  wire [31:0] _T_2229; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@137.4]
  wire [63:0] _T_2230; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@138.4]
  wire  _T_2231; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@139.4]
  wire [1:0] _T_2296; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@205.4]
  wire  _T_2297; // @[Bitwise.scala 50:65:@206.4]
  wire  _T_2298; // @[Bitwise.scala 50:65:@207.4]
  wire [1:0] _T_2299; // @[Bitwise.scala 48:55:@208.4]
  wire [2:0] _T_2363; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@273.4]
  wire  _T_2364; // @[Bitwise.scala 50:65:@274.4]
  wire  _T_2365; // @[Bitwise.scala 50:65:@275.4]
  wire  _T_2366; // @[Bitwise.scala 50:65:@276.4]
  wire [1:0] _T_2367; // @[Bitwise.scala 48:55:@277.4]
  wire [1:0] _GEN_544; // @[Bitwise.scala 48:55:@278.4]
  wire [2:0] _T_2368; // @[Bitwise.scala 48:55:@278.4]
  wire [3:0] _T_2432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@343.4]
  wire  _T_2433; // @[Bitwise.scala 50:65:@344.4]
  wire  _T_2434; // @[Bitwise.scala 50:65:@345.4]
  wire  _T_2435; // @[Bitwise.scala 50:65:@346.4]
  wire  _T_2436; // @[Bitwise.scala 50:65:@347.4]
  wire [1:0] _T_2437; // @[Bitwise.scala 48:55:@348.4]
  wire [1:0] _T_2438; // @[Bitwise.scala 48:55:@349.4]
  wire [2:0] _T_2439; // @[Bitwise.scala 48:55:@350.4]
  wire [4:0] _T_2503; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@415.4]
  wire  _T_2504; // @[Bitwise.scala 50:65:@416.4]
  wire  _T_2505; // @[Bitwise.scala 50:65:@417.4]
  wire  _T_2506; // @[Bitwise.scala 50:65:@418.4]
  wire  _T_2507; // @[Bitwise.scala 50:65:@419.4]
  wire  _T_2508; // @[Bitwise.scala 50:65:@420.4]
  wire [1:0] _T_2509; // @[Bitwise.scala 48:55:@421.4]
  wire [1:0] _T_2510; // @[Bitwise.scala 48:55:@422.4]
  wire [1:0] _GEN_545; // @[Bitwise.scala 48:55:@423.4]
  wire [2:0] _T_2511; // @[Bitwise.scala 48:55:@423.4]
  wire [2:0] _GEN_546; // @[Bitwise.scala 48:55:@424.4]
  wire [3:0] _T_2512; // @[Bitwise.scala 48:55:@424.4]
  wire [5:0] _T_2576; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@489.4]
  wire  _T_2577; // @[Bitwise.scala 50:65:@490.4]
  wire  _T_2578; // @[Bitwise.scala 50:65:@491.4]
  wire  _T_2579; // @[Bitwise.scala 50:65:@492.4]
  wire  _T_2580; // @[Bitwise.scala 50:65:@493.4]
  wire  _T_2581; // @[Bitwise.scala 50:65:@494.4]
  wire  _T_2582; // @[Bitwise.scala 50:65:@495.4]
  wire [1:0] _T_2583; // @[Bitwise.scala 48:55:@496.4]
  wire [1:0] _GEN_547; // @[Bitwise.scala 48:55:@497.4]
  wire [2:0] _T_2584; // @[Bitwise.scala 48:55:@497.4]
  wire [1:0] _T_2585; // @[Bitwise.scala 48:55:@498.4]
  wire [1:0] _GEN_548; // @[Bitwise.scala 48:55:@499.4]
  wire [2:0] _T_2586; // @[Bitwise.scala 48:55:@499.4]
  wire [3:0] _T_2587; // @[Bitwise.scala 48:55:@500.4]
  wire [6:0] _T_2651; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@565.4]
  wire  _T_2652; // @[Bitwise.scala 50:65:@566.4]
  wire  _T_2653; // @[Bitwise.scala 50:65:@567.4]
  wire  _T_2654; // @[Bitwise.scala 50:65:@568.4]
  wire  _T_2655; // @[Bitwise.scala 50:65:@569.4]
  wire  _T_2656; // @[Bitwise.scala 50:65:@570.4]
  wire  _T_2657; // @[Bitwise.scala 50:65:@571.4]
  wire  _T_2658; // @[Bitwise.scala 50:65:@572.4]
  wire [1:0] _T_2659; // @[Bitwise.scala 48:55:@573.4]
  wire [1:0] _GEN_549; // @[Bitwise.scala 48:55:@574.4]
  wire [2:0] _T_2660; // @[Bitwise.scala 48:55:@574.4]
  wire [1:0] _T_2661; // @[Bitwise.scala 48:55:@575.4]
  wire [1:0] _T_2662; // @[Bitwise.scala 48:55:@576.4]
  wire [2:0] _T_2663; // @[Bitwise.scala 48:55:@577.4]
  wire [3:0] _T_2664; // @[Bitwise.scala 48:55:@578.4]
  wire [7:0] _T_2728; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@643.4]
  wire  _T_2729; // @[Bitwise.scala 50:65:@644.4]
  wire  _T_2730; // @[Bitwise.scala 50:65:@645.4]
  wire  _T_2731; // @[Bitwise.scala 50:65:@646.4]
  wire  _T_2732; // @[Bitwise.scala 50:65:@647.4]
  wire  _T_2733; // @[Bitwise.scala 50:65:@648.4]
  wire  _T_2734; // @[Bitwise.scala 50:65:@649.4]
  wire  _T_2735; // @[Bitwise.scala 50:65:@650.4]
  wire  _T_2736; // @[Bitwise.scala 50:65:@651.4]
  wire [1:0] _T_2737; // @[Bitwise.scala 48:55:@652.4]
  wire [1:0] _T_2738; // @[Bitwise.scala 48:55:@653.4]
  wire [2:0] _T_2739; // @[Bitwise.scala 48:55:@654.4]
  wire [1:0] _T_2740; // @[Bitwise.scala 48:55:@655.4]
  wire [1:0] _T_2741; // @[Bitwise.scala 48:55:@656.4]
  wire [2:0] _T_2742; // @[Bitwise.scala 48:55:@657.4]
  wire [3:0] _T_2743; // @[Bitwise.scala 48:55:@658.4]
  wire [8:0] _T_2807; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@723.4]
  wire  _T_2808; // @[Bitwise.scala 50:65:@724.4]
  wire  _T_2809; // @[Bitwise.scala 50:65:@725.4]
  wire  _T_2810; // @[Bitwise.scala 50:65:@726.4]
  wire  _T_2811; // @[Bitwise.scala 50:65:@727.4]
  wire  _T_2812; // @[Bitwise.scala 50:65:@728.4]
  wire  _T_2813; // @[Bitwise.scala 50:65:@729.4]
  wire  _T_2814; // @[Bitwise.scala 50:65:@730.4]
  wire  _T_2815; // @[Bitwise.scala 50:65:@731.4]
  wire  _T_2816; // @[Bitwise.scala 50:65:@732.4]
  wire [1:0] _T_2817; // @[Bitwise.scala 48:55:@733.4]
  wire [1:0] _T_2818; // @[Bitwise.scala 48:55:@734.4]
  wire [2:0] _T_2819; // @[Bitwise.scala 48:55:@735.4]
  wire [1:0] _T_2820; // @[Bitwise.scala 48:55:@736.4]
  wire [1:0] _T_2821; // @[Bitwise.scala 48:55:@737.4]
  wire [1:0] _GEN_550; // @[Bitwise.scala 48:55:@738.4]
  wire [2:0] _T_2822; // @[Bitwise.scala 48:55:@738.4]
  wire [2:0] _GEN_551; // @[Bitwise.scala 48:55:@739.4]
  wire [3:0] _T_2823; // @[Bitwise.scala 48:55:@739.4]
  wire [3:0] _GEN_552; // @[Bitwise.scala 48:55:@740.4]
  wire [4:0] _T_2824; // @[Bitwise.scala 48:55:@740.4]
  wire [9:0] _T_2888; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@805.4]
  wire  _T_2889; // @[Bitwise.scala 50:65:@806.4]
  wire  _T_2890; // @[Bitwise.scala 50:65:@807.4]
  wire  _T_2891; // @[Bitwise.scala 50:65:@808.4]
  wire  _T_2892; // @[Bitwise.scala 50:65:@809.4]
  wire  _T_2893; // @[Bitwise.scala 50:65:@810.4]
  wire  _T_2894; // @[Bitwise.scala 50:65:@811.4]
  wire  _T_2895; // @[Bitwise.scala 50:65:@812.4]
  wire  _T_2896; // @[Bitwise.scala 50:65:@813.4]
  wire  _T_2897; // @[Bitwise.scala 50:65:@814.4]
  wire  _T_2898; // @[Bitwise.scala 50:65:@815.4]
  wire [1:0] _T_2899; // @[Bitwise.scala 48:55:@816.4]
  wire [1:0] _T_2900; // @[Bitwise.scala 48:55:@817.4]
  wire [1:0] _GEN_553; // @[Bitwise.scala 48:55:@818.4]
  wire [2:0] _T_2901; // @[Bitwise.scala 48:55:@818.4]
  wire [2:0] _GEN_554; // @[Bitwise.scala 48:55:@819.4]
  wire [3:0] _T_2902; // @[Bitwise.scala 48:55:@819.4]
  wire [1:0] _T_2903; // @[Bitwise.scala 48:55:@820.4]
  wire [1:0] _T_2904; // @[Bitwise.scala 48:55:@821.4]
  wire [1:0] _GEN_555; // @[Bitwise.scala 48:55:@822.4]
  wire [2:0] _T_2905; // @[Bitwise.scala 48:55:@822.4]
  wire [2:0] _GEN_556; // @[Bitwise.scala 48:55:@823.4]
  wire [3:0] _T_2906; // @[Bitwise.scala 48:55:@823.4]
  wire [4:0] _T_2907; // @[Bitwise.scala 48:55:@824.4]
  wire [10:0] _T_2971; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@889.4]
  wire  _T_2972; // @[Bitwise.scala 50:65:@890.4]
  wire  _T_2973; // @[Bitwise.scala 50:65:@891.4]
  wire  _T_2974; // @[Bitwise.scala 50:65:@892.4]
  wire  _T_2975; // @[Bitwise.scala 50:65:@893.4]
  wire  _T_2976; // @[Bitwise.scala 50:65:@894.4]
  wire  _T_2977; // @[Bitwise.scala 50:65:@895.4]
  wire  _T_2978; // @[Bitwise.scala 50:65:@896.4]
  wire  _T_2979; // @[Bitwise.scala 50:65:@897.4]
  wire  _T_2980; // @[Bitwise.scala 50:65:@898.4]
  wire  _T_2981; // @[Bitwise.scala 50:65:@899.4]
  wire  _T_2982; // @[Bitwise.scala 50:65:@900.4]
  wire [1:0] _T_2983; // @[Bitwise.scala 48:55:@901.4]
  wire [1:0] _T_2984; // @[Bitwise.scala 48:55:@902.4]
  wire [1:0] _GEN_557; // @[Bitwise.scala 48:55:@903.4]
  wire [2:0] _T_2985; // @[Bitwise.scala 48:55:@903.4]
  wire [2:0] _GEN_558; // @[Bitwise.scala 48:55:@904.4]
  wire [3:0] _T_2986; // @[Bitwise.scala 48:55:@904.4]
  wire [1:0] _T_2987; // @[Bitwise.scala 48:55:@905.4]
  wire [1:0] _GEN_559; // @[Bitwise.scala 48:55:@906.4]
  wire [2:0] _T_2988; // @[Bitwise.scala 48:55:@906.4]
  wire [1:0] _T_2989; // @[Bitwise.scala 48:55:@907.4]
  wire [1:0] _GEN_560; // @[Bitwise.scala 48:55:@908.4]
  wire [2:0] _T_2990; // @[Bitwise.scala 48:55:@908.4]
  wire [3:0] _T_2991; // @[Bitwise.scala 48:55:@909.4]
  wire [4:0] _T_2992; // @[Bitwise.scala 48:55:@910.4]
  wire [11:0] _T_3056; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@975.4]
  wire  _T_3057; // @[Bitwise.scala 50:65:@976.4]
  wire  _T_3058; // @[Bitwise.scala 50:65:@977.4]
  wire  _T_3059; // @[Bitwise.scala 50:65:@978.4]
  wire  _T_3060; // @[Bitwise.scala 50:65:@979.4]
  wire  _T_3061; // @[Bitwise.scala 50:65:@980.4]
  wire  _T_3062; // @[Bitwise.scala 50:65:@981.4]
  wire  _T_3063; // @[Bitwise.scala 50:65:@982.4]
  wire  _T_3064; // @[Bitwise.scala 50:65:@983.4]
  wire  _T_3065; // @[Bitwise.scala 50:65:@984.4]
  wire  _T_3066; // @[Bitwise.scala 50:65:@985.4]
  wire  _T_3067; // @[Bitwise.scala 50:65:@986.4]
  wire  _T_3068; // @[Bitwise.scala 50:65:@987.4]
  wire [1:0] _T_3069; // @[Bitwise.scala 48:55:@988.4]
  wire [1:0] _GEN_561; // @[Bitwise.scala 48:55:@989.4]
  wire [2:0] _T_3070; // @[Bitwise.scala 48:55:@989.4]
  wire [1:0] _T_3071; // @[Bitwise.scala 48:55:@990.4]
  wire [1:0] _GEN_562; // @[Bitwise.scala 48:55:@991.4]
  wire [2:0] _T_3072; // @[Bitwise.scala 48:55:@991.4]
  wire [3:0] _T_3073; // @[Bitwise.scala 48:55:@992.4]
  wire [1:0] _T_3074; // @[Bitwise.scala 48:55:@993.4]
  wire [1:0] _GEN_563; // @[Bitwise.scala 48:55:@994.4]
  wire [2:0] _T_3075; // @[Bitwise.scala 48:55:@994.4]
  wire [1:0] _T_3076; // @[Bitwise.scala 48:55:@995.4]
  wire [1:0] _GEN_564; // @[Bitwise.scala 48:55:@996.4]
  wire [2:0] _T_3077; // @[Bitwise.scala 48:55:@996.4]
  wire [3:0] _T_3078; // @[Bitwise.scala 48:55:@997.4]
  wire [4:0] _T_3079; // @[Bitwise.scala 48:55:@998.4]
  wire [12:0] _T_3143; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1063.4]
  wire  _T_3144; // @[Bitwise.scala 50:65:@1064.4]
  wire  _T_3145; // @[Bitwise.scala 50:65:@1065.4]
  wire  _T_3146; // @[Bitwise.scala 50:65:@1066.4]
  wire  _T_3147; // @[Bitwise.scala 50:65:@1067.4]
  wire  _T_3148; // @[Bitwise.scala 50:65:@1068.4]
  wire  _T_3149; // @[Bitwise.scala 50:65:@1069.4]
  wire  _T_3150; // @[Bitwise.scala 50:65:@1070.4]
  wire  _T_3151; // @[Bitwise.scala 50:65:@1071.4]
  wire  _T_3152; // @[Bitwise.scala 50:65:@1072.4]
  wire  _T_3153; // @[Bitwise.scala 50:65:@1073.4]
  wire  _T_3154; // @[Bitwise.scala 50:65:@1074.4]
  wire  _T_3155; // @[Bitwise.scala 50:65:@1075.4]
  wire  _T_3156; // @[Bitwise.scala 50:65:@1076.4]
  wire [1:0] _T_3157; // @[Bitwise.scala 48:55:@1077.4]
  wire [1:0] _GEN_565; // @[Bitwise.scala 48:55:@1078.4]
  wire [2:0] _T_3158; // @[Bitwise.scala 48:55:@1078.4]
  wire [1:0] _T_3159; // @[Bitwise.scala 48:55:@1079.4]
  wire [1:0] _GEN_566; // @[Bitwise.scala 48:55:@1080.4]
  wire [2:0] _T_3160; // @[Bitwise.scala 48:55:@1080.4]
  wire [3:0] _T_3161; // @[Bitwise.scala 48:55:@1081.4]
  wire [1:0] _T_3162; // @[Bitwise.scala 48:55:@1082.4]
  wire [1:0] _GEN_567; // @[Bitwise.scala 48:55:@1083.4]
  wire [2:0] _T_3163; // @[Bitwise.scala 48:55:@1083.4]
  wire [1:0] _T_3164; // @[Bitwise.scala 48:55:@1084.4]
  wire [1:0] _T_3165; // @[Bitwise.scala 48:55:@1085.4]
  wire [2:0] _T_3166; // @[Bitwise.scala 48:55:@1086.4]
  wire [3:0] _T_3167; // @[Bitwise.scala 48:55:@1087.4]
  wire [4:0] _T_3168; // @[Bitwise.scala 48:55:@1088.4]
  wire [13:0] _T_3232; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1153.4]
  wire  _T_3233; // @[Bitwise.scala 50:65:@1154.4]
  wire  _T_3234; // @[Bitwise.scala 50:65:@1155.4]
  wire  _T_3235; // @[Bitwise.scala 50:65:@1156.4]
  wire  _T_3236; // @[Bitwise.scala 50:65:@1157.4]
  wire  _T_3237; // @[Bitwise.scala 50:65:@1158.4]
  wire  _T_3238; // @[Bitwise.scala 50:65:@1159.4]
  wire  _T_3239; // @[Bitwise.scala 50:65:@1160.4]
  wire  _T_3240; // @[Bitwise.scala 50:65:@1161.4]
  wire  _T_3241; // @[Bitwise.scala 50:65:@1162.4]
  wire  _T_3242; // @[Bitwise.scala 50:65:@1163.4]
  wire  _T_3243; // @[Bitwise.scala 50:65:@1164.4]
  wire  _T_3244; // @[Bitwise.scala 50:65:@1165.4]
  wire  _T_3245; // @[Bitwise.scala 50:65:@1166.4]
  wire  _T_3246; // @[Bitwise.scala 50:65:@1167.4]
  wire [1:0] _T_3247; // @[Bitwise.scala 48:55:@1168.4]
  wire [1:0] _GEN_568; // @[Bitwise.scala 48:55:@1169.4]
  wire [2:0] _T_3248; // @[Bitwise.scala 48:55:@1169.4]
  wire [1:0] _T_3249; // @[Bitwise.scala 48:55:@1170.4]
  wire [1:0] _T_3250; // @[Bitwise.scala 48:55:@1171.4]
  wire [2:0] _T_3251; // @[Bitwise.scala 48:55:@1172.4]
  wire [3:0] _T_3252; // @[Bitwise.scala 48:55:@1173.4]
  wire [1:0] _T_3253; // @[Bitwise.scala 48:55:@1174.4]
  wire [1:0] _GEN_569; // @[Bitwise.scala 48:55:@1175.4]
  wire [2:0] _T_3254; // @[Bitwise.scala 48:55:@1175.4]
  wire [1:0] _T_3255; // @[Bitwise.scala 48:55:@1176.4]
  wire [1:0] _T_3256; // @[Bitwise.scala 48:55:@1177.4]
  wire [2:0] _T_3257; // @[Bitwise.scala 48:55:@1178.4]
  wire [3:0] _T_3258; // @[Bitwise.scala 48:55:@1179.4]
  wire [4:0] _T_3259; // @[Bitwise.scala 48:55:@1180.4]
  wire [14:0] _T_3323; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1245.4]
  wire  _T_3324; // @[Bitwise.scala 50:65:@1246.4]
  wire  _T_3325; // @[Bitwise.scala 50:65:@1247.4]
  wire  _T_3326; // @[Bitwise.scala 50:65:@1248.4]
  wire  _T_3327; // @[Bitwise.scala 50:65:@1249.4]
  wire  _T_3328; // @[Bitwise.scala 50:65:@1250.4]
  wire  _T_3329; // @[Bitwise.scala 50:65:@1251.4]
  wire  _T_3330; // @[Bitwise.scala 50:65:@1252.4]
  wire  _T_3331; // @[Bitwise.scala 50:65:@1253.4]
  wire  _T_3332; // @[Bitwise.scala 50:65:@1254.4]
  wire  _T_3333; // @[Bitwise.scala 50:65:@1255.4]
  wire  _T_3334; // @[Bitwise.scala 50:65:@1256.4]
  wire  _T_3335; // @[Bitwise.scala 50:65:@1257.4]
  wire  _T_3336; // @[Bitwise.scala 50:65:@1258.4]
  wire  _T_3337; // @[Bitwise.scala 50:65:@1259.4]
  wire  _T_3338; // @[Bitwise.scala 50:65:@1260.4]
  wire [1:0] _T_3339; // @[Bitwise.scala 48:55:@1261.4]
  wire [1:0] _GEN_570; // @[Bitwise.scala 48:55:@1262.4]
  wire [2:0] _T_3340; // @[Bitwise.scala 48:55:@1262.4]
  wire [1:0] _T_3341; // @[Bitwise.scala 48:55:@1263.4]
  wire [1:0] _T_3342; // @[Bitwise.scala 48:55:@1264.4]
  wire [2:0] _T_3343; // @[Bitwise.scala 48:55:@1265.4]
  wire [3:0] _T_3344; // @[Bitwise.scala 48:55:@1266.4]
  wire [1:0] _T_3345; // @[Bitwise.scala 48:55:@1267.4]
  wire [1:0] _T_3346; // @[Bitwise.scala 48:55:@1268.4]
  wire [2:0] _T_3347; // @[Bitwise.scala 48:55:@1269.4]
  wire [1:0] _T_3348; // @[Bitwise.scala 48:55:@1270.4]
  wire [1:0] _T_3349; // @[Bitwise.scala 48:55:@1271.4]
  wire [2:0] _T_3350; // @[Bitwise.scala 48:55:@1272.4]
  wire [3:0] _T_3351; // @[Bitwise.scala 48:55:@1273.4]
  wire [4:0] _T_3352; // @[Bitwise.scala 48:55:@1274.4]
  wire [15:0] _T_3416; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1339.4]
  wire  _T_3417; // @[Bitwise.scala 50:65:@1340.4]
  wire  _T_3418; // @[Bitwise.scala 50:65:@1341.4]
  wire  _T_3419; // @[Bitwise.scala 50:65:@1342.4]
  wire  _T_3420; // @[Bitwise.scala 50:65:@1343.4]
  wire  _T_3421; // @[Bitwise.scala 50:65:@1344.4]
  wire  _T_3422; // @[Bitwise.scala 50:65:@1345.4]
  wire  _T_3423; // @[Bitwise.scala 50:65:@1346.4]
  wire  _T_3424; // @[Bitwise.scala 50:65:@1347.4]
  wire  _T_3425; // @[Bitwise.scala 50:65:@1348.4]
  wire  _T_3426; // @[Bitwise.scala 50:65:@1349.4]
  wire  _T_3427; // @[Bitwise.scala 50:65:@1350.4]
  wire  _T_3428; // @[Bitwise.scala 50:65:@1351.4]
  wire  _T_3429; // @[Bitwise.scala 50:65:@1352.4]
  wire  _T_3430; // @[Bitwise.scala 50:65:@1353.4]
  wire  _T_3431; // @[Bitwise.scala 50:65:@1354.4]
  wire  _T_3432; // @[Bitwise.scala 50:65:@1355.4]
  wire [1:0] _T_3433; // @[Bitwise.scala 48:55:@1356.4]
  wire [1:0] _T_3434; // @[Bitwise.scala 48:55:@1357.4]
  wire [2:0] _T_3435; // @[Bitwise.scala 48:55:@1358.4]
  wire [1:0] _T_3436; // @[Bitwise.scala 48:55:@1359.4]
  wire [1:0] _T_3437; // @[Bitwise.scala 48:55:@1360.4]
  wire [2:0] _T_3438; // @[Bitwise.scala 48:55:@1361.4]
  wire [3:0] _T_3439; // @[Bitwise.scala 48:55:@1362.4]
  wire [1:0] _T_3440; // @[Bitwise.scala 48:55:@1363.4]
  wire [1:0] _T_3441; // @[Bitwise.scala 48:55:@1364.4]
  wire [2:0] _T_3442; // @[Bitwise.scala 48:55:@1365.4]
  wire [1:0] _T_3443; // @[Bitwise.scala 48:55:@1366.4]
  wire [1:0] _T_3444; // @[Bitwise.scala 48:55:@1367.4]
  wire [2:0] _T_3445; // @[Bitwise.scala 48:55:@1368.4]
  wire [3:0] _T_3446; // @[Bitwise.scala 48:55:@1369.4]
  wire [4:0] _T_3447; // @[Bitwise.scala 48:55:@1370.4]
  wire [16:0] _T_3511; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1435.4]
  wire  _T_3512; // @[Bitwise.scala 50:65:@1436.4]
  wire  _T_3513; // @[Bitwise.scala 50:65:@1437.4]
  wire  _T_3514; // @[Bitwise.scala 50:65:@1438.4]
  wire  _T_3515; // @[Bitwise.scala 50:65:@1439.4]
  wire  _T_3516; // @[Bitwise.scala 50:65:@1440.4]
  wire  _T_3517; // @[Bitwise.scala 50:65:@1441.4]
  wire  _T_3518; // @[Bitwise.scala 50:65:@1442.4]
  wire  _T_3519; // @[Bitwise.scala 50:65:@1443.4]
  wire  _T_3520; // @[Bitwise.scala 50:65:@1444.4]
  wire  _T_3521; // @[Bitwise.scala 50:65:@1445.4]
  wire  _T_3522; // @[Bitwise.scala 50:65:@1446.4]
  wire  _T_3523; // @[Bitwise.scala 50:65:@1447.4]
  wire  _T_3524; // @[Bitwise.scala 50:65:@1448.4]
  wire  _T_3525; // @[Bitwise.scala 50:65:@1449.4]
  wire  _T_3526; // @[Bitwise.scala 50:65:@1450.4]
  wire  _T_3527; // @[Bitwise.scala 50:65:@1451.4]
  wire  _T_3528; // @[Bitwise.scala 50:65:@1452.4]
  wire [1:0] _T_3529; // @[Bitwise.scala 48:55:@1453.4]
  wire [1:0] _T_3530; // @[Bitwise.scala 48:55:@1454.4]
  wire [2:0] _T_3531; // @[Bitwise.scala 48:55:@1455.4]
  wire [1:0] _T_3532; // @[Bitwise.scala 48:55:@1456.4]
  wire [1:0] _T_3533; // @[Bitwise.scala 48:55:@1457.4]
  wire [2:0] _T_3534; // @[Bitwise.scala 48:55:@1458.4]
  wire [3:0] _T_3535; // @[Bitwise.scala 48:55:@1459.4]
  wire [1:0] _T_3536; // @[Bitwise.scala 48:55:@1460.4]
  wire [1:0] _T_3537; // @[Bitwise.scala 48:55:@1461.4]
  wire [2:0] _T_3538; // @[Bitwise.scala 48:55:@1462.4]
  wire [1:0] _T_3539; // @[Bitwise.scala 48:55:@1463.4]
  wire [1:0] _T_3540; // @[Bitwise.scala 48:55:@1464.4]
  wire [1:0] _GEN_571; // @[Bitwise.scala 48:55:@1465.4]
  wire [2:0] _T_3541; // @[Bitwise.scala 48:55:@1465.4]
  wire [2:0] _GEN_572; // @[Bitwise.scala 48:55:@1466.4]
  wire [3:0] _T_3542; // @[Bitwise.scala 48:55:@1466.4]
  wire [3:0] _GEN_573; // @[Bitwise.scala 48:55:@1467.4]
  wire [4:0] _T_3543; // @[Bitwise.scala 48:55:@1467.4]
  wire [4:0] _GEN_574; // @[Bitwise.scala 48:55:@1468.4]
  wire [5:0] _T_3544; // @[Bitwise.scala 48:55:@1468.4]
  wire [17:0] _T_3608; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1533.4]
  wire  _T_3609; // @[Bitwise.scala 50:65:@1534.4]
  wire  _T_3610; // @[Bitwise.scala 50:65:@1535.4]
  wire  _T_3611; // @[Bitwise.scala 50:65:@1536.4]
  wire  _T_3612; // @[Bitwise.scala 50:65:@1537.4]
  wire  _T_3613; // @[Bitwise.scala 50:65:@1538.4]
  wire  _T_3614; // @[Bitwise.scala 50:65:@1539.4]
  wire  _T_3615; // @[Bitwise.scala 50:65:@1540.4]
  wire  _T_3616; // @[Bitwise.scala 50:65:@1541.4]
  wire  _T_3617; // @[Bitwise.scala 50:65:@1542.4]
  wire  _T_3618; // @[Bitwise.scala 50:65:@1543.4]
  wire  _T_3619; // @[Bitwise.scala 50:65:@1544.4]
  wire  _T_3620; // @[Bitwise.scala 50:65:@1545.4]
  wire  _T_3621; // @[Bitwise.scala 50:65:@1546.4]
  wire  _T_3622; // @[Bitwise.scala 50:65:@1547.4]
  wire  _T_3623; // @[Bitwise.scala 50:65:@1548.4]
  wire  _T_3624; // @[Bitwise.scala 50:65:@1549.4]
  wire  _T_3625; // @[Bitwise.scala 50:65:@1550.4]
  wire  _T_3626; // @[Bitwise.scala 50:65:@1551.4]
  wire [1:0] _T_3627; // @[Bitwise.scala 48:55:@1552.4]
  wire [1:0] _T_3628; // @[Bitwise.scala 48:55:@1553.4]
  wire [2:0] _T_3629; // @[Bitwise.scala 48:55:@1554.4]
  wire [1:0] _T_3630; // @[Bitwise.scala 48:55:@1555.4]
  wire [1:0] _T_3631; // @[Bitwise.scala 48:55:@1556.4]
  wire [1:0] _GEN_575; // @[Bitwise.scala 48:55:@1557.4]
  wire [2:0] _T_3632; // @[Bitwise.scala 48:55:@1557.4]
  wire [2:0] _GEN_576; // @[Bitwise.scala 48:55:@1558.4]
  wire [3:0] _T_3633; // @[Bitwise.scala 48:55:@1558.4]
  wire [3:0] _GEN_577; // @[Bitwise.scala 48:55:@1559.4]
  wire [4:0] _T_3634; // @[Bitwise.scala 48:55:@1559.4]
  wire [1:0] _T_3635; // @[Bitwise.scala 48:55:@1560.4]
  wire [1:0] _T_3636; // @[Bitwise.scala 48:55:@1561.4]
  wire [2:0] _T_3637; // @[Bitwise.scala 48:55:@1562.4]
  wire [1:0] _T_3638; // @[Bitwise.scala 48:55:@1563.4]
  wire [1:0] _T_3639; // @[Bitwise.scala 48:55:@1564.4]
  wire [1:0] _GEN_578; // @[Bitwise.scala 48:55:@1565.4]
  wire [2:0] _T_3640; // @[Bitwise.scala 48:55:@1565.4]
  wire [2:0] _GEN_579; // @[Bitwise.scala 48:55:@1566.4]
  wire [3:0] _T_3641; // @[Bitwise.scala 48:55:@1566.4]
  wire [3:0] _GEN_580; // @[Bitwise.scala 48:55:@1567.4]
  wire [4:0] _T_3642; // @[Bitwise.scala 48:55:@1567.4]
  wire [5:0] _T_3643; // @[Bitwise.scala 48:55:@1568.4]
  wire [18:0] _T_3707; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1633.4]
  wire  _T_3708; // @[Bitwise.scala 50:65:@1634.4]
  wire  _T_3709; // @[Bitwise.scala 50:65:@1635.4]
  wire  _T_3710; // @[Bitwise.scala 50:65:@1636.4]
  wire  _T_3711; // @[Bitwise.scala 50:65:@1637.4]
  wire  _T_3712; // @[Bitwise.scala 50:65:@1638.4]
  wire  _T_3713; // @[Bitwise.scala 50:65:@1639.4]
  wire  _T_3714; // @[Bitwise.scala 50:65:@1640.4]
  wire  _T_3715; // @[Bitwise.scala 50:65:@1641.4]
  wire  _T_3716; // @[Bitwise.scala 50:65:@1642.4]
  wire  _T_3717; // @[Bitwise.scala 50:65:@1643.4]
  wire  _T_3718; // @[Bitwise.scala 50:65:@1644.4]
  wire  _T_3719; // @[Bitwise.scala 50:65:@1645.4]
  wire  _T_3720; // @[Bitwise.scala 50:65:@1646.4]
  wire  _T_3721; // @[Bitwise.scala 50:65:@1647.4]
  wire  _T_3722; // @[Bitwise.scala 50:65:@1648.4]
  wire  _T_3723; // @[Bitwise.scala 50:65:@1649.4]
  wire  _T_3724; // @[Bitwise.scala 50:65:@1650.4]
  wire  _T_3725; // @[Bitwise.scala 50:65:@1651.4]
  wire  _T_3726; // @[Bitwise.scala 50:65:@1652.4]
  wire [1:0] _T_3727; // @[Bitwise.scala 48:55:@1653.4]
  wire [1:0] _T_3728; // @[Bitwise.scala 48:55:@1654.4]
  wire [2:0] _T_3729; // @[Bitwise.scala 48:55:@1655.4]
  wire [1:0] _T_3730; // @[Bitwise.scala 48:55:@1656.4]
  wire [1:0] _T_3731; // @[Bitwise.scala 48:55:@1657.4]
  wire [1:0] _GEN_581; // @[Bitwise.scala 48:55:@1658.4]
  wire [2:0] _T_3732; // @[Bitwise.scala 48:55:@1658.4]
  wire [2:0] _GEN_582; // @[Bitwise.scala 48:55:@1659.4]
  wire [3:0] _T_3733; // @[Bitwise.scala 48:55:@1659.4]
  wire [3:0] _GEN_583; // @[Bitwise.scala 48:55:@1660.4]
  wire [4:0] _T_3734; // @[Bitwise.scala 48:55:@1660.4]
  wire [1:0] _T_3735; // @[Bitwise.scala 48:55:@1661.4]
  wire [1:0] _T_3736; // @[Bitwise.scala 48:55:@1662.4]
  wire [1:0] _GEN_584; // @[Bitwise.scala 48:55:@1663.4]
  wire [2:0] _T_3737; // @[Bitwise.scala 48:55:@1663.4]
  wire [2:0] _GEN_585; // @[Bitwise.scala 48:55:@1664.4]
  wire [3:0] _T_3738; // @[Bitwise.scala 48:55:@1664.4]
  wire [1:0] _T_3739; // @[Bitwise.scala 48:55:@1665.4]
  wire [1:0] _T_3740; // @[Bitwise.scala 48:55:@1666.4]
  wire [1:0] _GEN_586; // @[Bitwise.scala 48:55:@1667.4]
  wire [2:0] _T_3741; // @[Bitwise.scala 48:55:@1667.4]
  wire [2:0] _GEN_587; // @[Bitwise.scala 48:55:@1668.4]
  wire [3:0] _T_3742; // @[Bitwise.scala 48:55:@1668.4]
  wire [4:0] _T_3743; // @[Bitwise.scala 48:55:@1669.4]
  wire [5:0] _T_3744; // @[Bitwise.scala 48:55:@1670.4]
  wire [19:0] _T_3808; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1735.4]
  wire  _T_3809; // @[Bitwise.scala 50:65:@1736.4]
  wire  _T_3810; // @[Bitwise.scala 50:65:@1737.4]
  wire  _T_3811; // @[Bitwise.scala 50:65:@1738.4]
  wire  _T_3812; // @[Bitwise.scala 50:65:@1739.4]
  wire  _T_3813; // @[Bitwise.scala 50:65:@1740.4]
  wire  _T_3814; // @[Bitwise.scala 50:65:@1741.4]
  wire  _T_3815; // @[Bitwise.scala 50:65:@1742.4]
  wire  _T_3816; // @[Bitwise.scala 50:65:@1743.4]
  wire  _T_3817; // @[Bitwise.scala 50:65:@1744.4]
  wire  _T_3818; // @[Bitwise.scala 50:65:@1745.4]
  wire  _T_3819; // @[Bitwise.scala 50:65:@1746.4]
  wire  _T_3820; // @[Bitwise.scala 50:65:@1747.4]
  wire  _T_3821; // @[Bitwise.scala 50:65:@1748.4]
  wire  _T_3822; // @[Bitwise.scala 50:65:@1749.4]
  wire  _T_3823; // @[Bitwise.scala 50:65:@1750.4]
  wire  _T_3824; // @[Bitwise.scala 50:65:@1751.4]
  wire  _T_3825; // @[Bitwise.scala 50:65:@1752.4]
  wire  _T_3826; // @[Bitwise.scala 50:65:@1753.4]
  wire  _T_3827; // @[Bitwise.scala 50:65:@1754.4]
  wire  _T_3828; // @[Bitwise.scala 50:65:@1755.4]
  wire [1:0] _T_3829; // @[Bitwise.scala 48:55:@1756.4]
  wire [1:0] _T_3830; // @[Bitwise.scala 48:55:@1757.4]
  wire [1:0] _GEN_588; // @[Bitwise.scala 48:55:@1758.4]
  wire [2:0] _T_3831; // @[Bitwise.scala 48:55:@1758.4]
  wire [2:0] _GEN_589; // @[Bitwise.scala 48:55:@1759.4]
  wire [3:0] _T_3832; // @[Bitwise.scala 48:55:@1759.4]
  wire [1:0] _T_3833; // @[Bitwise.scala 48:55:@1760.4]
  wire [1:0] _T_3834; // @[Bitwise.scala 48:55:@1761.4]
  wire [1:0] _GEN_590; // @[Bitwise.scala 48:55:@1762.4]
  wire [2:0] _T_3835; // @[Bitwise.scala 48:55:@1762.4]
  wire [2:0] _GEN_591; // @[Bitwise.scala 48:55:@1763.4]
  wire [3:0] _T_3836; // @[Bitwise.scala 48:55:@1763.4]
  wire [4:0] _T_3837; // @[Bitwise.scala 48:55:@1764.4]
  wire [1:0] _T_3838; // @[Bitwise.scala 48:55:@1765.4]
  wire [1:0] _T_3839; // @[Bitwise.scala 48:55:@1766.4]
  wire [1:0] _GEN_592; // @[Bitwise.scala 48:55:@1767.4]
  wire [2:0] _T_3840; // @[Bitwise.scala 48:55:@1767.4]
  wire [2:0] _GEN_593; // @[Bitwise.scala 48:55:@1768.4]
  wire [3:0] _T_3841; // @[Bitwise.scala 48:55:@1768.4]
  wire [1:0] _T_3842; // @[Bitwise.scala 48:55:@1769.4]
  wire [1:0] _T_3843; // @[Bitwise.scala 48:55:@1770.4]
  wire [1:0] _GEN_594; // @[Bitwise.scala 48:55:@1771.4]
  wire [2:0] _T_3844; // @[Bitwise.scala 48:55:@1771.4]
  wire [2:0] _GEN_595; // @[Bitwise.scala 48:55:@1772.4]
  wire [3:0] _T_3845; // @[Bitwise.scala 48:55:@1772.4]
  wire [4:0] _T_3846; // @[Bitwise.scala 48:55:@1773.4]
  wire [5:0] _T_3847; // @[Bitwise.scala 48:55:@1774.4]
  wire [20:0] _T_3911; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1839.4]
  wire  _T_3912; // @[Bitwise.scala 50:65:@1840.4]
  wire  _T_3913; // @[Bitwise.scala 50:65:@1841.4]
  wire  _T_3914; // @[Bitwise.scala 50:65:@1842.4]
  wire  _T_3915; // @[Bitwise.scala 50:65:@1843.4]
  wire  _T_3916; // @[Bitwise.scala 50:65:@1844.4]
  wire  _T_3917; // @[Bitwise.scala 50:65:@1845.4]
  wire  _T_3918; // @[Bitwise.scala 50:65:@1846.4]
  wire  _T_3919; // @[Bitwise.scala 50:65:@1847.4]
  wire  _T_3920; // @[Bitwise.scala 50:65:@1848.4]
  wire  _T_3921; // @[Bitwise.scala 50:65:@1849.4]
  wire  _T_3922; // @[Bitwise.scala 50:65:@1850.4]
  wire  _T_3923; // @[Bitwise.scala 50:65:@1851.4]
  wire  _T_3924; // @[Bitwise.scala 50:65:@1852.4]
  wire  _T_3925; // @[Bitwise.scala 50:65:@1853.4]
  wire  _T_3926; // @[Bitwise.scala 50:65:@1854.4]
  wire  _T_3927; // @[Bitwise.scala 50:65:@1855.4]
  wire  _T_3928; // @[Bitwise.scala 50:65:@1856.4]
  wire  _T_3929; // @[Bitwise.scala 50:65:@1857.4]
  wire  _T_3930; // @[Bitwise.scala 50:65:@1858.4]
  wire  _T_3931; // @[Bitwise.scala 50:65:@1859.4]
  wire  _T_3932; // @[Bitwise.scala 50:65:@1860.4]
  wire [1:0] _T_3933; // @[Bitwise.scala 48:55:@1861.4]
  wire [1:0] _T_3934; // @[Bitwise.scala 48:55:@1862.4]
  wire [1:0] _GEN_596; // @[Bitwise.scala 48:55:@1863.4]
  wire [2:0] _T_3935; // @[Bitwise.scala 48:55:@1863.4]
  wire [2:0] _GEN_597; // @[Bitwise.scala 48:55:@1864.4]
  wire [3:0] _T_3936; // @[Bitwise.scala 48:55:@1864.4]
  wire [1:0] _T_3937; // @[Bitwise.scala 48:55:@1865.4]
  wire [1:0] _T_3938; // @[Bitwise.scala 48:55:@1866.4]
  wire [1:0] _GEN_598; // @[Bitwise.scala 48:55:@1867.4]
  wire [2:0] _T_3939; // @[Bitwise.scala 48:55:@1867.4]
  wire [2:0] _GEN_599; // @[Bitwise.scala 48:55:@1868.4]
  wire [3:0] _T_3940; // @[Bitwise.scala 48:55:@1868.4]
  wire [4:0] _T_3941; // @[Bitwise.scala 48:55:@1869.4]
  wire [1:0] _T_3942; // @[Bitwise.scala 48:55:@1870.4]
  wire [1:0] _T_3943; // @[Bitwise.scala 48:55:@1871.4]
  wire [1:0] _GEN_600; // @[Bitwise.scala 48:55:@1872.4]
  wire [2:0] _T_3944; // @[Bitwise.scala 48:55:@1872.4]
  wire [2:0] _GEN_601; // @[Bitwise.scala 48:55:@1873.4]
  wire [3:0] _T_3945; // @[Bitwise.scala 48:55:@1873.4]
  wire [1:0] _T_3946; // @[Bitwise.scala 48:55:@1874.4]
  wire [1:0] _GEN_602; // @[Bitwise.scala 48:55:@1875.4]
  wire [2:0] _T_3947; // @[Bitwise.scala 48:55:@1875.4]
  wire [1:0] _T_3948; // @[Bitwise.scala 48:55:@1876.4]
  wire [1:0] _GEN_603; // @[Bitwise.scala 48:55:@1877.4]
  wire [2:0] _T_3949; // @[Bitwise.scala 48:55:@1877.4]
  wire [3:0] _T_3950; // @[Bitwise.scala 48:55:@1878.4]
  wire [4:0] _T_3951; // @[Bitwise.scala 48:55:@1879.4]
  wire [5:0] _T_3952; // @[Bitwise.scala 48:55:@1880.4]
  wire [21:0] _T_4016; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1945.4]
  wire  _T_4017; // @[Bitwise.scala 50:65:@1946.4]
  wire  _T_4018; // @[Bitwise.scala 50:65:@1947.4]
  wire  _T_4019; // @[Bitwise.scala 50:65:@1948.4]
  wire  _T_4020; // @[Bitwise.scala 50:65:@1949.4]
  wire  _T_4021; // @[Bitwise.scala 50:65:@1950.4]
  wire  _T_4022; // @[Bitwise.scala 50:65:@1951.4]
  wire  _T_4023; // @[Bitwise.scala 50:65:@1952.4]
  wire  _T_4024; // @[Bitwise.scala 50:65:@1953.4]
  wire  _T_4025; // @[Bitwise.scala 50:65:@1954.4]
  wire  _T_4026; // @[Bitwise.scala 50:65:@1955.4]
  wire  _T_4027; // @[Bitwise.scala 50:65:@1956.4]
  wire  _T_4028; // @[Bitwise.scala 50:65:@1957.4]
  wire  _T_4029; // @[Bitwise.scala 50:65:@1958.4]
  wire  _T_4030; // @[Bitwise.scala 50:65:@1959.4]
  wire  _T_4031; // @[Bitwise.scala 50:65:@1960.4]
  wire  _T_4032; // @[Bitwise.scala 50:65:@1961.4]
  wire  _T_4033; // @[Bitwise.scala 50:65:@1962.4]
  wire  _T_4034; // @[Bitwise.scala 50:65:@1963.4]
  wire  _T_4035; // @[Bitwise.scala 50:65:@1964.4]
  wire  _T_4036; // @[Bitwise.scala 50:65:@1965.4]
  wire  _T_4037; // @[Bitwise.scala 50:65:@1966.4]
  wire  _T_4038; // @[Bitwise.scala 50:65:@1967.4]
  wire [1:0] _T_4039; // @[Bitwise.scala 48:55:@1968.4]
  wire [1:0] _T_4040; // @[Bitwise.scala 48:55:@1969.4]
  wire [1:0] _GEN_604; // @[Bitwise.scala 48:55:@1970.4]
  wire [2:0] _T_4041; // @[Bitwise.scala 48:55:@1970.4]
  wire [2:0] _GEN_605; // @[Bitwise.scala 48:55:@1971.4]
  wire [3:0] _T_4042; // @[Bitwise.scala 48:55:@1971.4]
  wire [1:0] _T_4043; // @[Bitwise.scala 48:55:@1972.4]
  wire [1:0] _GEN_606; // @[Bitwise.scala 48:55:@1973.4]
  wire [2:0] _T_4044; // @[Bitwise.scala 48:55:@1973.4]
  wire [1:0] _T_4045; // @[Bitwise.scala 48:55:@1974.4]
  wire [1:0] _GEN_607; // @[Bitwise.scala 48:55:@1975.4]
  wire [2:0] _T_4046; // @[Bitwise.scala 48:55:@1975.4]
  wire [3:0] _T_4047; // @[Bitwise.scala 48:55:@1976.4]
  wire [4:0] _T_4048; // @[Bitwise.scala 48:55:@1977.4]
  wire [1:0] _T_4049; // @[Bitwise.scala 48:55:@1978.4]
  wire [1:0] _T_4050; // @[Bitwise.scala 48:55:@1979.4]
  wire [1:0] _GEN_608; // @[Bitwise.scala 48:55:@1980.4]
  wire [2:0] _T_4051; // @[Bitwise.scala 48:55:@1980.4]
  wire [2:0] _GEN_609; // @[Bitwise.scala 48:55:@1981.4]
  wire [3:0] _T_4052; // @[Bitwise.scala 48:55:@1981.4]
  wire [1:0] _T_4053; // @[Bitwise.scala 48:55:@1982.4]
  wire [1:0] _GEN_610; // @[Bitwise.scala 48:55:@1983.4]
  wire [2:0] _T_4054; // @[Bitwise.scala 48:55:@1983.4]
  wire [1:0] _T_4055; // @[Bitwise.scala 48:55:@1984.4]
  wire [1:0] _GEN_611; // @[Bitwise.scala 48:55:@1985.4]
  wire [2:0] _T_4056; // @[Bitwise.scala 48:55:@1985.4]
  wire [3:0] _T_4057; // @[Bitwise.scala 48:55:@1986.4]
  wire [4:0] _T_4058; // @[Bitwise.scala 48:55:@1987.4]
  wire [5:0] _T_4059; // @[Bitwise.scala 48:55:@1988.4]
  wire [22:0] _T_4123; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2053.4]
  wire  _T_4124; // @[Bitwise.scala 50:65:@2054.4]
  wire  _T_4125; // @[Bitwise.scala 50:65:@2055.4]
  wire  _T_4126; // @[Bitwise.scala 50:65:@2056.4]
  wire  _T_4127; // @[Bitwise.scala 50:65:@2057.4]
  wire  _T_4128; // @[Bitwise.scala 50:65:@2058.4]
  wire  _T_4129; // @[Bitwise.scala 50:65:@2059.4]
  wire  _T_4130; // @[Bitwise.scala 50:65:@2060.4]
  wire  _T_4131; // @[Bitwise.scala 50:65:@2061.4]
  wire  _T_4132; // @[Bitwise.scala 50:65:@2062.4]
  wire  _T_4133; // @[Bitwise.scala 50:65:@2063.4]
  wire  _T_4134; // @[Bitwise.scala 50:65:@2064.4]
  wire  _T_4135; // @[Bitwise.scala 50:65:@2065.4]
  wire  _T_4136; // @[Bitwise.scala 50:65:@2066.4]
  wire  _T_4137; // @[Bitwise.scala 50:65:@2067.4]
  wire  _T_4138; // @[Bitwise.scala 50:65:@2068.4]
  wire  _T_4139; // @[Bitwise.scala 50:65:@2069.4]
  wire  _T_4140; // @[Bitwise.scala 50:65:@2070.4]
  wire  _T_4141; // @[Bitwise.scala 50:65:@2071.4]
  wire  _T_4142; // @[Bitwise.scala 50:65:@2072.4]
  wire  _T_4143; // @[Bitwise.scala 50:65:@2073.4]
  wire  _T_4144; // @[Bitwise.scala 50:65:@2074.4]
  wire  _T_4145; // @[Bitwise.scala 50:65:@2075.4]
  wire  _T_4146; // @[Bitwise.scala 50:65:@2076.4]
  wire [1:0] _T_4147; // @[Bitwise.scala 48:55:@2077.4]
  wire [1:0] _T_4148; // @[Bitwise.scala 48:55:@2078.4]
  wire [1:0] _GEN_612; // @[Bitwise.scala 48:55:@2079.4]
  wire [2:0] _T_4149; // @[Bitwise.scala 48:55:@2079.4]
  wire [2:0] _GEN_613; // @[Bitwise.scala 48:55:@2080.4]
  wire [3:0] _T_4150; // @[Bitwise.scala 48:55:@2080.4]
  wire [1:0] _T_4151; // @[Bitwise.scala 48:55:@2081.4]
  wire [1:0] _GEN_614; // @[Bitwise.scala 48:55:@2082.4]
  wire [2:0] _T_4152; // @[Bitwise.scala 48:55:@2082.4]
  wire [1:0] _T_4153; // @[Bitwise.scala 48:55:@2083.4]
  wire [1:0] _GEN_615; // @[Bitwise.scala 48:55:@2084.4]
  wire [2:0] _T_4154; // @[Bitwise.scala 48:55:@2084.4]
  wire [3:0] _T_4155; // @[Bitwise.scala 48:55:@2085.4]
  wire [4:0] _T_4156; // @[Bitwise.scala 48:55:@2086.4]
  wire [1:0] _T_4157; // @[Bitwise.scala 48:55:@2087.4]
  wire [1:0] _GEN_616; // @[Bitwise.scala 48:55:@2088.4]
  wire [2:0] _T_4158; // @[Bitwise.scala 48:55:@2088.4]
  wire [1:0] _T_4159; // @[Bitwise.scala 48:55:@2089.4]
  wire [1:0] _GEN_617; // @[Bitwise.scala 48:55:@2090.4]
  wire [2:0] _T_4160; // @[Bitwise.scala 48:55:@2090.4]
  wire [3:0] _T_4161; // @[Bitwise.scala 48:55:@2091.4]
  wire [1:0] _T_4162; // @[Bitwise.scala 48:55:@2092.4]
  wire [1:0] _GEN_618; // @[Bitwise.scala 48:55:@2093.4]
  wire [2:0] _T_4163; // @[Bitwise.scala 48:55:@2093.4]
  wire [1:0] _T_4164; // @[Bitwise.scala 48:55:@2094.4]
  wire [1:0] _GEN_619; // @[Bitwise.scala 48:55:@2095.4]
  wire [2:0] _T_4165; // @[Bitwise.scala 48:55:@2095.4]
  wire [3:0] _T_4166; // @[Bitwise.scala 48:55:@2096.4]
  wire [4:0] _T_4167; // @[Bitwise.scala 48:55:@2097.4]
  wire [5:0] _T_4168; // @[Bitwise.scala 48:55:@2098.4]
  wire [23:0] _T_4232; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2163.4]
  wire  _T_4233; // @[Bitwise.scala 50:65:@2164.4]
  wire  _T_4234; // @[Bitwise.scala 50:65:@2165.4]
  wire  _T_4235; // @[Bitwise.scala 50:65:@2166.4]
  wire  _T_4236; // @[Bitwise.scala 50:65:@2167.4]
  wire  _T_4237; // @[Bitwise.scala 50:65:@2168.4]
  wire  _T_4238; // @[Bitwise.scala 50:65:@2169.4]
  wire  _T_4239; // @[Bitwise.scala 50:65:@2170.4]
  wire  _T_4240; // @[Bitwise.scala 50:65:@2171.4]
  wire  _T_4241; // @[Bitwise.scala 50:65:@2172.4]
  wire  _T_4242; // @[Bitwise.scala 50:65:@2173.4]
  wire  _T_4243; // @[Bitwise.scala 50:65:@2174.4]
  wire  _T_4244; // @[Bitwise.scala 50:65:@2175.4]
  wire  _T_4245; // @[Bitwise.scala 50:65:@2176.4]
  wire  _T_4246; // @[Bitwise.scala 50:65:@2177.4]
  wire  _T_4247; // @[Bitwise.scala 50:65:@2178.4]
  wire  _T_4248; // @[Bitwise.scala 50:65:@2179.4]
  wire  _T_4249; // @[Bitwise.scala 50:65:@2180.4]
  wire  _T_4250; // @[Bitwise.scala 50:65:@2181.4]
  wire  _T_4251; // @[Bitwise.scala 50:65:@2182.4]
  wire  _T_4252; // @[Bitwise.scala 50:65:@2183.4]
  wire  _T_4253; // @[Bitwise.scala 50:65:@2184.4]
  wire  _T_4254; // @[Bitwise.scala 50:65:@2185.4]
  wire  _T_4255; // @[Bitwise.scala 50:65:@2186.4]
  wire  _T_4256; // @[Bitwise.scala 50:65:@2187.4]
  wire [1:0] _T_4257; // @[Bitwise.scala 48:55:@2188.4]
  wire [1:0] _GEN_620; // @[Bitwise.scala 48:55:@2189.4]
  wire [2:0] _T_4258; // @[Bitwise.scala 48:55:@2189.4]
  wire [1:0] _T_4259; // @[Bitwise.scala 48:55:@2190.4]
  wire [1:0] _GEN_621; // @[Bitwise.scala 48:55:@2191.4]
  wire [2:0] _T_4260; // @[Bitwise.scala 48:55:@2191.4]
  wire [3:0] _T_4261; // @[Bitwise.scala 48:55:@2192.4]
  wire [1:0] _T_4262; // @[Bitwise.scala 48:55:@2193.4]
  wire [1:0] _GEN_622; // @[Bitwise.scala 48:55:@2194.4]
  wire [2:0] _T_4263; // @[Bitwise.scala 48:55:@2194.4]
  wire [1:0] _T_4264; // @[Bitwise.scala 48:55:@2195.4]
  wire [1:0] _GEN_623; // @[Bitwise.scala 48:55:@2196.4]
  wire [2:0] _T_4265; // @[Bitwise.scala 48:55:@2196.4]
  wire [3:0] _T_4266; // @[Bitwise.scala 48:55:@2197.4]
  wire [4:0] _T_4267; // @[Bitwise.scala 48:55:@2198.4]
  wire [1:0] _T_4268; // @[Bitwise.scala 48:55:@2199.4]
  wire [1:0] _GEN_624; // @[Bitwise.scala 48:55:@2200.4]
  wire [2:0] _T_4269; // @[Bitwise.scala 48:55:@2200.4]
  wire [1:0] _T_4270; // @[Bitwise.scala 48:55:@2201.4]
  wire [1:0] _GEN_625; // @[Bitwise.scala 48:55:@2202.4]
  wire [2:0] _T_4271; // @[Bitwise.scala 48:55:@2202.4]
  wire [3:0] _T_4272; // @[Bitwise.scala 48:55:@2203.4]
  wire [1:0] _T_4273; // @[Bitwise.scala 48:55:@2204.4]
  wire [1:0] _GEN_626; // @[Bitwise.scala 48:55:@2205.4]
  wire [2:0] _T_4274; // @[Bitwise.scala 48:55:@2205.4]
  wire [1:0] _T_4275; // @[Bitwise.scala 48:55:@2206.4]
  wire [1:0] _GEN_627; // @[Bitwise.scala 48:55:@2207.4]
  wire [2:0] _T_4276; // @[Bitwise.scala 48:55:@2207.4]
  wire [3:0] _T_4277; // @[Bitwise.scala 48:55:@2208.4]
  wire [4:0] _T_4278; // @[Bitwise.scala 48:55:@2209.4]
  wire [5:0] _T_4279; // @[Bitwise.scala 48:55:@2210.4]
  wire [24:0] _T_4343; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2275.4]
  wire  _T_4344; // @[Bitwise.scala 50:65:@2276.4]
  wire  _T_4345; // @[Bitwise.scala 50:65:@2277.4]
  wire  _T_4346; // @[Bitwise.scala 50:65:@2278.4]
  wire  _T_4347; // @[Bitwise.scala 50:65:@2279.4]
  wire  _T_4348; // @[Bitwise.scala 50:65:@2280.4]
  wire  _T_4349; // @[Bitwise.scala 50:65:@2281.4]
  wire  _T_4350; // @[Bitwise.scala 50:65:@2282.4]
  wire  _T_4351; // @[Bitwise.scala 50:65:@2283.4]
  wire  _T_4352; // @[Bitwise.scala 50:65:@2284.4]
  wire  _T_4353; // @[Bitwise.scala 50:65:@2285.4]
  wire  _T_4354; // @[Bitwise.scala 50:65:@2286.4]
  wire  _T_4355; // @[Bitwise.scala 50:65:@2287.4]
  wire  _T_4356; // @[Bitwise.scala 50:65:@2288.4]
  wire  _T_4357; // @[Bitwise.scala 50:65:@2289.4]
  wire  _T_4358; // @[Bitwise.scala 50:65:@2290.4]
  wire  _T_4359; // @[Bitwise.scala 50:65:@2291.4]
  wire  _T_4360; // @[Bitwise.scala 50:65:@2292.4]
  wire  _T_4361; // @[Bitwise.scala 50:65:@2293.4]
  wire  _T_4362; // @[Bitwise.scala 50:65:@2294.4]
  wire  _T_4363; // @[Bitwise.scala 50:65:@2295.4]
  wire  _T_4364; // @[Bitwise.scala 50:65:@2296.4]
  wire  _T_4365; // @[Bitwise.scala 50:65:@2297.4]
  wire  _T_4366; // @[Bitwise.scala 50:65:@2298.4]
  wire  _T_4367; // @[Bitwise.scala 50:65:@2299.4]
  wire  _T_4368; // @[Bitwise.scala 50:65:@2300.4]
  wire [1:0] _T_4369; // @[Bitwise.scala 48:55:@2301.4]
  wire [1:0] _GEN_628; // @[Bitwise.scala 48:55:@2302.4]
  wire [2:0] _T_4370; // @[Bitwise.scala 48:55:@2302.4]
  wire [1:0] _T_4371; // @[Bitwise.scala 48:55:@2303.4]
  wire [1:0] _GEN_629; // @[Bitwise.scala 48:55:@2304.4]
  wire [2:0] _T_4372; // @[Bitwise.scala 48:55:@2304.4]
  wire [3:0] _T_4373; // @[Bitwise.scala 48:55:@2305.4]
  wire [1:0] _T_4374; // @[Bitwise.scala 48:55:@2306.4]
  wire [1:0] _GEN_630; // @[Bitwise.scala 48:55:@2307.4]
  wire [2:0] _T_4375; // @[Bitwise.scala 48:55:@2307.4]
  wire [1:0] _T_4376; // @[Bitwise.scala 48:55:@2308.4]
  wire [1:0] _GEN_631; // @[Bitwise.scala 48:55:@2309.4]
  wire [2:0] _T_4377; // @[Bitwise.scala 48:55:@2309.4]
  wire [3:0] _T_4378; // @[Bitwise.scala 48:55:@2310.4]
  wire [4:0] _T_4379; // @[Bitwise.scala 48:55:@2311.4]
  wire [1:0] _T_4380; // @[Bitwise.scala 48:55:@2312.4]
  wire [1:0] _GEN_632; // @[Bitwise.scala 48:55:@2313.4]
  wire [2:0] _T_4381; // @[Bitwise.scala 48:55:@2313.4]
  wire [1:0] _T_4382; // @[Bitwise.scala 48:55:@2314.4]
  wire [1:0] _GEN_633; // @[Bitwise.scala 48:55:@2315.4]
  wire [2:0] _T_4383; // @[Bitwise.scala 48:55:@2315.4]
  wire [3:0] _T_4384; // @[Bitwise.scala 48:55:@2316.4]
  wire [1:0] _T_4385; // @[Bitwise.scala 48:55:@2317.4]
  wire [1:0] _GEN_634; // @[Bitwise.scala 48:55:@2318.4]
  wire [2:0] _T_4386; // @[Bitwise.scala 48:55:@2318.4]
  wire [1:0] _T_4387; // @[Bitwise.scala 48:55:@2319.4]
  wire [1:0] _T_4388; // @[Bitwise.scala 48:55:@2320.4]
  wire [2:0] _T_4389; // @[Bitwise.scala 48:55:@2321.4]
  wire [3:0] _T_4390; // @[Bitwise.scala 48:55:@2322.4]
  wire [4:0] _T_4391; // @[Bitwise.scala 48:55:@2323.4]
  wire [5:0] _T_4392; // @[Bitwise.scala 48:55:@2324.4]
  wire [25:0] _T_4456; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2389.4]
  wire  _T_4457; // @[Bitwise.scala 50:65:@2390.4]
  wire  _T_4458; // @[Bitwise.scala 50:65:@2391.4]
  wire  _T_4459; // @[Bitwise.scala 50:65:@2392.4]
  wire  _T_4460; // @[Bitwise.scala 50:65:@2393.4]
  wire  _T_4461; // @[Bitwise.scala 50:65:@2394.4]
  wire  _T_4462; // @[Bitwise.scala 50:65:@2395.4]
  wire  _T_4463; // @[Bitwise.scala 50:65:@2396.4]
  wire  _T_4464; // @[Bitwise.scala 50:65:@2397.4]
  wire  _T_4465; // @[Bitwise.scala 50:65:@2398.4]
  wire  _T_4466; // @[Bitwise.scala 50:65:@2399.4]
  wire  _T_4467; // @[Bitwise.scala 50:65:@2400.4]
  wire  _T_4468; // @[Bitwise.scala 50:65:@2401.4]
  wire  _T_4469; // @[Bitwise.scala 50:65:@2402.4]
  wire  _T_4470; // @[Bitwise.scala 50:65:@2403.4]
  wire  _T_4471; // @[Bitwise.scala 50:65:@2404.4]
  wire  _T_4472; // @[Bitwise.scala 50:65:@2405.4]
  wire  _T_4473; // @[Bitwise.scala 50:65:@2406.4]
  wire  _T_4474; // @[Bitwise.scala 50:65:@2407.4]
  wire  _T_4475; // @[Bitwise.scala 50:65:@2408.4]
  wire  _T_4476; // @[Bitwise.scala 50:65:@2409.4]
  wire  _T_4477; // @[Bitwise.scala 50:65:@2410.4]
  wire  _T_4478; // @[Bitwise.scala 50:65:@2411.4]
  wire  _T_4479; // @[Bitwise.scala 50:65:@2412.4]
  wire  _T_4480; // @[Bitwise.scala 50:65:@2413.4]
  wire  _T_4481; // @[Bitwise.scala 50:65:@2414.4]
  wire  _T_4482; // @[Bitwise.scala 50:65:@2415.4]
  wire [1:0] _T_4483; // @[Bitwise.scala 48:55:@2416.4]
  wire [1:0] _GEN_635; // @[Bitwise.scala 48:55:@2417.4]
  wire [2:0] _T_4484; // @[Bitwise.scala 48:55:@2417.4]
  wire [1:0] _T_4485; // @[Bitwise.scala 48:55:@2418.4]
  wire [1:0] _GEN_636; // @[Bitwise.scala 48:55:@2419.4]
  wire [2:0] _T_4486; // @[Bitwise.scala 48:55:@2419.4]
  wire [3:0] _T_4487; // @[Bitwise.scala 48:55:@2420.4]
  wire [1:0] _T_4488; // @[Bitwise.scala 48:55:@2421.4]
  wire [1:0] _GEN_637; // @[Bitwise.scala 48:55:@2422.4]
  wire [2:0] _T_4489; // @[Bitwise.scala 48:55:@2422.4]
  wire [1:0] _T_4490; // @[Bitwise.scala 48:55:@2423.4]
  wire [1:0] _T_4491; // @[Bitwise.scala 48:55:@2424.4]
  wire [2:0] _T_4492; // @[Bitwise.scala 48:55:@2425.4]
  wire [3:0] _T_4493; // @[Bitwise.scala 48:55:@2426.4]
  wire [4:0] _T_4494; // @[Bitwise.scala 48:55:@2427.4]
  wire [1:0] _T_4495; // @[Bitwise.scala 48:55:@2428.4]
  wire [1:0] _GEN_638; // @[Bitwise.scala 48:55:@2429.4]
  wire [2:0] _T_4496; // @[Bitwise.scala 48:55:@2429.4]
  wire [1:0] _T_4497; // @[Bitwise.scala 48:55:@2430.4]
  wire [1:0] _GEN_639; // @[Bitwise.scala 48:55:@2431.4]
  wire [2:0] _T_4498; // @[Bitwise.scala 48:55:@2431.4]
  wire [3:0] _T_4499; // @[Bitwise.scala 48:55:@2432.4]
  wire [1:0] _T_4500; // @[Bitwise.scala 48:55:@2433.4]
  wire [1:0] _GEN_640; // @[Bitwise.scala 48:55:@2434.4]
  wire [2:0] _T_4501; // @[Bitwise.scala 48:55:@2434.4]
  wire [1:0] _T_4502; // @[Bitwise.scala 48:55:@2435.4]
  wire [1:0] _T_4503; // @[Bitwise.scala 48:55:@2436.4]
  wire [2:0] _T_4504; // @[Bitwise.scala 48:55:@2437.4]
  wire [3:0] _T_4505; // @[Bitwise.scala 48:55:@2438.4]
  wire [4:0] _T_4506; // @[Bitwise.scala 48:55:@2439.4]
  wire [5:0] _T_4507; // @[Bitwise.scala 48:55:@2440.4]
  wire [26:0] _T_4571; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2505.4]
  wire  _T_4572; // @[Bitwise.scala 50:65:@2506.4]
  wire  _T_4573; // @[Bitwise.scala 50:65:@2507.4]
  wire  _T_4574; // @[Bitwise.scala 50:65:@2508.4]
  wire  _T_4575; // @[Bitwise.scala 50:65:@2509.4]
  wire  _T_4576; // @[Bitwise.scala 50:65:@2510.4]
  wire  _T_4577; // @[Bitwise.scala 50:65:@2511.4]
  wire  _T_4578; // @[Bitwise.scala 50:65:@2512.4]
  wire  _T_4579; // @[Bitwise.scala 50:65:@2513.4]
  wire  _T_4580; // @[Bitwise.scala 50:65:@2514.4]
  wire  _T_4581; // @[Bitwise.scala 50:65:@2515.4]
  wire  _T_4582; // @[Bitwise.scala 50:65:@2516.4]
  wire  _T_4583; // @[Bitwise.scala 50:65:@2517.4]
  wire  _T_4584; // @[Bitwise.scala 50:65:@2518.4]
  wire  _T_4585; // @[Bitwise.scala 50:65:@2519.4]
  wire  _T_4586; // @[Bitwise.scala 50:65:@2520.4]
  wire  _T_4587; // @[Bitwise.scala 50:65:@2521.4]
  wire  _T_4588; // @[Bitwise.scala 50:65:@2522.4]
  wire  _T_4589; // @[Bitwise.scala 50:65:@2523.4]
  wire  _T_4590; // @[Bitwise.scala 50:65:@2524.4]
  wire  _T_4591; // @[Bitwise.scala 50:65:@2525.4]
  wire  _T_4592; // @[Bitwise.scala 50:65:@2526.4]
  wire  _T_4593; // @[Bitwise.scala 50:65:@2527.4]
  wire  _T_4594; // @[Bitwise.scala 50:65:@2528.4]
  wire  _T_4595; // @[Bitwise.scala 50:65:@2529.4]
  wire  _T_4596; // @[Bitwise.scala 50:65:@2530.4]
  wire  _T_4597; // @[Bitwise.scala 50:65:@2531.4]
  wire  _T_4598; // @[Bitwise.scala 50:65:@2532.4]
  wire [1:0] _T_4599; // @[Bitwise.scala 48:55:@2533.4]
  wire [1:0] _GEN_641; // @[Bitwise.scala 48:55:@2534.4]
  wire [2:0] _T_4600; // @[Bitwise.scala 48:55:@2534.4]
  wire [1:0] _T_4601; // @[Bitwise.scala 48:55:@2535.4]
  wire [1:0] _GEN_642; // @[Bitwise.scala 48:55:@2536.4]
  wire [2:0] _T_4602; // @[Bitwise.scala 48:55:@2536.4]
  wire [3:0] _T_4603; // @[Bitwise.scala 48:55:@2537.4]
  wire [1:0] _T_4604; // @[Bitwise.scala 48:55:@2538.4]
  wire [1:0] _GEN_643; // @[Bitwise.scala 48:55:@2539.4]
  wire [2:0] _T_4605; // @[Bitwise.scala 48:55:@2539.4]
  wire [1:0] _T_4606; // @[Bitwise.scala 48:55:@2540.4]
  wire [1:0] _T_4607; // @[Bitwise.scala 48:55:@2541.4]
  wire [2:0] _T_4608; // @[Bitwise.scala 48:55:@2542.4]
  wire [3:0] _T_4609; // @[Bitwise.scala 48:55:@2543.4]
  wire [4:0] _T_4610; // @[Bitwise.scala 48:55:@2544.4]
  wire [1:0] _T_4611; // @[Bitwise.scala 48:55:@2545.4]
  wire [1:0] _GEN_644; // @[Bitwise.scala 48:55:@2546.4]
  wire [2:0] _T_4612; // @[Bitwise.scala 48:55:@2546.4]
  wire [1:0] _T_4613; // @[Bitwise.scala 48:55:@2547.4]
  wire [1:0] _T_4614; // @[Bitwise.scala 48:55:@2548.4]
  wire [2:0] _T_4615; // @[Bitwise.scala 48:55:@2549.4]
  wire [3:0] _T_4616; // @[Bitwise.scala 48:55:@2550.4]
  wire [1:0] _T_4617; // @[Bitwise.scala 48:55:@2551.4]
  wire [1:0] _GEN_645; // @[Bitwise.scala 48:55:@2552.4]
  wire [2:0] _T_4618; // @[Bitwise.scala 48:55:@2552.4]
  wire [1:0] _T_4619; // @[Bitwise.scala 48:55:@2553.4]
  wire [1:0] _T_4620; // @[Bitwise.scala 48:55:@2554.4]
  wire [2:0] _T_4621; // @[Bitwise.scala 48:55:@2555.4]
  wire [3:0] _T_4622; // @[Bitwise.scala 48:55:@2556.4]
  wire [4:0] _T_4623; // @[Bitwise.scala 48:55:@2557.4]
  wire [5:0] _T_4624; // @[Bitwise.scala 48:55:@2558.4]
  wire [27:0] _T_4688; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2623.4]
  wire  _T_4689; // @[Bitwise.scala 50:65:@2624.4]
  wire  _T_4690; // @[Bitwise.scala 50:65:@2625.4]
  wire  _T_4691; // @[Bitwise.scala 50:65:@2626.4]
  wire  _T_4692; // @[Bitwise.scala 50:65:@2627.4]
  wire  _T_4693; // @[Bitwise.scala 50:65:@2628.4]
  wire  _T_4694; // @[Bitwise.scala 50:65:@2629.4]
  wire  _T_4695; // @[Bitwise.scala 50:65:@2630.4]
  wire  _T_4696; // @[Bitwise.scala 50:65:@2631.4]
  wire  _T_4697; // @[Bitwise.scala 50:65:@2632.4]
  wire  _T_4698; // @[Bitwise.scala 50:65:@2633.4]
  wire  _T_4699; // @[Bitwise.scala 50:65:@2634.4]
  wire  _T_4700; // @[Bitwise.scala 50:65:@2635.4]
  wire  _T_4701; // @[Bitwise.scala 50:65:@2636.4]
  wire  _T_4702; // @[Bitwise.scala 50:65:@2637.4]
  wire  _T_4703; // @[Bitwise.scala 50:65:@2638.4]
  wire  _T_4704; // @[Bitwise.scala 50:65:@2639.4]
  wire  _T_4705; // @[Bitwise.scala 50:65:@2640.4]
  wire  _T_4706; // @[Bitwise.scala 50:65:@2641.4]
  wire  _T_4707; // @[Bitwise.scala 50:65:@2642.4]
  wire  _T_4708; // @[Bitwise.scala 50:65:@2643.4]
  wire  _T_4709; // @[Bitwise.scala 50:65:@2644.4]
  wire  _T_4710; // @[Bitwise.scala 50:65:@2645.4]
  wire  _T_4711; // @[Bitwise.scala 50:65:@2646.4]
  wire  _T_4712; // @[Bitwise.scala 50:65:@2647.4]
  wire  _T_4713; // @[Bitwise.scala 50:65:@2648.4]
  wire  _T_4714; // @[Bitwise.scala 50:65:@2649.4]
  wire  _T_4715; // @[Bitwise.scala 50:65:@2650.4]
  wire  _T_4716; // @[Bitwise.scala 50:65:@2651.4]
  wire [1:0] _T_4717; // @[Bitwise.scala 48:55:@2652.4]
  wire [1:0] _GEN_646; // @[Bitwise.scala 48:55:@2653.4]
  wire [2:0] _T_4718; // @[Bitwise.scala 48:55:@2653.4]
  wire [1:0] _T_4719; // @[Bitwise.scala 48:55:@2654.4]
  wire [1:0] _T_4720; // @[Bitwise.scala 48:55:@2655.4]
  wire [2:0] _T_4721; // @[Bitwise.scala 48:55:@2656.4]
  wire [3:0] _T_4722; // @[Bitwise.scala 48:55:@2657.4]
  wire [1:0] _T_4723; // @[Bitwise.scala 48:55:@2658.4]
  wire [1:0] _GEN_647; // @[Bitwise.scala 48:55:@2659.4]
  wire [2:0] _T_4724; // @[Bitwise.scala 48:55:@2659.4]
  wire [1:0] _T_4725; // @[Bitwise.scala 48:55:@2660.4]
  wire [1:0] _T_4726; // @[Bitwise.scala 48:55:@2661.4]
  wire [2:0] _T_4727; // @[Bitwise.scala 48:55:@2662.4]
  wire [3:0] _T_4728; // @[Bitwise.scala 48:55:@2663.4]
  wire [4:0] _T_4729; // @[Bitwise.scala 48:55:@2664.4]
  wire [1:0] _T_4730; // @[Bitwise.scala 48:55:@2665.4]
  wire [1:0] _GEN_648; // @[Bitwise.scala 48:55:@2666.4]
  wire [2:0] _T_4731; // @[Bitwise.scala 48:55:@2666.4]
  wire [1:0] _T_4732; // @[Bitwise.scala 48:55:@2667.4]
  wire [1:0] _T_4733; // @[Bitwise.scala 48:55:@2668.4]
  wire [2:0] _T_4734; // @[Bitwise.scala 48:55:@2669.4]
  wire [3:0] _T_4735; // @[Bitwise.scala 48:55:@2670.4]
  wire [1:0] _T_4736; // @[Bitwise.scala 48:55:@2671.4]
  wire [1:0] _GEN_649; // @[Bitwise.scala 48:55:@2672.4]
  wire [2:0] _T_4737; // @[Bitwise.scala 48:55:@2672.4]
  wire [1:0] _T_4738; // @[Bitwise.scala 48:55:@2673.4]
  wire [1:0] _T_4739; // @[Bitwise.scala 48:55:@2674.4]
  wire [2:0] _T_4740; // @[Bitwise.scala 48:55:@2675.4]
  wire [3:0] _T_4741; // @[Bitwise.scala 48:55:@2676.4]
  wire [4:0] _T_4742; // @[Bitwise.scala 48:55:@2677.4]
  wire [5:0] _T_4743; // @[Bitwise.scala 48:55:@2678.4]
  wire [28:0] _T_4807; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2743.4]
  wire  _T_4808; // @[Bitwise.scala 50:65:@2744.4]
  wire  _T_4809; // @[Bitwise.scala 50:65:@2745.4]
  wire  _T_4810; // @[Bitwise.scala 50:65:@2746.4]
  wire  _T_4811; // @[Bitwise.scala 50:65:@2747.4]
  wire  _T_4812; // @[Bitwise.scala 50:65:@2748.4]
  wire  _T_4813; // @[Bitwise.scala 50:65:@2749.4]
  wire  _T_4814; // @[Bitwise.scala 50:65:@2750.4]
  wire  _T_4815; // @[Bitwise.scala 50:65:@2751.4]
  wire  _T_4816; // @[Bitwise.scala 50:65:@2752.4]
  wire  _T_4817; // @[Bitwise.scala 50:65:@2753.4]
  wire  _T_4818; // @[Bitwise.scala 50:65:@2754.4]
  wire  _T_4819; // @[Bitwise.scala 50:65:@2755.4]
  wire  _T_4820; // @[Bitwise.scala 50:65:@2756.4]
  wire  _T_4821; // @[Bitwise.scala 50:65:@2757.4]
  wire  _T_4822; // @[Bitwise.scala 50:65:@2758.4]
  wire  _T_4823; // @[Bitwise.scala 50:65:@2759.4]
  wire  _T_4824; // @[Bitwise.scala 50:65:@2760.4]
  wire  _T_4825; // @[Bitwise.scala 50:65:@2761.4]
  wire  _T_4826; // @[Bitwise.scala 50:65:@2762.4]
  wire  _T_4827; // @[Bitwise.scala 50:65:@2763.4]
  wire  _T_4828; // @[Bitwise.scala 50:65:@2764.4]
  wire  _T_4829; // @[Bitwise.scala 50:65:@2765.4]
  wire  _T_4830; // @[Bitwise.scala 50:65:@2766.4]
  wire  _T_4831; // @[Bitwise.scala 50:65:@2767.4]
  wire  _T_4832; // @[Bitwise.scala 50:65:@2768.4]
  wire  _T_4833; // @[Bitwise.scala 50:65:@2769.4]
  wire  _T_4834; // @[Bitwise.scala 50:65:@2770.4]
  wire  _T_4835; // @[Bitwise.scala 50:65:@2771.4]
  wire  _T_4836; // @[Bitwise.scala 50:65:@2772.4]
  wire [1:0] _T_4837; // @[Bitwise.scala 48:55:@2773.4]
  wire [1:0] _GEN_650; // @[Bitwise.scala 48:55:@2774.4]
  wire [2:0] _T_4838; // @[Bitwise.scala 48:55:@2774.4]
  wire [1:0] _T_4839; // @[Bitwise.scala 48:55:@2775.4]
  wire [1:0] _T_4840; // @[Bitwise.scala 48:55:@2776.4]
  wire [2:0] _T_4841; // @[Bitwise.scala 48:55:@2777.4]
  wire [3:0] _T_4842; // @[Bitwise.scala 48:55:@2778.4]
  wire [1:0] _T_4843; // @[Bitwise.scala 48:55:@2779.4]
  wire [1:0] _GEN_651; // @[Bitwise.scala 48:55:@2780.4]
  wire [2:0] _T_4844; // @[Bitwise.scala 48:55:@2780.4]
  wire [1:0] _T_4845; // @[Bitwise.scala 48:55:@2781.4]
  wire [1:0] _T_4846; // @[Bitwise.scala 48:55:@2782.4]
  wire [2:0] _T_4847; // @[Bitwise.scala 48:55:@2783.4]
  wire [3:0] _T_4848; // @[Bitwise.scala 48:55:@2784.4]
  wire [4:0] _T_4849; // @[Bitwise.scala 48:55:@2785.4]
  wire [1:0] _T_4850; // @[Bitwise.scala 48:55:@2786.4]
  wire [1:0] _GEN_652; // @[Bitwise.scala 48:55:@2787.4]
  wire [2:0] _T_4851; // @[Bitwise.scala 48:55:@2787.4]
  wire [1:0] _T_4852; // @[Bitwise.scala 48:55:@2788.4]
  wire [1:0] _T_4853; // @[Bitwise.scala 48:55:@2789.4]
  wire [2:0] _T_4854; // @[Bitwise.scala 48:55:@2790.4]
  wire [3:0] _T_4855; // @[Bitwise.scala 48:55:@2791.4]
  wire [1:0] _T_4856; // @[Bitwise.scala 48:55:@2792.4]
  wire [1:0] _T_4857; // @[Bitwise.scala 48:55:@2793.4]
  wire [2:0] _T_4858; // @[Bitwise.scala 48:55:@2794.4]
  wire [1:0] _T_4859; // @[Bitwise.scala 48:55:@2795.4]
  wire [1:0] _T_4860; // @[Bitwise.scala 48:55:@2796.4]
  wire [2:0] _T_4861; // @[Bitwise.scala 48:55:@2797.4]
  wire [3:0] _T_4862; // @[Bitwise.scala 48:55:@2798.4]
  wire [4:0] _T_4863; // @[Bitwise.scala 48:55:@2799.4]
  wire [5:0] _T_4864; // @[Bitwise.scala 48:55:@2800.4]
  wire [29:0] _T_4928; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2865.4]
  wire  _T_4929; // @[Bitwise.scala 50:65:@2866.4]
  wire  _T_4930; // @[Bitwise.scala 50:65:@2867.4]
  wire  _T_4931; // @[Bitwise.scala 50:65:@2868.4]
  wire  _T_4932; // @[Bitwise.scala 50:65:@2869.4]
  wire  _T_4933; // @[Bitwise.scala 50:65:@2870.4]
  wire  _T_4934; // @[Bitwise.scala 50:65:@2871.4]
  wire  _T_4935; // @[Bitwise.scala 50:65:@2872.4]
  wire  _T_4936; // @[Bitwise.scala 50:65:@2873.4]
  wire  _T_4937; // @[Bitwise.scala 50:65:@2874.4]
  wire  _T_4938; // @[Bitwise.scala 50:65:@2875.4]
  wire  _T_4939; // @[Bitwise.scala 50:65:@2876.4]
  wire  _T_4940; // @[Bitwise.scala 50:65:@2877.4]
  wire  _T_4941; // @[Bitwise.scala 50:65:@2878.4]
  wire  _T_4942; // @[Bitwise.scala 50:65:@2879.4]
  wire  _T_4943; // @[Bitwise.scala 50:65:@2880.4]
  wire  _T_4944; // @[Bitwise.scala 50:65:@2881.4]
  wire  _T_4945; // @[Bitwise.scala 50:65:@2882.4]
  wire  _T_4946; // @[Bitwise.scala 50:65:@2883.4]
  wire  _T_4947; // @[Bitwise.scala 50:65:@2884.4]
  wire  _T_4948; // @[Bitwise.scala 50:65:@2885.4]
  wire  _T_4949; // @[Bitwise.scala 50:65:@2886.4]
  wire  _T_4950; // @[Bitwise.scala 50:65:@2887.4]
  wire  _T_4951; // @[Bitwise.scala 50:65:@2888.4]
  wire  _T_4952; // @[Bitwise.scala 50:65:@2889.4]
  wire  _T_4953; // @[Bitwise.scala 50:65:@2890.4]
  wire  _T_4954; // @[Bitwise.scala 50:65:@2891.4]
  wire  _T_4955; // @[Bitwise.scala 50:65:@2892.4]
  wire  _T_4956; // @[Bitwise.scala 50:65:@2893.4]
  wire  _T_4957; // @[Bitwise.scala 50:65:@2894.4]
  wire  _T_4958; // @[Bitwise.scala 50:65:@2895.4]
  wire [1:0] _T_4959; // @[Bitwise.scala 48:55:@2896.4]
  wire [1:0] _GEN_653; // @[Bitwise.scala 48:55:@2897.4]
  wire [2:0] _T_4960; // @[Bitwise.scala 48:55:@2897.4]
  wire [1:0] _T_4961; // @[Bitwise.scala 48:55:@2898.4]
  wire [1:0] _T_4962; // @[Bitwise.scala 48:55:@2899.4]
  wire [2:0] _T_4963; // @[Bitwise.scala 48:55:@2900.4]
  wire [3:0] _T_4964; // @[Bitwise.scala 48:55:@2901.4]
  wire [1:0] _T_4965; // @[Bitwise.scala 48:55:@2902.4]
  wire [1:0] _T_4966; // @[Bitwise.scala 48:55:@2903.4]
  wire [2:0] _T_4967; // @[Bitwise.scala 48:55:@2904.4]
  wire [1:0] _T_4968; // @[Bitwise.scala 48:55:@2905.4]
  wire [1:0] _T_4969; // @[Bitwise.scala 48:55:@2906.4]
  wire [2:0] _T_4970; // @[Bitwise.scala 48:55:@2907.4]
  wire [3:0] _T_4971; // @[Bitwise.scala 48:55:@2908.4]
  wire [4:0] _T_4972; // @[Bitwise.scala 48:55:@2909.4]
  wire [1:0] _T_4973; // @[Bitwise.scala 48:55:@2910.4]
  wire [1:0] _GEN_654; // @[Bitwise.scala 48:55:@2911.4]
  wire [2:0] _T_4974; // @[Bitwise.scala 48:55:@2911.4]
  wire [1:0] _T_4975; // @[Bitwise.scala 48:55:@2912.4]
  wire [1:0] _T_4976; // @[Bitwise.scala 48:55:@2913.4]
  wire [2:0] _T_4977; // @[Bitwise.scala 48:55:@2914.4]
  wire [3:0] _T_4978; // @[Bitwise.scala 48:55:@2915.4]
  wire [1:0] _T_4979; // @[Bitwise.scala 48:55:@2916.4]
  wire [1:0] _T_4980; // @[Bitwise.scala 48:55:@2917.4]
  wire [2:0] _T_4981; // @[Bitwise.scala 48:55:@2918.4]
  wire [1:0] _T_4982; // @[Bitwise.scala 48:55:@2919.4]
  wire [1:0] _T_4983; // @[Bitwise.scala 48:55:@2920.4]
  wire [2:0] _T_4984; // @[Bitwise.scala 48:55:@2921.4]
  wire [3:0] _T_4985; // @[Bitwise.scala 48:55:@2922.4]
  wire [4:0] _T_4986; // @[Bitwise.scala 48:55:@2923.4]
  wire [5:0] _T_4987; // @[Bitwise.scala 48:55:@2924.4]
  wire [30:0] _T_5051; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2989.4]
  wire  _T_5052; // @[Bitwise.scala 50:65:@2990.4]
  wire  _T_5053; // @[Bitwise.scala 50:65:@2991.4]
  wire  _T_5054; // @[Bitwise.scala 50:65:@2992.4]
  wire  _T_5055; // @[Bitwise.scala 50:65:@2993.4]
  wire  _T_5056; // @[Bitwise.scala 50:65:@2994.4]
  wire  _T_5057; // @[Bitwise.scala 50:65:@2995.4]
  wire  _T_5058; // @[Bitwise.scala 50:65:@2996.4]
  wire  _T_5059; // @[Bitwise.scala 50:65:@2997.4]
  wire  _T_5060; // @[Bitwise.scala 50:65:@2998.4]
  wire  _T_5061; // @[Bitwise.scala 50:65:@2999.4]
  wire  _T_5062; // @[Bitwise.scala 50:65:@3000.4]
  wire  _T_5063; // @[Bitwise.scala 50:65:@3001.4]
  wire  _T_5064; // @[Bitwise.scala 50:65:@3002.4]
  wire  _T_5065; // @[Bitwise.scala 50:65:@3003.4]
  wire  _T_5066; // @[Bitwise.scala 50:65:@3004.4]
  wire  _T_5067; // @[Bitwise.scala 50:65:@3005.4]
  wire  _T_5068; // @[Bitwise.scala 50:65:@3006.4]
  wire  _T_5069; // @[Bitwise.scala 50:65:@3007.4]
  wire  _T_5070; // @[Bitwise.scala 50:65:@3008.4]
  wire  _T_5071; // @[Bitwise.scala 50:65:@3009.4]
  wire  _T_5072; // @[Bitwise.scala 50:65:@3010.4]
  wire  _T_5073; // @[Bitwise.scala 50:65:@3011.4]
  wire  _T_5074; // @[Bitwise.scala 50:65:@3012.4]
  wire  _T_5075; // @[Bitwise.scala 50:65:@3013.4]
  wire  _T_5076; // @[Bitwise.scala 50:65:@3014.4]
  wire  _T_5077; // @[Bitwise.scala 50:65:@3015.4]
  wire  _T_5078; // @[Bitwise.scala 50:65:@3016.4]
  wire  _T_5079; // @[Bitwise.scala 50:65:@3017.4]
  wire  _T_5080; // @[Bitwise.scala 50:65:@3018.4]
  wire  _T_5081; // @[Bitwise.scala 50:65:@3019.4]
  wire  _T_5082; // @[Bitwise.scala 50:65:@3020.4]
  wire [1:0] _T_5083; // @[Bitwise.scala 48:55:@3021.4]
  wire [1:0] _GEN_655; // @[Bitwise.scala 48:55:@3022.4]
  wire [2:0] _T_5084; // @[Bitwise.scala 48:55:@3022.4]
  wire [1:0] _T_5085; // @[Bitwise.scala 48:55:@3023.4]
  wire [1:0] _T_5086; // @[Bitwise.scala 48:55:@3024.4]
  wire [2:0] _T_5087; // @[Bitwise.scala 48:55:@3025.4]
  wire [3:0] _T_5088; // @[Bitwise.scala 48:55:@3026.4]
  wire [1:0] _T_5089; // @[Bitwise.scala 48:55:@3027.4]
  wire [1:0] _T_5090; // @[Bitwise.scala 48:55:@3028.4]
  wire [2:0] _T_5091; // @[Bitwise.scala 48:55:@3029.4]
  wire [1:0] _T_5092; // @[Bitwise.scala 48:55:@3030.4]
  wire [1:0] _T_5093; // @[Bitwise.scala 48:55:@3031.4]
  wire [2:0] _T_5094; // @[Bitwise.scala 48:55:@3032.4]
  wire [3:0] _T_5095; // @[Bitwise.scala 48:55:@3033.4]
  wire [4:0] _T_5096; // @[Bitwise.scala 48:55:@3034.4]
  wire [1:0] _T_5097; // @[Bitwise.scala 48:55:@3035.4]
  wire [1:0] _T_5098; // @[Bitwise.scala 48:55:@3036.4]
  wire [2:0] _T_5099; // @[Bitwise.scala 48:55:@3037.4]
  wire [1:0] _T_5100; // @[Bitwise.scala 48:55:@3038.4]
  wire [1:0] _T_5101; // @[Bitwise.scala 48:55:@3039.4]
  wire [2:0] _T_5102; // @[Bitwise.scala 48:55:@3040.4]
  wire [3:0] _T_5103; // @[Bitwise.scala 48:55:@3041.4]
  wire [1:0] _T_5104; // @[Bitwise.scala 48:55:@3042.4]
  wire [1:0] _T_5105; // @[Bitwise.scala 48:55:@3043.4]
  wire [2:0] _T_5106; // @[Bitwise.scala 48:55:@3044.4]
  wire [1:0] _T_5107; // @[Bitwise.scala 48:55:@3045.4]
  wire [1:0] _T_5108; // @[Bitwise.scala 48:55:@3046.4]
  wire [2:0] _T_5109; // @[Bitwise.scala 48:55:@3047.4]
  wire [3:0] _T_5110; // @[Bitwise.scala 48:55:@3048.4]
  wire [4:0] _T_5111; // @[Bitwise.scala 48:55:@3049.4]
  wire [5:0] _T_5112; // @[Bitwise.scala 48:55:@3050.4]
  wire [31:0] _T_5176; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3115.4]
  wire  _T_5177; // @[Bitwise.scala 50:65:@3116.4]
  wire  _T_5178; // @[Bitwise.scala 50:65:@3117.4]
  wire  _T_5179; // @[Bitwise.scala 50:65:@3118.4]
  wire  _T_5180; // @[Bitwise.scala 50:65:@3119.4]
  wire  _T_5181; // @[Bitwise.scala 50:65:@3120.4]
  wire  _T_5182; // @[Bitwise.scala 50:65:@3121.4]
  wire  _T_5183; // @[Bitwise.scala 50:65:@3122.4]
  wire  _T_5184; // @[Bitwise.scala 50:65:@3123.4]
  wire  _T_5185; // @[Bitwise.scala 50:65:@3124.4]
  wire  _T_5186; // @[Bitwise.scala 50:65:@3125.4]
  wire  _T_5187; // @[Bitwise.scala 50:65:@3126.4]
  wire  _T_5188; // @[Bitwise.scala 50:65:@3127.4]
  wire  _T_5189; // @[Bitwise.scala 50:65:@3128.4]
  wire  _T_5190; // @[Bitwise.scala 50:65:@3129.4]
  wire  _T_5191; // @[Bitwise.scala 50:65:@3130.4]
  wire  _T_5192; // @[Bitwise.scala 50:65:@3131.4]
  wire  _T_5193; // @[Bitwise.scala 50:65:@3132.4]
  wire  _T_5194; // @[Bitwise.scala 50:65:@3133.4]
  wire  _T_5195; // @[Bitwise.scala 50:65:@3134.4]
  wire  _T_5196; // @[Bitwise.scala 50:65:@3135.4]
  wire  _T_5197; // @[Bitwise.scala 50:65:@3136.4]
  wire  _T_5198; // @[Bitwise.scala 50:65:@3137.4]
  wire  _T_5199; // @[Bitwise.scala 50:65:@3138.4]
  wire  _T_5200; // @[Bitwise.scala 50:65:@3139.4]
  wire  _T_5201; // @[Bitwise.scala 50:65:@3140.4]
  wire  _T_5202; // @[Bitwise.scala 50:65:@3141.4]
  wire  _T_5203; // @[Bitwise.scala 50:65:@3142.4]
  wire  _T_5204; // @[Bitwise.scala 50:65:@3143.4]
  wire  _T_5205; // @[Bitwise.scala 50:65:@3144.4]
  wire  _T_5206; // @[Bitwise.scala 50:65:@3145.4]
  wire  _T_5207; // @[Bitwise.scala 50:65:@3146.4]
  wire  _T_5208; // @[Bitwise.scala 50:65:@3147.4]
  wire [1:0] _T_5209; // @[Bitwise.scala 48:55:@3148.4]
  wire [1:0] _T_5210; // @[Bitwise.scala 48:55:@3149.4]
  wire [2:0] _T_5211; // @[Bitwise.scala 48:55:@3150.4]
  wire [1:0] _T_5212; // @[Bitwise.scala 48:55:@3151.4]
  wire [1:0] _T_5213; // @[Bitwise.scala 48:55:@3152.4]
  wire [2:0] _T_5214; // @[Bitwise.scala 48:55:@3153.4]
  wire [3:0] _T_5215; // @[Bitwise.scala 48:55:@3154.4]
  wire [1:0] _T_5216; // @[Bitwise.scala 48:55:@3155.4]
  wire [1:0] _T_5217; // @[Bitwise.scala 48:55:@3156.4]
  wire [2:0] _T_5218; // @[Bitwise.scala 48:55:@3157.4]
  wire [1:0] _T_5219; // @[Bitwise.scala 48:55:@3158.4]
  wire [1:0] _T_5220; // @[Bitwise.scala 48:55:@3159.4]
  wire [2:0] _T_5221; // @[Bitwise.scala 48:55:@3160.4]
  wire [3:0] _T_5222; // @[Bitwise.scala 48:55:@3161.4]
  wire [4:0] _T_5223; // @[Bitwise.scala 48:55:@3162.4]
  wire [1:0] _T_5224; // @[Bitwise.scala 48:55:@3163.4]
  wire [1:0] _T_5225; // @[Bitwise.scala 48:55:@3164.4]
  wire [2:0] _T_5226; // @[Bitwise.scala 48:55:@3165.4]
  wire [1:0] _T_5227; // @[Bitwise.scala 48:55:@3166.4]
  wire [1:0] _T_5228; // @[Bitwise.scala 48:55:@3167.4]
  wire [2:0] _T_5229; // @[Bitwise.scala 48:55:@3168.4]
  wire [3:0] _T_5230; // @[Bitwise.scala 48:55:@3169.4]
  wire [1:0] _T_5231; // @[Bitwise.scala 48:55:@3170.4]
  wire [1:0] _T_5232; // @[Bitwise.scala 48:55:@3171.4]
  wire [2:0] _T_5233; // @[Bitwise.scala 48:55:@3172.4]
  wire [1:0] _T_5234; // @[Bitwise.scala 48:55:@3173.4]
  wire [1:0] _T_5235; // @[Bitwise.scala 48:55:@3174.4]
  wire [2:0] _T_5236; // @[Bitwise.scala 48:55:@3175.4]
  wire [3:0] _T_5237; // @[Bitwise.scala 48:55:@3176.4]
  wire [4:0] _T_5238; // @[Bitwise.scala 48:55:@3177.4]
  wire [5:0] _T_5239; // @[Bitwise.scala 48:55:@3178.4]
  wire [32:0] _T_5303; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3243.4]
  wire  _T_5304; // @[Bitwise.scala 50:65:@3244.4]
  wire  _T_5305; // @[Bitwise.scala 50:65:@3245.4]
  wire  _T_5306; // @[Bitwise.scala 50:65:@3246.4]
  wire  _T_5307; // @[Bitwise.scala 50:65:@3247.4]
  wire  _T_5308; // @[Bitwise.scala 50:65:@3248.4]
  wire  _T_5309; // @[Bitwise.scala 50:65:@3249.4]
  wire  _T_5310; // @[Bitwise.scala 50:65:@3250.4]
  wire  _T_5311; // @[Bitwise.scala 50:65:@3251.4]
  wire  _T_5312; // @[Bitwise.scala 50:65:@3252.4]
  wire  _T_5313; // @[Bitwise.scala 50:65:@3253.4]
  wire  _T_5314; // @[Bitwise.scala 50:65:@3254.4]
  wire  _T_5315; // @[Bitwise.scala 50:65:@3255.4]
  wire  _T_5316; // @[Bitwise.scala 50:65:@3256.4]
  wire  _T_5317; // @[Bitwise.scala 50:65:@3257.4]
  wire  _T_5318; // @[Bitwise.scala 50:65:@3258.4]
  wire  _T_5319; // @[Bitwise.scala 50:65:@3259.4]
  wire  _T_5320; // @[Bitwise.scala 50:65:@3260.4]
  wire  _T_5321; // @[Bitwise.scala 50:65:@3261.4]
  wire  _T_5322; // @[Bitwise.scala 50:65:@3262.4]
  wire  _T_5323; // @[Bitwise.scala 50:65:@3263.4]
  wire  _T_5324; // @[Bitwise.scala 50:65:@3264.4]
  wire  _T_5325; // @[Bitwise.scala 50:65:@3265.4]
  wire  _T_5326; // @[Bitwise.scala 50:65:@3266.4]
  wire  _T_5327; // @[Bitwise.scala 50:65:@3267.4]
  wire  _T_5328; // @[Bitwise.scala 50:65:@3268.4]
  wire  _T_5329; // @[Bitwise.scala 50:65:@3269.4]
  wire  _T_5330; // @[Bitwise.scala 50:65:@3270.4]
  wire  _T_5331; // @[Bitwise.scala 50:65:@3271.4]
  wire  _T_5332; // @[Bitwise.scala 50:65:@3272.4]
  wire  _T_5333; // @[Bitwise.scala 50:65:@3273.4]
  wire  _T_5334; // @[Bitwise.scala 50:65:@3274.4]
  wire  _T_5335; // @[Bitwise.scala 50:65:@3275.4]
  wire  _T_5336; // @[Bitwise.scala 50:65:@3276.4]
  wire [1:0] _T_5337; // @[Bitwise.scala 48:55:@3277.4]
  wire [1:0] _T_5338; // @[Bitwise.scala 48:55:@3278.4]
  wire [2:0] _T_5339; // @[Bitwise.scala 48:55:@3279.4]
  wire [1:0] _T_5340; // @[Bitwise.scala 48:55:@3280.4]
  wire [1:0] _T_5341; // @[Bitwise.scala 48:55:@3281.4]
  wire [2:0] _T_5342; // @[Bitwise.scala 48:55:@3282.4]
  wire [3:0] _T_5343; // @[Bitwise.scala 48:55:@3283.4]
  wire [1:0] _T_5344; // @[Bitwise.scala 48:55:@3284.4]
  wire [1:0] _T_5345; // @[Bitwise.scala 48:55:@3285.4]
  wire [2:0] _T_5346; // @[Bitwise.scala 48:55:@3286.4]
  wire [1:0] _T_5347; // @[Bitwise.scala 48:55:@3287.4]
  wire [1:0] _T_5348; // @[Bitwise.scala 48:55:@3288.4]
  wire [2:0] _T_5349; // @[Bitwise.scala 48:55:@3289.4]
  wire [3:0] _T_5350; // @[Bitwise.scala 48:55:@3290.4]
  wire [4:0] _T_5351; // @[Bitwise.scala 48:55:@3291.4]
  wire [1:0] _T_5352; // @[Bitwise.scala 48:55:@3292.4]
  wire [1:0] _T_5353; // @[Bitwise.scala 48:55:@3293.4]
  wire [2:0] _T_5354; // @[Bitwise.scala 48:55:@3294.4]
  wire [1:0] _T_5355; // @[Bitwise.scala 48:55:@3295.4]
  wire [1:0] _T_5356; // @[Bitwise.scala 48:55:@3296.4]
  wire [2:0] _T_5357; // @[Bitwise.scala 48:55:@3297.4]
  wire [3:0] _T_5358; // @[Bitwise.scala 48:55:@3298.4]
  wire [1:0] _T_5359; // @[Bitwise.scala 48:55:@3299.4]
  wire [1:0] _T_5360; // @[Bitwise.scala 48:55:@3300.4]
  wire [2:0] _T_5361; // @[Bitwise.scala 48:55:@3301.4]
  wire [1:0] _T_5362; // @[Bitwise.scala 48:55:@3302.4]
  wire [1:0] _T_5363; // @[Bitwise.scala 48:55:@3303.4]
  wire [1:0] _GEN_656; // @[Bitwise.scala 48:55:@3304.4]
  wire [2:0] _T_5364; // @[Bitwise.scala 48:55:@3304.4]
  wire [2:0] _GEN_657; // @[Bitwise.scala 48:55:@3305.4]
  wire [3:0] _T_5365; // @[Bitwise.scala 48:55:@3305.4]
  wire [3:0] _GEN_658; // @[Bitwise.scala 48:55:@3306.4]
  wire [4:0] _T_5366; // @[Bitwise.scala 48:55:@3306.4]
  wire [4:0] _GEN_659; // @[Bitwise.scala 48:55:@3307.4]
  wire [5:0] _T_5367; // @[Bitwise.scala 48:55:@3307.4]
  wire [5:0] _GEN_660; // @[Bitwise.scala 48:55:@3308.4]
  wire [6:0] _T_5368; // @[Bitwise.scala 48:55:@3308.4]
  wire [33:0] _T_5432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3373.4]
  wire  _T_5433; // @[Bitwise.scala 50:65:@3374.4]
  wire  _T_5434; // @[Bitwise.scala 50:65:@3375.4]
  wire  _T_5435; // @[Bitwise.scala 50:65:@3376.4]
  wire  _T_5436; // @[Bitwise.scala 50:65:@3377.4]
  wire  _T_5437; // @[Bitwise.scala 50:65:@3378.4]
  wire  _T_5438; // @[Bitwise.scala 50:65:@3379.4]
  wire  _T_5439; // @[Bitwise.scala 50:65:@3380.4]
  wire  _T_5440; // @[Bitwise.scala 50:65:@3381.4]
  wire  _T_5441; // @[Bitwise.scala 50:65:@3382.4]
  wire  _T_5442; // @[Bitwise.scala 50:65:@3383.4]
  wire  _T_5443; // @[Bitwise.scala 50:65:@3384.4]
  wire  _T_5444; // @[Bitwise.scala 50:65:@3385.4]
  wire  _T_5445; // @[Bitwise.scala 50:65:@3386.4]
  wire  _T_5446; // @[Bitwise.scala 50:65:@3387.4]
  wire  _T_5447; // @[Bitwise.scala 50:65:@3388.4]
  wire  _T_5448; // @[Bitwise.scala 50:65:@3389.4]
  wire  _T_5449; // @[Bitwise.scala 50:65:@3390.4]
  wire  _T_5450; // @[Bitwise.scala 50:65:@3391.4]
  wire  _T_5451; // @[Bitwise.scala 50:65:@3392.4]
  wire  _T_5452; // @[Bitwise.scala 50:65:@3393.4]
  wire  _T_5453; // @[Bitwise.scala 50:65:@3394.4]
  wire  _T_5454; // @[Bitwise.scala 50:65:@3395.4]
  wire  _T_5455; // @[Bitwise.scala 50:65:@3396.4]
  wire  _T_5456; // @[Bitwise.scala 50:65:@3397.4]
  wire  _T_5457; // @[Bitwise.scala 50:65:@3398.4]
  wire  _T_5458; // @[Bitwise.scala 50:65:@3399.4]
  wire  _T_5459; // @[Bitwise.scala 50:65:@3400.4]
  wire  _T_5460; // @[Bitwise.scala 50:65:@3401.4]
  wire  _T_5461; // @[Bitwise.scala 50:65:@3402.4]
  wire  _T_5462; // @[Bitwise.scala 50:65:@3403.4]
  wire  _T_5463; // @[Bitwise.scala 50:65:@3404.4]
  wire  _T_5464; // @[Bitwise.scala 50:65:@3405.4]
  wire  _T_5465; // @[Bitwise.scala 50:65:@3406.4]
  wire  _T_5466; // @[Bitwise.scala 50:65:@3407.4]
  wire [1:0] _T_5467; // @[Bitwise.scala 48:55:@3408.4]
  wire [1:0] _T_5468; // @[Bitwise.scala 48:55:@3409.4]
  wire [2:0] _T_5469; // @[Bitwise.scala 48:55:@3410.4]
  wire [1:0] _T_5470; // @[Bitwise.scala 48:55:@3411.4]
  wire [1:0] _T_5471; // @[Bitwise.scala 48:55:@3412.4]
  wire [2:0] _T_5472; // @[Bitwise.scala 48:55:@3413.4]
  wire [3:0] _T_5473; // @[Bitwise.scala 48:55:@3414.4]
  wire [1:0] _T_5474; // @[Bitwise.scala 48:55:@3415.4]
  wire [1:0] _T_5475; // @[Bitwise.scala 48:55:@3416.4]
  wire [2:0] _T_5476; // @[Bitwise.scala 48:55:@3417.4]
  wire [1:0] _T_5477; // @[Bitwise.scala 48:55:@3418.4]
  wire [1:0] _T_5478; // @[Bitwise.scala 48:55:@3419.4]
  wire [1:0] _GEN_661; // @[Bitwise.scala 48:55:@3420.4]
  wire [2:0] _T_5479; // @[Bitwise.scala 48:55:@3420.4]
  wire [2:0] _GEN_662; // @[Bitwise.scala 48:55:@3421.4]
  wire [3:0] _T_5480; // @[Bitwise.scala 48:55:@3421.4]
  wire [3:0] _GEN_663; // @[Bitwise.scala 48:55:@3422.4]
  wire [4:0] _T_5481; // @[Bitwise.scala 48:55:@3422.4]
  wire [4:0] _GEN_664; // @[Bitwise.scala 48:55:@3423.4]
  wire [5:0] _T_5482; // @[Bitwise.scala 48:55:@3423.4]
  wire [1:0] _T_5483; // @[Bitwise.scala 48:55:@3424.4]
  wire [1:0] _T_5484; // @[Bitwise.scala 48:55:@3425.4]
  wire [2:0] _T_5485; // @[Bitwise.scala 48:55:@3426.4]
  wire [1:0] _T_5486; // @[Bitwise.scala 48:55:@3427.4]
  wire [1:0] _T_5487; // @[Bitwise.scala 48:55:@3428.4]
  wire [2:0] _T_5488; // @[Bitwise.scala 48:55:@3429.4]
  wire [3:0] _T_5489; // @[Bitwise.scala 48:55:@3430.4]
  wire [1:0] _T_5490; // @[Bitwise.scala 48:55:@3431.4]
  wire [1:0] _T_5491; // @[Bitwise.scala 48:55:@3432.4]
  wire [2:0] _T_5492; // @[Bitwise.scala 48:55:@3433.4]
  wire [1:0] _T_5493; // @[Bitwise.scala 48:55:@3434.4]
  wire [1:0] _T_5494; // @[Bitwise.scala 48:55:@3435.4]
  wire [1:0] _GEN_665; // @[Bitwise.scala 48:55:@3436.4]
  wire [2:0] _T_5495; // @[Bitwise.scala 48:55:@3436.4]
  wire [2:0] _GEN_666; // @[Bitwise.scala 48:55:@3437.4]
  wire [3:0] _T_5496; // @[Bitwise.scala 48:55:@3437.4]
  wire [3:0] _GEN_667; // @[Bitwise.scala 48:55:@3438.4]
  wire [4:0] _T_5497; // @[Bitwise.scala 48:55:@3438.4]
  wire [4:0] _GEN_668; // @[Bitwise.scala 48:55:@3439.4]
  wire [5:0] _T_5498; // @[Bitwise.scala 48:55:@3439.4]
  wire [6:0] _T_5499; // @[Bitwise.scala 48:55:@3440.4]
  wire [34:0] _T_5563; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3505.4]
  wire  _T_5564; // @[Bitwise.scala 50:65:@3506.4]
  wire  _T_5565; // @[Bitwise.scala 50:65:@3507.4]
  wire  _T_5566; // @[Bitwise.scala 50:65:@3508.4]
  wire  _T_5567; // @[Bitwise.scala 50:65:@3509.4]
  wire  _T_5568; // @[Bitwise.scala 50:65:@3510.4]
  wire  _T_5569; // @[Bitwise.scala 50:65:@3511.4]
  wire  _T_5570; // @[Bitwise.scala 50:65:@3512.4]
  wire  _T_5571; // @[Bitwise.scala 50:65:@3513.4]
  wire  _T_5572; // @[Bitwise.scala 50:65:@3514.4]
  wire  _T_5573; // @[Bitwise.scala 50:65:@3515.4]
  wire  _T_5574; // @[Bitwise.scala 50:65:@3516.4]
  wire  _T_5575; // @[Bitwise.scala 50:65:@3517.4]
  wire  _T_5576; // @[Bitwise.scala 50:65:@3518.4]
  wire  _T_5577; // @[Bitwise.scala 50:65:@3519.4]
  wire  _T_5578; // @[Bitwise.scala 50:65:@3520.4]
  wire  _T_5579; // @[Bitwise.scala 50:65:@3521.4]
  wire  _T_5580; // @[Bitwise.scala 50:65:@3522.4]
  wire  _T_5581; // @[Bitwise.scala 50:65:@3523.4]
  wire  _T_5582; // @[Bitwise.scala 50:65:@3524.4]
  wire  _T_5583; // @[Bitwise.scala 50:65:@3525.4]
  wire  _T_5584; // @[Bitwise.scala 50:65:@3526.4]
  wire  _T_5585; // @[Bitwise.scala 50:65:@3527.4]
  wire  _T_5586; // @[Bitwise.scala 50:65:@3528.4]
  wire  _T_5587; // @[Bitwise.scala 50:65:@3529.4]
  wire  _T_5588; // @[Bitwise.scala 50:65:@3530.4]
  wire  _T_5589; // @[Bitwise.scala 50:65:@3531.4]
  wire  _T_5590; // @[Bitwise.scala 50:65:@3532.4]
  wire  _T_5591; // @[Bitwise.scala 50:65:@3533.4]
  wire  _T_5592; // @[Bitwise.scala 50:65:@3534.4]
  wire  _T_5593; // @[Bitwise.scala 50:65:@3535.4]
  wire  _T_5594; // @[Bitwise.scala 50:65:@3536.4]
  wire  _T_5595; // @[Bitwise.scala 50:65:@3537.4]
  wire  _T_5596; // @[Bitwise.scala 50:65:@3538.4]
  wire  _T_5597; // @[Bitwise.scala 50:65:@3539.4]
  wire  _T_5598; // @[Bitwise.scala 50:65:@3540.4]
  wire [1:0] _T_5599; // @[Bitwise.scala 48:55:@3541.4]
  wire [1:0] _T_5600; // @[Bitwise.scala 48:55:@3542.4]
  wire [2:0] _T_5601; // @[Bitwise.scala 48:55:@3543.4]
  wire [1:0] _T_5602; // @[Bitwise.scala 48:55:@3544.4]
  wire [1:0] _T_5603; // @[Bitwise.scala 48:55:@3545.4]
  wire [2:0] _T_5604; // @[Bitwise.scala 48:55:@3546.4]
  wire [3:0] _T_5605; // @[Bitwise.scala 48:55:@3547.4]
  wire [1:0] _T_5606; // @[Bitwise.scala 48:55:@3548.4]
  wire [1:0] _T_5607; // @[Bitwise.scala 48:55:@3549.4]
  wire [2:0] _T_5608; // @[Bitwise.scala 48:55:@3550.4]
  wire [1:0] _T_5609; // @[Bitwise.scala 48:55:@3551.4]
  wire [1:0] _T_5610; // @[Bitwise.scala 48:55:@3552.4]
  wire [1:0] _GEN_669; // @[Bitwise.scala 48:55:@3553.4]
  wire [2:0] _T_5611; // @[Bitwise.scala 48:55:@3553.4]
  wire [2:0] _GEN_670; // @[Bitwise.scala 48:55:@3554.4]
  wire [3:0] _T_5612; // @[Bitwise.scala 48:55:@3554.4]
  wire [3:0] _GEN_671; // @[Bitwise.scala 48:55:@3555.4]
  wire [4:0] _T_5613; // @[Bitwise.scala 48:55:@3555.4]
  wire [4:0] _GEN_672; // @[Bitwise.scala 48:55:@3556.4]
  wire [5:0] _T_5614; // @[Bitwise.scala 48:55:@3556.4]
  wire [1:0] _T_5615; // @[Bitwise.scala 48:55:@3557.4]
  wire [1:0] _T_5616; // @[Bitwise.scala 48:55:@3558.4]
  wire [2:0] _T_5617; // @[Bitwise.scala 48:55:@3559.4]
  wire [1:0] _T_5618; // @[Bitwise.scala 48:55:@3560.4]
  wire [1:0] _T_5619; // @[Bitwise.scala 48:55:@3561.4]
  wire [1:0] _GEN_673; // @[Bitwise.scala 48:55:@3562.4]
  wire [2:0] _T_5620; // @[Bitwise.scala 48:55:@3562.4]
  wire [2:0] _GEN_674; // @[Bitwise.scala 48:55:@3563.4]
  wire [3:0] _T_5621; // @[Bitwise.scala 48:55:@3563.4]
  wire [3:0] _GEN_675; // @[Bitwise.scala 48:55:@3564.4]
  wire [4:0] _T_5622; // @[Bitwise.scala 48:55:@3564.4]
  wire [1:0] _T_5623; // @[Bitwise.scala 48:55:@3565.4]
  wire [1:0] _T_5624; // @[Bitwise.scala 48:55:@3566.4]
  wire [2:0] _T_5625; // @[Bitwise.scala 48:55:@3567.4]
  wire [1:0] _T_5626; // @[Bitwise.scala 48:55:@3568.4]
  wire [1:0] _T_5627; // @[Bitwise.scala 48:55:@3569.4]
  wire [1:0] _GEN_676; // @[Bitwise.scala 48:55:@3570.4]
  wire [2:0] _T_5628; // @[Bitwise.scala 48:55:@3570.4]
  wire [2:0] _GEN_677; // @[Bitwise.scala 48:55:@3571.4]
  wire [3:0] _T_5629; // @[Bitwise.scala 48:55:@3571.4]
  wire [3:0] _GEN_678; // @[Bitwise.scala 48:55:@3572.4]
  wire [4:0] _T_5630; // @[Bitwise.scala 48:55:@3572.4]
  wire [5:0] _T_5631; // @[Bitwise.scala 48:55:@3573.4]
  wire [6:0] _T_5632; // @[Bitwise.scala 48:55:@3574.4]
  wire [35:0] _T_5696; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3639.4]
  wire  _T_5697; // @[Bitwise.scala 50:65:@3640.4]
  wire  _T_5698; // @[Bitwise.scala 50:65:@3641.4]
  wire  _T_5699; // @[Bitwise.scala 50:65:@3642.4]
  wire  _T_5700; // @[Bitwise.scala 50:65:@3643.4]
  wire  _T_5701; // @[Bitwise.scala 50:65:@3644.4]
  wire  _T_5702; // @[Bitwise.scala 50:65:@3645.4]
  wire  _T_5703; // @[Bitwise.scala 50:65:@3646.4]
  wire  _T_5704; // @[Bitwise.scala 50:65:@3647.4]
  wire  _T_5705; // @[Bitwise.scala 50:65:@3648.4]
  wire  _T_5706; // @[Bitwise.scala 50:65:@3649.4]
  wire  _T_5707; // @[Bitwise.scala 50:65:@3650.4]
  wire  _T_5708; // @[Bitwise.scala 50:65:@3651.4]
  wire  _T_5709; // @[Bitwise.scala 50:65:@3652.4]
  wire  _T_5710; // @[Bitwise.scala 50:65:@3653.4]
  wire  _T_5711; // @[Bitwise.scala 50:65:@3654.4]
  wire  _T_5712; // @[Bitwise.scala 50:65:@3655.4]
  wire  _T_5713; // @[Bitwise.scala 50:65:@3656.4]
  wire  _T_5714; // @[Bitwise.scala 50:65:@3657.4]
  wire  _T_5715; // @[Bitwise.scala 50:65:@3658.4]
  wire  _T_5716; // @[Bitwise.scala 50:65:@3659.4]
  wire  _T_5717; // @[Bitwise.scala 50:65:@3660.4]
  wire  _T_5718; // @[Bitwise.scala 50:65:@3661.4]
  wire  _T_5719; // @[Bitwise.scala 50:65:@3662.4]
  wire  _T_5720; // @[Bitwise.scala 50:65:@3663.4]
  wire  _T_5721; // @[Bitwise.scala 50:65:@3664.4]
  wire  _T_5722; // @[Bitwise.scala 50:65:@3665.4]
  wire  _T_5723; // @[Bitwise.scala 50:65:@3666.4]
  wire  _T_5724; // @[Bitwise.scala 50:65:@3667.4]
  wire  _T_5725; // @[Bitwise.scala 50:65:@3668.4]
  wire  _T_5726; // @[Bitwise.scala 50:65:@3669.4]
  wire  _T_5727; // @[Bitwise.scala 50:65:@3670.4]
  wire  _T_5728; // @[Bitwise.scala 50:65:@3671.4]
  wire  _T_5729; // @[Bitwise.scala 50:65:@3672.4]
  wire  _T_5730; // @[Bitwise.scala 50:65:@3673.4]
  wire  _T_5731; // @[Bitwise.scala 50:65:@3674.4]
  wire  _T_5732; // @[Bitwise.scala 50:65:@3675.4]
  wire [1:0] _T_5733; // @[Bitwise.scala 48:55:@3676.4]
  wire [1:0] _T_5734; // @[Bitwise.scala 48:55:@3677.4]
  wire [2:0] _T_5735; // @[Bitwise.scala 48:55:@3678.4]
  wire [1:0] _T_5736; // @[Bitwise.scala 48:55:@3679.4]
  wire [1:0] _T_5737; // @[Bitwise.scala 48:55:@3680.4]
  wire [1:0] _GEN_679; // @[Bitwise.scala 48:55:@3681.4]
  wire [2:0] _T_5738; // @[Bitwise.scala 48:55:@3681.4]
  wire [2:0] _GEN_680; // @[Bitwise.scala 48:55:@3682.4]
  wire [3:0] _T_5739; // @[Bitwise.scala 48:55:@3682.4]
  wire [3:0] _GEN_681; // @[Bitwise.scala 48:55:@3683.4]
  wire [4:0] _T_5740; // @[Bitwise.scala 48:55:@3683.4]
  wire [1:0] _T_5741; // @[Bitwise.scala 48:55:@3684.4]
  wire [1:0] _T_5742; // @[Bitwise.scala 48:55:@3685.4]
  wire [2:0] _T_5743; // @[Bitwise.scala 48:55:@3686.4]
  wire [1:0] _T_5744; // @[Bitwise.scala 48:55:@3687.4]
  wire [1:0] _T_5745; // @[Bitwise.scala 48:55:@3688.4]
  wire [1:0] _GEN_682; // @[Bitwise.scala 48:55:@3689.4]
  wire [2:0] _T_5746; // @[Bitwise.scala 48:55:@3689.4]
  wire [2:0] _GEN_683; // @[Bitwise.scala 48:55:@3690.4]
  wire [3:0] _T_5747; // @[Bitwise.scala 48:55:@3690.4]
  wire [3:0] _GEN_684; // @[Bitwise.scala 48:55:@3691.4]
  wire [4:0] _T_5748; // @[Bitwise.scala 48:55:@3691.4]
  wire [5:0] _T_5749; // @[Bitwise.scala 48:55:@3692.4]
  wire [1:0] _T_5750; // @[Bitwise.scala 48:55:@3693.4]
  wire [1:0] _T_5751; // @[Bitwise.scala 48:55:@3694.4]
  wire [2:0] _T_5752; // @[Bitwise.scala 48:55:@3695.4]
  wire [1:0] _T_5753; // @[Bitwise.scala 48:55:@3696.4]
  wire [1:0] _T_5754; // @[Bitwise.scala 48:55:@3697.4]
  wire [1:0] _GEN_685; // @[Bitwise.scala 48:55:@3698.4]
  wire [2:0] _T_5755; // @[Bitwise.scala 48:55:@3698.4]
  wire [2:0] _GEN_686; // @[Bitwise.scala 48:55:@3699.4]
  wire [3:0] _T_5756; // @[Bitwise.scala 48:55:@3699.4]
  wire [3:0] _GEN_687; // @[Bitwise.scala 48:55:@3700.4]
  wire [4:0] _T_5757; // @[Bitwise.scala 48:55:@3700.4]
  wire [1:0] _T_5758; // @[Bitwise.scala 48:55:@3701.4]
  wire [1:0] _T_5759; // @[Bitwise.scala 48:55:@3702.4]
  wire [2:0] _T_5760; // @[Bitwise.scala 48:55:@3703.4]
  wire [1:0] _T_5761; // @[Bitwise.scala 48:55:@3704.4]
  wire [1:0] _T_5762; // @[Bitwise.scala 48:55:@3705.4]
  wire [1:0] _GEN_688; // @[Bitwise.scala 48:55:@3706.4]
  wire [2:0] _T_5763; // @[Bitwise.scala 48:55:@3706.4]
  wire [2:0] _GEN_689; // @[Bitwise.scala 48:55:@3707.4]
  wire [3:0] _T_5764; // @[Bitwise.scala 48:55:@3707.4]
  wire [3:0] _GEN_690; // @[Bitwise.scala 48:55:@3708.4]
  wire [4:0] _T_5765; // @[Bitwise.scala 48:55:@3708.4]
  wire [5:0] _T_5766; // @[Bitwise.scala 48:55:@3709.4]
  wire [6:0] _T_5767; // @[Bitwise.scala 48:55:@3710.4]
  wire [36:0] _T_5831; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3775.4]
  wire  _T_5832; // @[Bitwise.scala 50:65:@3776.4]
  wire  _T_5833; // @[Bitwise.scala 50:65:@3777.4]
  wire  _T_5834; // @[Bitwise.scala 50:65:@3778.4]
  wire  _T_5835; // @[Bitwise.scala 50:65:@3779.4]
  wire  _T_5836; // @[Bitwise.scala 50:65:@3780.4]
  wire  _T_5837; // @[Bitwise.scala 50:65:@3781.4]
  wire  _T_5838; // @[Bitwise.scala 50:65:@3782.4]
  wire  _T_5839; // @[Bitwise.scala 50:65:@3783.4]
  wire  _T_5840; // @[Bitwise.scala 50:65:@3784.4]
  wire  _T_5841; // @[Bitwise.scala 50:65:@3785.4]
  wire  _T_5842; // @[Bitwise.scala 50:65:@3786.4]
  wire  _T_5843; // @[Bitwise.scala 50:65:@3787.4]
  wire  _T_5844; // @[Bitwise.scala 50:65:@3788.4]
  wire  _T_5845; // @[Bitwise.scala 50:65:@3789.4]
  wire  _T_5846; // @[Bitwise.scala 50:65:@3790.4]
  wire  _T_5847; // @[Bitwise.scala 50:65:@3791.4]
  wire  _T_5848; // @[Bitwise.scala 50:65:@3792.4]
  wire  _T_5849; // @[Bitwise.scala 50:65:@3793.4]
  wire  _T_5850; // @[Bitwise.scala 50:65:@3794.4]
  wire  _T_5851; // @[Bitwise.scala 50:65:@3795.4]
  wire  _T_5852; // @[Bitwise.scala 50:65:@3796.4]
  wire  _T_5853; // @[Bitwise.scala 50:65:@3797.4]
  wire  _T_5854; // @[Bitwise.scala 50:65:@3798.4]
  wire  _T_5855; // @[Bitwise.scala 50:65:@3799.4]
  wire  _T_5856; // @[Bitwise.scala 50:65:@3800.4]
  wire  _T_5857; // @[Bitwise.scala 50:65:@3801.4]
  wire  _T_5858; // @[Bitwise.scala 50:65:@3802.4]
  wire  _T_5859; // @[Bitwise.scala 50:65:@3803.4]
  wire  _T_5860; // @[Bitwise.scala 50:65:@3804.4]
  wire  _T_5861; // @[Bitwise.scala 50:65:@3805.4]
  wire  _T_5862; // @[Bitwise.scala 50:65:@3806.4]
  wire  _T_5863; // @[Bitwise.scala 50:65:@3807.4]
  wire  _T_5864; // @[Bitwise.scala 50:65:@3808.4]
  wire  _T_5865; // @[Bitwise.scala 50:65:@3809.4]
  wire  _T_5866; // @[Bitwise.scala 50:65:@3810.4]
  wire  _T_5867; // @[Bitwise.scala 50:65:@3811.4]
  wire  _T_5868; // @[Bitwise.scala 50:65:@3812.4]
  wire [1:0] _T_5869; // @[Bitwise.scala 48:55:@3813.4]
  wire [1:0] _T_5870; // @[Bitwise.scala 48:55:@3814.4]
  wire [2:0] _T_5871; // @[Bitwise.scala 48:55:@3815.4]
  wire [1:0] _T_5872; // @[Bitwise.scala 48:55:@3816.4]
  wire [1:0] _T_5873; // @[Bitwise.scala 48:55:@3817.4]
  wire [1:0] _GEN_691; // @[Bitwise.scala 48:55:@3818.4]
  wire [2:0] _T_5874; // @[Bitwise.scala 48:55:@3818.4]
  wire [2:0] _GEN_692; // @[Bitwise.scala 48:55:@3819.4]
  wire [3:0] _T_5875; // @[Bitwise.scala 48:55:@3819.4]
  wire [3:0] _GEN_693; // @[Bitwise.scala 48:55:@3820.4]
  wire [4:0] _T_5876; // @[Bitwise.scala 48:55:@3820.4]
  wire [1:0] _T_5877; // @[Bitwise.scala 48:55:@3821.4]
  wire [1:0] _T_5878; // @[Bitwise.scala 48:55:@3822.4]
  wire [2:0] _T_5879; // @[Bitwise.scala 48:55:@3823.4]
  wire [1:0] _T_5880; // @[Bitwise.scala 48:55:@3824.4]
  wire [1:0] _T_5881; // @[Bitwise.scala 48:55:@3825.4]
  wire [1:0] _GEN_694; // @[Bitwise.scala 48:55:@3826.4]
  wire [2:0] _T_5882; // @[Bitwise.scala 48:55:@3826.4]
  wire [2:0] _GEN_695; // @[Bitwise.scala 48:55:@3827.4]
  wire [3:0] _T_5883; // @[Bitwise.scala 48:55:@3827.4]
  wire [3:0] _GEN_696; // @[Bitwise.scala 48:55:@3828.4]
  wire [4:0] _T_5884; // @[Bitwise.scala 48:55:@3828.4]
  wire [5:0] _T_5885; // @[Bitwise.scala 48:55:@3829.4]
  wire [1:0] _T_5886; // @[Bitwise.scala 48:55:@3830.4]
  wire [1:0] _T_5887; // @[Bitwise.scala 48:55:@3831.4]
  wire [2:0] _T_5888; // @[Bitwise.scala 48:55:@3832.4]
  wire [1:0] _T_5889; // @[Bitwise.scala 48:55:@3833.4]
  wire [1:0] _T_5890; // @[Bitwise.scala 48:55:@3834.4]
  wire [1:0] _GEN_697; // @[Bitwise.scala 48:55:@3835.4]
  wire [2:0] _T_5891; // @[Bitwise.scala 48:55:@3835.4]
  wire [2:0] _GEN_698; // @[Bitwise.scala 48:55:@3836.4]
  wire [3:0] _T_5892; // @[Bitwise.scala 48:55:@3836.4]
  wire [3:0] _GEN_699; // @[Bitwise.scala 48:55:@3837.4]
  wire [4:0] _T_5893; // @[Bitwise.scala 48:55:@3837.4]
  wire [1:0] _T_5894; // @[Bitwise.scala 48:55:@3838.4]
  wire [1:0] _T_5895; // @[Bitwise.scala 48:55:@3839.4]
  wire [1:0] _GEN_700; // @[Bitwise.scala 48:55:@3840.4]
  wire [2:0] _T_5896; // @[Bitwise.scala 48:55:@3840.4]
  wire [2:0] _GEN_701; // @[Bitwise.scala 48:55:@3841.4]
  wire [3:0] _T_5897; // @[Bitwise.scala 48:55:@3841.4]
  wire [1:0] _T_5898; // @[Bitwise.scala 48:55:@3842.4]
  wire [1:0] _T_5899; // @[Bitwise.scala 48:55:@3843.4]
  wire [1:0] _GEN_702; // @[Bitwise.scala 48:55:@3844.4]
  wire [2:0] _T_5900; // @[Bitwise.scala 48:55:@3844.4]
  wire [2:0] _GEN_703; // @[Bitwise.scala 48:55:@3845.4]
  wire [3:0] _T_5901; // @[Bitwise.scala 48:55:@3845.4]
  wire [4:0] _T_5902; // @[Bitwise.scala 48:55:@3846.4]
  wire [5:0] _T_5903; // @[Bitwise.scala 48:55:@3847.4]
  wire [6:0] _T_5904; // @[Bitwise.scala 48:55:@3848.4]
  wire [37:0] _T_5968; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3913.4]
  wire  _T_5969; // @[Bitwise.scala 50:65:@3914.4]
  wire  _T_5970; // @[Bitwise.scala 50:65:@3915.4]
  wire  _T_5971; // @[Bitwise.scala 50:65:@3916.4]
  wire  _T_5972; // @[Bitwise.scala 50:65:@3917.4]
  wire  _T_5973; // @[Bitwise.scala 50:65:@3918.4]
  wire  _T_5974; // @[Bitwise.scala 50:65:@3919.4]
  wire  _T_5975; // @[Bitwise.scala 50:65:@3920.4]
  wire  _T_5976; // @[Bitwise.scala 50:65:@3921.4]
  wire  _T_5977; // @[Bitwise.scala 50:65:@3922.4]
  wire  _T_5978; // @[Bitwise.scala 50:65:@3923.4]
  wire  _T_5979; // @[Bitwise.scala 50:65:@3924.4]
  wire  _T_5980; // @[Bitwise.scala 50:65:@3925.4]
  wire  _T_5981; // @[Bitwise.scala 50:65:@3926.4]
  wire  _T_5982; // @[Bitwise.scala 50:65:@3927.4]
  wire  _T_5983; // @[Bitwise.scala 50:65:@3928.4]
  wire  _T_5984; // @[Bitwise.scala 50:65:@3929.4]
  wire  _T_5985; // @[Bitwise.scala 50:65:@3930.4]
  wire  _T_5986; // @[Bitwise.scala 50:65:@3931.4]
  wire  _T_5987; // @[Bitwise.scala 50:65:@3932.4]
  wire  _T_5988; // @[Bitwise.scala 50:65:@3933.4]
  wire  _T_5989; // @[Bitwise.scala 50:65:@3934.4]
  wire  _T_5990; // @[Bitwise.scala 50:65:@3935.4]
  wire  _T_5991; // @[Bitwise.scala 50:65:@3936.4]
  wire  _T_5992; // @[Bitwise.scala 50:65:@3937.4]
  wire  _T_5993; // @[Bitwise.scala 50:65:@3938.4]
  wire  _T_5994; // @[Bitwise.scala 50:65:@3939.4]
  wire  _T_5995; // @[Bitwise.scala 50:65:@3940.4]
  wire  _T_5996; // @[Bitwise.scala 50:65:@3941.4]
  wire  _T_5997; // @[Bitwise.scala 50:65:@3942.4]
  wire  _T_5998; // @[Bitwise.scala 50:65:@3943.4]
  wire  _T_5999; // @[Bitwise.scala 50:65:@3944.4]
  wire  _T_6000; // @[Bitwise.scala 50:65:@3945.4]
  wire  _T_6001; // @[Bitwise.scala 50:65:@3946.4]
  wire  _T_6002; // @[Bitwise.scala 50:65:@3947.4]
  wire  _T_6003; // @[Bitwise.scala 50:65:@3948.4]
  wire  _T_6004; // @[Bitwise.scala 50:65:@3949.4]
  wire  _T_6005; // @[Bitwise.scala 50:65:@3950.4]
  wire  _T_6006; // @[Bitwise.scala 50:65:@3951.4]
  wire [1:0] _T_6007; // @[Bitwise.scala 48:55:@3952.4]
  wire [1:0] _T_6008; // @[Bitwise.scala 48:55:@3953.4]
  wire [2:0] _T_6009; // @[Bitwise.scala 48:55:@3954.4]
  wire [1:0] _T_6010; // @[Bitwise.scala 48:55:@3955.4]
  wire [1:0] _T_6011; // @[Bitwise.scala 48:55:@3956.4]
  wire [1:0] _GEN_704; // @[Bitwise.scala 48:55:@3957.4]
  wire [2:0] _T_6012; // @[Bitwise.scala 48:55:@3957.4]
  wire [2:0] _GEN_705; // @[Bitwise.scala 48:55:@3958.4]
  wire [3:0] _T_6013; // @[Bitwise.scala 48:55:@3958.4]
  wire [3:0] _GEN_706; // @[Bitwise.scala 48:55:@3959.4]
  wire [4:0] _T_6014; // @[Bitwise.scala 48:55:@3959.4]
  wire [1:0] _T_6015; // @[Bitwise.scala 48:55:@3960.4]
  wire [1:0] _T_6016; // @[Bitwise.scala 48:55:@3961.4]
  wire [1:0] _GEN_707; // @[Bitwise.scala 48:55:@3962.4]
  wire [2:0] _T_6017; // @[Bitwise.scala 48:55:@3962.4]
  wire [2:0] _GEN_708; // @[Bitwise.scala 48:55:@3963.4]
  wire [3:0] _T_6018; // @[Bitwise.scala 48:55:@3963.4]
  wire [1:0] _T_6019; // @[Bitwise.scala 48:55:@3964.4]
  wire [1:0] _T_6020; // @[Bitwise.scala 48:55:@3965.4]
  wire [1:0] _GEN_709; // @[Bitwise.scala 48:55:@3966.4]
  wire [2:0] _T_6021; // @[Bitwise.scala 48:55:@3966.4]
  wire [2:0] _GEN_710; // @[Bitwise.scala 48:55:@3967.4]
  wire [3:0] _T_6022; // @[Bitwise.scala 48:55:@3967.4]
  wire [4:0] _T_6023; // @[Bitwise.scala 48:55:@3968.4]
  wire [5:0] _T_6024; // @[Bitwise.scala 48:55:@3969.4]
  wire [1:0] _T_6025; // @[Bitwise.scala 48:55:@3970.4]
  wire [1:0] _T_6026; // @[Bitwise.scala 48:55:@3971.4]
  wire [2:0] _T_6027; // @[Bitwise.scala 48:55:@3972.4]
  wire [1:0] _T_6028; // @[Bitwise.scala 48:55:@3973.4]
  wire [1:0] _T_6029; // @[Bitwise.scala 48:55:@3974.4]
  wire [1:0] _GEN_711; // @[Bitwise.scala 48:55:@3975.4]
  wire [2:0] _T_6030; // @[Bitwise.scala 48:55:@3975.4]
  wire [2:0] _GEN_712; // @[Bitwise.scala 48:55:@3976.4]
  wire [3:0] _T_6031; // @[Bitwise.scala 48:55:@3976.4]
  wire [3:0] _GEN_713; // @[Bitwise.scala 48:55:@3977.4]
  wire [4:0] _T_6032; // @[Bitwise.scala 48:55:@3977.4]
  wire [1:0] _T_6033; // @[Bitwise.scala 48:55:@3978.4]
  wire [1:0] _T_6034; // @[Bitwise.scala 48:55:@3979.4]
  wire [1:0] _GEN_714; // @[Bitwise.scala 48:55:@3980.4]
  wire [2:0] _T_6035; // @[Bitwise.scala 48:55:@3980.4]
  wire [2:0] _GEN_715; // @[Bitwise.scala 48:55:@3981.4]
  wire [3:0] _T_6036; // @[Bitwise.scala 48:55:@3981.4]
  wire [1:0] _T_6037; // @[Bitwise.scala 48:55:@3982.4]
  wire [1:0] _T_6038; // @[Bitwise.scala 48:55:@3983.4]
  wire [1:0] _GEN_716; // @[Bitwise.scala 48:55:@3984.4]
  wire [2:0] _T_6039; // @[Bitwise.scala 48:55:@3984.4]
  wire [2:0] _GEN_717; // @[Bitwise.scala 48:55:@3985.4]
  wire [3:0] _T_6040; // @[Bitwise.scala 48:55:@3985.4]
  wire [4:0] _T_6041; // @[Bitwise.scala 48:55:@3986.4]
  wire [5:0] _T_6042; // @[Bitwise.scala 48:55:@3987.4]
  wire [6:0] _T_6043; // @[Bitwise.scala 48:55:@3988.4]
  wire [38:0] _T_6107; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4053.4]
  wire  _T_6108; // @[Bitwise.scala 50:65:@4054.4]
  wire  _T_6109; // @[Bitwise.scala 50:65:@4055.4]
  wire  _T_6110; // @[Bitwise.scala 50:65:@4056.4]
  wire  _T_6111; // @[Bitwise.scala 50:65:@4057.4]
  wire  _T_6112; // @[Bitwise.scala 50:65:@4058.4]
  wire  _T_6113; // @[Bitwise.scala 50:65:@4059.4]
  wire  _T_6114; // @[Bitwise.scala 50:65:@4060.4]
  wire  _T_6115; // @[Bitwise.scala 50:65:@4061.4]
  wire  _T_6116; // @[Bitwise.scala 50:65:@4062.4]
  wire  _T_6117; // @[Bitwise.scala 50:65:@4063.4]
  wire  _T_6118; // @[Bitwise.scala 50:65:@4064.4]
  wire  _T_6119; // @[Bitwise.scala 50:65:@4065.4]
  wire  _T_6120; // @[Bitwise.scala 50:65:@4066.4]
  wire  _T_6121; // @[Bitwise.scala 50:65:@4067.4]
  wire  _T_6122; // @[Bitwise.scala 50:65:@4068.4]
  wire  _T_6123; // @[Bitwise.scala 50:65:@4069.4]
  wire  _T_6124; // @[Bitwise.scala 50:65:@4070.4]
  wire  _T_6125; // @[Bitwise.scala 50:65:@4071.4]
  wire  _T_6126; // @[Bitwise.scala 50:65:@4072.4]
  wire  _T_6127; // @[Bitwise.scala 50:65:@4073.4]
  wire  _T_6128; // @[Bitwise.scala 50:65:@4074.4]
  wire  _T_6129; // @[Bitwise.scala 50:65:@4075.4]
  wire  _T_6130; // @[Bitwise.scala 50:65:@4076.4]
  wire  _T_6131; // @[Bitwise.scala 50:65:@4077.4]
  wire  _T_6132; // @[Bitwise.scala 50:65:@4078.4]
  wire  _T_6133; // @[Bitwise.scala 50:65:@4079.4]
  wire  _T_6134; // @[Bitwise.scala 50:65:@4080.4]
  wire  _T_6135; // @[Bitwise.scala 50:65:@4081.4]
  wire  _T_6136; // @[Bitwise.scala 50:65:@4082.4]
  wire  _T_6137; // @[Bitwise.scala 50:65:@4083.4]
  wire  _T_6138; // @[Bitwise.scala 50:65:@4084.4]
  wire  _T_6139; // @[Bitwise.scala 50:65:@4085.4]
  wire  _T_6140; // @[Bitwise.scala 50:65:@4086.4]
  wire  _T_6141; // @[Bitwise.scala 50:65:@4087.4]
  wire  _T_6142; // @[Bitwise.scala 50:65:@4088.4]
  wire  _T_6143; // @[Bitwise.scala 50:65:@4089.4]
  wire  _T_6144; // @[Bitwise.scala 50:65:@4090.4]
  wire  _T_6145; // @[Bitwise.scala 50:65:@4091.4]
  wire  _T_6146; // @[Bitwise.scala 50:65:@4092.4]
  wire [1:0] _T_6147; // @[Bitwise.scala 48:55:@4093.4]
  wire [1:0] _T_6148; // @[Bitwise.scala 48:55:@4094.4]
  wire [2:0] _T_6149; // @[Bitwise.scala 48:55:@4095.4]
  wire [1:0] _T_6150; // @[Bitwise.scala 48:55:@4096.4]
  wire [1:0] _T_6151; // @[Bitwise.scala 48:55:@4097.4]
  wire [1:0] _GEN_718; // @[Bitwise.scala 48:55:@4098.4]
  wire [2:0] _T_6152; // @[Bitwise.scala 48:55:@4098.4]
  wire [2:0] _GEN_719; // @[Bitwise.scala 48:55:@4099.4]
  wire [3:0] _T_6153; // @[Bitwise.scala 48:55:@4099.4]
  wire [3:0] _GEN_720; // @[Bitwise.scala 48:55:@4100.4]
  wire [4:0] _T_6154; // @[Bitwise.scala 48:55:@4100.4]
  wire [1:0] _T_6155; // @[Bitwise.scala 48:55:@4101.4]
  wire [1:0] _T_6156; // @[Bitwise.scala 48:55:@4102.4]
  wire [1:0] _GEN_721; // @[Bitwise.scala 48:55:@4103.4]
  wire [2:0] _T_6157; // @[Bitwise.scala 48:55:@4103.4]
  wire [2:0] _GEN_722; // @[Bitwise.scala 48:55:@4104.4]
  wire [3:0] _T_6158; // @[Bitwise.scala 48:55:@4104.4]
  wire [1:0] _T_6159; // @[Bitwise.scala 48:55:@4105.4]
  wire [1:0] _T_6160; // @[Bitwise.scala 48:55:@4106.4]
  wire [1:0] _GEN_723; // @[Bitwise.scala 48:55:@4107.4]
  wire [2:0] _T_6161; // @[Bitwise.scala 48:55:@4107.4]
  wire [2:0] _GEN_724; // @[Bitwise.scala 48:55:@4108.4]
  wire [3:0] _T_6162; // @[Bitwise.scala 48:55:@4108.4]
  wire [4:0] _T_6163; // @[Bitwise.scala 48:55:@4109.4]
  wire [5:0] _T_6164; // @[Bitwise.scala 48:55:@4110.4]
  wire [1:0] _T_6165; // @[Bitwise.scala 48:55:@4111.4]
  wire [1:0] _T_6166; // @[Bitwise.scala 48:55:@4112.4]
  wire [1:0] _GEN_725; // @[Bitwise.scala 48:55:@4113.4]
  wire [2:0] _T_6167; // @[Bitwise.scala 48:55:@4113.4]
  wire [2:0] _GEN_726; // @[Bitwise.scala 48:55:@4114.4]
  wire [3:0] _T_6168; // @[Bitwise.scala 48:55:@4114.4]
  wire [1:0] _T_6169; // @[Bitwise.scala 48:55:@4115.4]
  wire [1:0] _T_6170; // @[Bitwise.scala 48:55:@4116.4]
  wire [1:0] _GEN_727; // @[Bitwise.scala 48:55:@4117.4]
  wire [2:0] _T_6171; // @[Bitwise.scala 48:55:@4117.4]
  wire [2:0] _GEN_728; // @[Bitwise.scala 48:55:@4118.4]
  wire [3:0] _T_6172; // @[Bitwise.scala 48:55:@4118.4]
  wire [4:0] _T_6173; // @[Bitwise.scala 48:55:@4119.4]
  wire [1:0] _T_6174; // @[Bitwise.scala 48:55:@4120.4]
  wire [1:0] _T_6175; // @[Bitwise.scala 48:55:@4121.4]
  wire [1:0] _GEN_729; // @[Bitwise.scala 48:55:@4122.4]
  wire [2:0] _T_6176; // @[Bitwise.scala 48:55:@4122.4]
  wire [2:0] _GEN_730; // @[Bitwise.scala 48:55:@4123.4]
  wire [3:0] _T_6177; // @[Bitwise.scala 48:55:@4123.4]
  wire [1:0] _T_6178; // @[Bitwise.scala 48:55:@4124.4]
  wire [1:0] _T_6179; // @[Bitwise.scala 48:55:@4125.4]
  wire [1:0] _GEN_731; // @[Bitwise.scala 48:55:@4126.4]
  wire [2:0] _T_6180; // @[Bitwise.scala 48:55:@4126.4]
  wire [2:0] _GEN_732; // @[Bitwise.scala 48:55:@4127.4]
  wire [3:0] _T_6181; // @[Bitwise.scala 48:55:@4127.4]
  wire [4:0] _T_6182; // @[Bitwise.scala 48:55:@4128.4]
  wire [5:0] _T_6183; // @[Bitwise.scala 48:55:@4129.4]
  wire [6:0] _T_6184; // @[Bitwise.scala 48:55:@4130.4]
  wire [39:0] _T_6248; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4195.4]
  wire  _T_6249; // @[Bitwise.scala 50:65:@4196.4]
  wire  _T_6250; // @[Bitwise.scala 50:65:@4197.4]
  wire  _T_6251; // @[Bitwise.scala 50:65:@4198.4]
  wire  _T_6252; // @[Bitwise.scala 50:65:@4199.4]
  wire  _T_6253; // @[Bitwise.scala 50:65:@4200.4]
  wire  _T_6254; // @[Bitwise.scala 50:65:@4201.4]
  wire  _T_6255; // @[Bitwise.scala 50:65:@4202.4]
  wire  _T_6256; // @[Bitwise.scala 50:65:@4203.4]
  wire  _T_6257; // @[Bitwise.scala 50:65:@4204.4]
  wire  _T_6258; // @[Bitwise.scala 50:65:@4205.4]
  wire  _T_6259; // @[Bitwise.scala 50:65:@4206.4]
  wire  _T_6260; // @[Bitwise.scala 50:65:@4207.4]
  wire  _T_6261; // @[Bitwise.scala 50:65:@4208.4]
  wire  _T_6262; // @[Bitwise.scala 50:65:@4209.4]
  wire  _T_6263; // @[Bitwise.scala 50:65:@4210.4]
  wire  _T_6264; // @[Bitwise.scala 50:65:@4211.4]
  wire  _T_6265; // @[Bitwise.scala 50:65:@4212.4]
  wire  _T_6266; // @[Bitwise.scala 50:65:@4213.4]
  wire  _T_6267; // @[Bitwise.scala 50:65:@4214.4]
  wire  _T_6268; // @[Bitwise.scala 50:65:@4215.4]
  wire  _T_6269; // @[Bitwise.scala 50:65:@4216.4]
  wire  _T_6270; // @[Bitwise.scala 50:65:@4217.4]
  wire  _T_6271; // @[Bitwise.scala 50:65:@4218.4]
  wire  _T_6272; // @[Bitwise.scala 50:65:@4219.4]
  wire  _T_6273; // @[Bitwise.scala 50:65:@4220.4]
  wire  _T_6274; // @[Bitwise.scala 50:65:@4221.4]
  wire  _T_6275; // @[Bitwise.scala 50:65:@4222.4]
  wire  _T_6276; // @[Bitwise.scala 50:65:@4223.4]
  wire  _T_6277; // @[Bitwise.scala 50:65:@4224.4]
  wire  _T_6278; // @[Bitwise.scala 50:65:@4225.4]
  wire  _T_6279; // @[Bitwise.scala 50:65:@4226.4]
  wire  _T_6280; // @[Bitwise.scala 50:65:@4227.4]
  wire  _T_6281; // @[Bitwise.scala 50:65:@4228.4]
  wire  _T_6282; // @[Bitwise.scala 50:65:@4229.4]
  wire  _T_6283; // @[Bitwise.scala 50:65:@4230.4]
  wire  _T_6284; // @[Bitwise.scala 50:65:@4231.4]
  wire  _T_6285; // @[Bitwise.scala 50:65:@4232.4]
  wire  _T_6286; // @[Bitwise.scala 50:65:@4233.4]
  wire  _T_6287; // @[Bitwise.scala 50:65:@4234.4]
  wire  _T_6288; // @[Bitwise.scala 50:65:@4235.4]
  wire [1:0] _T_6289; // @[Bitwise.scala 48:55:@4236.4]
  wire [1:0] _T_6290; // @[Bitwise.scala 48:55:@4237.4]
  wire [1:0] _GEN_733; // @[Bitwise.scala 48:55:@4238.4]
  wire [2:0] _T_6291; // @[Bitwise.scala 48:55:@4238.4]
  wire [2:0] _GEN_734; // @[Bitwise.scala 48:55:@4239.4]
  wire [3:0] _T_6292; // @[Bitwise.scala 48:55:@4239.4]
  wire [1:0] _T_6293; // @[Bitwise.scala 48:55:@4240.4]
  wire [1:0] _T_6294; // @[Bitwise.scala 48:55:@4241.4]
  wire [1:0] _GEN_735; // @[Bitwise.scala 48:55:@4242.4]
  wire [2:0] _T_6295; // @[Bitwise.scala 48:55:@4242.4]
  wire [2:0] _GEN_736; // @[Bitwise.scala 48:55:@4243.4]
  wire [3:0] _T_6296; // @[Bitwise.scala 48:55:@4243.4]
  wire [4:0] _T_6297; // @[Bitwise.scala 48:55:@4244.4]
  wire [1:0] _T_6298; // @[Bitwise.scala 48:55:@4245.4]
  wire [1:0] _T_6299; // @[Bitwise.scala 48:55:@4246.4]
  wire [1:0] _GEN_737; // @[Bitwise.scala 48:55:@4247.4]
  wire [2:0] _T_6300; // @[Bitwise.scala 48:55:@4247.4]
  wire [2:0] _GEN_738; // @[Bitwise.scala 48:55:@4248.4]
  wire [3:0] _T_6301; // @[Bitwise.scala 48:55:@4248.4]
  wire [1:0] _T_6302; // @[Bitwise.scala 48:55:@4249.4]
  wire [1:0] _T_6303; // @[Bitwise.scala 48:55:@4250.4]
  wire [1:0] _GEN_739; // @[Bitwise.scala 48:55:@4251.4]
  wire [2:0] _T_6304; // @[Bitwise.scala 48:55:@4251.4]
  wire [2:0] _GEN_740; // @[Bitwise.scala 48:55:@4252.4]
  wire [3:0] _T_6305; // @[Bitwise.scala 48:55:@4252.4]
  wire [4:0] _T_6306; // @[Bitwise.scala 48:55:@4253.4]
  wire [5:0] _T_6307; // @[Bitwise.scala 48:55:@4254.4]
  wire [1:0] _T_6308; // @[Bitwise.scala 48:55:@4255.4]
  wire [1:0] _T_6309; // @[Bitwise.scala 48:55:@4256.4]
  wire [1:0] _GEN_741; // @[Bitwise.scala 48:55:@4257.4]
  wire [2:0] _T_6310; // @[Bitwise.scala 48:55:@4257.4]
  wire [2:0] _GEN_742; // @[Bitwise.scala 48:55:@4258.4]
  wire [3:0] _T_6311; // @[Bitwise.scala 48:55:@4258.4]
  wire [1:0] _T_6312; // @[Bitwise.scala 48:55:@4259.4]
  wire [1:0] _T_6313; // @[Bitwise.scala 48:55:@4260.4]
  wire [1:0] _GEN_743; // @[Bitwise.scala 48:55:@4261.4]
  wire [2:0] _T_6314; // @[Bitwise.scala 48:55:@4261.4]
  wire [2:0] _GEN_744; // @[Bitwise.scala 48:55:@4262.4]
  wire [3:0] _T_6315; // @[Bitwise.scala 48:55:@4262.4]
  wire [4:0] _T_6316; // @[Bitwise.scala 48:55:@4263.4]
  wire [1:0] _T_6317; // @[Bitwise.scala 48:55:@4264.4]
  wire [1:0] _T_6318; // @[Bitwise.scala 48:55:@4265.4]
  wire [1:0] _GEN_745; // @[Bitwise.scala 48:55:@4266.4]
  wire [2:0] _T_6319; // @[Bitwise.scala 48:55:@4266.4]
  wire [2:0] _GEN_746; // @[Bitwise.scala 48:55:@4267.4]
  wire [3:0] _T_6320; // @[Bitwise.scala 48:55:@4267.4]
  wire [1:0] _T_6321; // @[Bitwise.scala 48:55:@4268.4]
  wire [1:0] _T_6322; // @[Bitwise.scala 48:55:@4269.4]
  wire [1:0] _GEN_747; // @[Bitwise.scala 48:55:@4270.4]
  wire [2:0] _T_6323; // @[Bitwise.scala 48:55:@4270.4]
  wire [2:0] _GEN_748; // @[Bitwise.scala 48:55:@4271.4]
  wire [3:0] _T_6324; // @[Bitwise.scala 48:55:@4271.4]
  wire [4:0] _T_6325; // @[Bitwise.scala 48:55:@4272.4]
  wire [5:0] _T_6326; // @[Bitwise.scala 48:55:@4273.4]
  wire [6:0] _T_6327; // @[Bitwise.scala 48:55:@4274.4]
  wire [40:0] _T_6391; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4339.4]
  wire  _T_6392; // @[Bitwise.scala 50:65:@4340.4]
  wire  _T_6393; // @[Bitwise.scala 50:65:@4341.4]
  wire  _T_6394; // @[Bitwise.scala 50:65:@4342.4]
  wire  _T_6395; // @[Bitwise.scala 50:65:@4343.4]
  wire  _T_6396; // @[Bitwise.scala 50:65:@4344.4]
  wire  _T_6397; // @[Bitwise.scala 50:65:@4345.4]
  wire  _T_6398; // @[Bitwise.scala 50:65:@4346.4]
  wire  _T_6399; // @[Bitwise.scala 50:65:@4347.4]
  wire  _T_6400; // @[Bitwise.scala 50:65:@4348.4]
  wire  _T_6401; // @[Bitwise.scala 50:65:@4349.4]
  wire  _T_6402; // @[Bitwise.scala 50:65:@4350.4]
  wire  _T_6403; // @[Bitwise.scala 50:65:@4351.4]
  wire  _T_6404; // @[Bitwise.scala 50:65:@4352.4]
  wire  _T_6405; // @[Bitwise.scala 50:65:@4353.4]
  wire  _T_6406; // @[Bitwise.scala 50:65:@4354.4]
  wire  _T_6407; // @[Bitwise.scala 50:65:@4355.4]
  wire  _T_6408; // @[Bitwise.scala 50:65:@4356.4]
  wire  _T_6409; // @[Bitwise.scala 50:65:@4357.4]
  wire  _T_6410; // @[Bitwise.scala 50:65:@4358.4]
  wire  _T_6411; // @[Bitwise.scala 50:65:@4359.4]
  wire  _T_6412; // @[Bitwise.scala 50:65:@4360.4]
  wire  _T_6413; // @[Bitwise.scala 50:65:@4361.4]
  wire  _T_6414; // @[Bitwise.scala 50:65:@4362.4]
  wire  _T_6415; // @[Bitwise.scala 50:65:@4363.4]
  wire  _T_6416; // @[Bitwise.scala 50:65:@4364.4]
  wire  _T_6417; // @[Bitwise.scala 50:65:@4365.4]
  wire  _T_6418; // @[Bitwise.scala 50:65:@4366.4]
  wire  _T_6419; // @[Bitwise.scala 50:65:@4367.4]
  wire  _T_6420; // @[Bitwise.scala 50:65:@4368.4]
  wire  _T_6421; // @[Bitwise.scala 50:65:@4369.4]
  wire  _T_6422; // @[Bitwise.scala 50:65:@4370.4]
  wire  _T_6423; // @[Bitwise.scala 50:65:@4371.4]
  wire  _T_6424; // @[Bitwise.scala 50:65:@4372.4]
  wire  _T_6425; // @[Bitwise.scala 50:65:@4373.4]
  wire  _T_6426; // @[Bitwise.scala 50:65:@4374.4]
  wire  _T_6427; // @[Bitwise.scala 50:65:@4375.4]
  wire  _T_6428; // @[Bitwise.scala 50:65:@4376.4]
  wire  _T_6429; // @[Bitwise.scala 50:65:@4377.4]
  wire  _T_6430; // @[Bitwise.scala 50:65:@4378.4]
  wire  _T_6431; // @[Bitwise.scala 50:65:@4379.4]
  wire  _T_6432; // @[Bitwise.scala 50:65:@4380.4]
  wire [1:0] _T_6433; // @[Bitwise.scala 48:55:@4381.4]
  wire [1:0] _T_6434; // @[Bitwise.scala 48:55:@4382.4]
  wire [1:0] _GEN_749; // @[Bitwise.scala 48:55:@4383.4]
  wire [2:0] _T_6435; // @[Bitwise.scala 48:55:@4383.4]
  wire [2:0] _GEN_750; // @[Bitwise.scala 48:55:@4384.4]
  wire [3:0] _T_6436; // @[Bitwise.scala 48:55:@4384.4]
  wire [1:0] _T_6437; // @[Bitwise.scala 48:55:@4385.4]
  wire [1:0] _T_6438; // @[Bitwise.scala 48:55:@4386.4]
  wire [1:0] _GEN_751; // @[Bitwise.scala 48:55:@4387.4]
  wire [2:0] _T_6439; // @[Bitwise.scala 48:55:@4387.4]
  wire [2:0] _GEN_752; // @[Bitwise.scala 48:55:@4388.4]
  wire [3:0] _T_6440; // @[Bitwise.scala 48:55:@4388.4]
  wire [4:0] _T_6441; // @[Bitwise.scala 48:55:@4389.4]
  wire [1:0] _T_6442; // @[Bitwise.scala 48:55:@4390.4]
  wire [1:0] _T_6443; // @[Bitwise.scala 48:55:@4391.4]
  wire [1:0] _GEN_753; // @[Bitwise.scala 48:55:@4392.4]
  wire [2:0] _T_6444; // @[Bitwise.scala 48:55:@4392.4]
  wire [2:0] _GEN_754; // @[Bitwise.scala 48:55:@4393.4]
  wire [3:0] _T_6445; // @[Bitwise.scala 48:55:@4393.4]
  wire [1:0] _T_6446; // @[Bitwise.scala 48:55:@4394.4]
  wire [1:0] _T_6447; // @[Bitwise.scala 48:55:@4395.4]
  wire [1:0] _GEN_755; // @[Bitwise.scala 48:55:@4396.4]
  wire [2:0] _T_6448; // @[Bitwise.scala 48:55:@4396.4]
  wire [2:0] _GEN_756; // @[Bitwise.scala 48:55:@4397.4]
  wire [3:0] _T_6449; // @[Bitwise.scala 48:55:@4397.4]
  wire [4:0] _T_6450; // @[Bitwise.scala 48:55:@4398.4]
  wire [5:0] _T_6451; // @[Bitwise.scala 48:55:@4399.4]
  wire [1:0] _T_6452; // @[Bitwise.scala 48:55:@4400.4]
  wire [1:0] _T_6453; // @[Bitwise.scala 48:55:@4401.4]
  wire [1:0] _GEN_757; // @[Bitwise.scala 48:55:@4402.4]
  wire [2:0] _T_6454; // @[Bitwise.scala 48:55:@4402.4]
  wire [2:0] _GEN_758; // @[Bitwise.scala 48:55:@4403.4]
  wire [3:0] _T_6455; // @[Bitwise.scala 48:55:@4403.4]
  wire [1:0] _T_6456; // @[Bitwise.scala 48:55:@4404.4]
  wire [1:0] _T_6457; // @[Bitwise.scala 48:55:@4405.4]
  wire [1:0] _GEN_759; // @[Bitwise.scala 48:55:@4406.4]
  wire [2:0] _T_6458; // @[Bitwise.scala 48:55:@4406.4]
  wire [2:0] _GEN_760; // @[Bitwise.scala 48:55:@4407.4]
  wire [3:0] _T_6459; // @[Bitwise.scala 48:55:@4407.4]
  wire [4:0] _T_6460; // @[Bitwise.scala 48:55:@4408.4]
  wire [1:0] _T_6461; // @[Bitwise.scala 48:55:@4409.4]
  wire [1:0] _T_6462; // @[Bitwise.scala 48:55:@4410.4]
  wire [1:0] _GEN_761; // @[Bitwise.scala 48:55:@4411.4]
  wire [2:0] _T_6463; // @[Bitwise.scala 48:55:@4411.4]
  wire [2:0] _GEN_762; // @[Bitwise.scala 48:55:@4412.4]
  wire [3:0] _T_6464; // @[Bitwise.scala 48:55:@4412.4]
  wire [1:0] _T_6465; // @[Bitwise.scala 48:55:@4413.4]
  wire [1:0] _GEN_763; // @[Bitwise.scala 48:55:@4414.4]
  wire [2:0] _T_6466; // @[Bitwise.scala 48:55:@4414.4]
  wire [1:0] _T_6467; // @[Bitwise.scala 48:55:@4415.4]
  wire [1:0] _GEN_764; // @[Bitwise.scala 48:55:@4416.4]
  wire [2:0] _T_6468; // @[Bitwise.scala 48:55:@4416.4]
  wire [3:0] _T_6469; // @[Bitwise.scala 48:55:@4417.4]
  wire [4:0] _T_6470; // @[Bitwise.scala 48:55:@4418.4]
  wire [5:0] _T_6471; // @[Bitwise.scala 48:55:@4419.4]
  wire [6:0] _T_6472; // @[Bitwise.scala 48:55:@4420.4]
  wire [41:0] _T_6536; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4485.4]
  wire  _T_6537; // @[Bitwise.scala 50:65:@4486.4]
  wire  _T_6538; // @[Bitwise.scala 50:65:@4487.4]
  wire  _T_6539; // @[Bitwise.scala 50:65:@4488.4]
  wire  _T_6540; // @[Bitwise.scala 50:65:@4489.4]
  wire  _T_6541; // @[Bitwise.scala 50:65:@4490.4]
  wire  _T_6542; // @[Bitwise.scala 50:65:@4491.4]
  wire  _T_6543; // @[Bitwise.scala 50:65:@4492.4]
  wire  _T_6544; // @[Bitwise.scala 50:65:@4493.4]
  wire  _T_6545; // @[Bitwise.scala 50:65:@4494.4]
  wire  _T_6546; // @[Bitwise.scala 50:65:@4495.4]
  wire  _T_6547; // @[Bitwise.scala 50:65:@4496.4]
  wire  _T_6548; // @[Bitwise.scala 50:65:@4497.4]
  wire  _T_6549; // @[Bitwise.scala 50:65:@4498.4]
  wire  _T_6550; // @[Bitwise.scala 50:65:@4499.4]
  wire  _T_6551; // @[Bitwise.scala 50:65:@4500.4]
  wire  _T_6552; // @[Bitwise.scala 50:65:@4501.4]
  wire  _T_6553; // @[Bitwise.scala 50:65:@4502.4]
  wire  _T_6554; // @[Bitwise.scala 50:65:@4503.4]
  wire  _T_6555; // @[Bitwise.scala 50:65:@4504.4]
  wire  _T_6556; // @[Bitwise.scala 50:65:@4505.4]
  wire  _T_6557; // @[Bitwise.scala 50:65:@4506.4]
  wire  _T_6558; // @[Bitwise.scala 50:65:@4507.4]
  wire  _T_6559; // @[Bitwise.scala 50:65:@4508.4]
  wire  _T_6560; // @[Bitwise.scala 50:65:@4509.4]
  wire  _T_6561; // @[Bitwise.scala 50:65:@4510.4]
  wire  _T_6562; // @[Bitwise.scala 50:65:@4511.4]
  wire  _T_6563; // @[Bitwise.scala 50:65:@4512.4]
  wire  _T_6564; // @[Bitwise.scala 50:65:@4513.4]
  wire  _T_6565; // @[Bitwise.scala 50:65:@4514.4]
  wire  _T_6566; // @[Bitwise.scala 50:65:@4515.4]
  wire  _T_6567; // @[Bitwise.scala 50:65:@4516.4]
  wire  _T_6568; // @[Bitwise.scala 50:65:@4517.4]
  wire  _T_6569; // @[Bitwise.scala 50:65:@4518.4]
  wire  _T_6570; // @[Bitwise.scala 50:65:@4519.4]
  wire  _T_6571; // @[Bitwise.scala 50:65:@4520.4]
  wire  _T_6572; // @[Bitwise.scala 50:65:@4521.4]
  wire  _T_6573; // @[Bitwise.scala 50:65:@4522.4]
  wire  _T_6574; // @[Bitwise.scala 50:65:@4523.4]
  wire  _T_6575; // @[Bitwise.scala 50:65:@4524.4]
  wire  _T_6576; // @[Bitwise.scala 50:65:@4525.4]
  wire  _T_6577; // @[Bitwise.scala 50:65:@4526.4]
  wire  _T_6578; // @[Bitwise.scala 50:65:@4527.4]
  wire [1:0] _T_6579; // @[Bitwise.scala 48:55:@4528.4]
  wire [1:0] _T_6580; // @[Bitwise.scala 48:55:@4529.4]
  wire [1:0] _GEN_765; // @[Bitwise.scala 48:55:@4530.4]
  wire [2:0] _T_6581; // @[Bitwise.scala 48:55:@4530.4]
  wire [2:0] _GEN_766; // @[Bitwise.scala 48:55:@4531.4]
  wire [3:0] _T_6582; // @[Bitwise.scala 48:55:@4531.4]
  wire [1:0] _T_6583; // @[Bitwise.scala 48:55:@4532.4]
  wire [1:0] _T_6584; // @[Bitwise.scala 48:55:@4533.4]
  wire [1:0] _GEN_767; // @[Bitwise.scala 48:55:@4534.4]
  wire [2:0] _T_6585; // @[Bitwise.scala 48:55:@4534.4]
  wire [2:0] _GEN_768; // @[Bitwise.scala 48:55:@4535.4]
  wire [3:0] _T_6586; // @[Bitwise.scala 48:55:@4535.4]
  wire [4:0] _T_6587; // @[Bitwise.scala 48:55:@4536.4]
  wire [1:0] _T_6588; // @[Bitwise.scala 48:55:@4537.4]
  wire [1:0] _T_6589; // @[Bitwise.scala 48:55:@4538.4]
  wire [1:0] _GEN_769; // @[Bitwise.scala 48:55:@4539.4]
  wire [2:0] _T_6590; // @[Bitwise.scala 48:55:@4539.4]
  wire [2:0] _GEN_770; // @[Bitwise.scala 48:55:@4540.4]
  wire [3:0] _T_6591; // @[Bitwise.scala 48:55:@4540.4]
  wire [1:0] _T_6592; // @[Bitwise.scala 48:55:@4541.4]
  wire [1:0] _GEN_771; // @[Bitwise.scala 48:55:@4542.4]
  wire [2:0] _T_6593; // @[Bitwise.scala 48:55:@4542.4]
  wire [1:0] _T_6594; // @[Bitwise.scala 48:55:@4543.4]
  wire [1:0] _GEN_772; // @[Bitwise.scala 48:55:@4544.4]
  wire [2:0] _T_6595; // @[Bitwise.scala 48:55:@4544.4]
  wire [3:0] _T_6596; // @[Bitwise.scala 48:55:@4545.4]
  wire [4:0] _T_6597; // @[Bitwise.scala 48:55:@4546.4]
  wire [5:0] _T_6598; // @[Bitwise.scala 48:55:@4547.4]
  wire [1:0] _T_6599; // @[Bitwise.scala 48:55:@4548.4]
  wire [1:0] _T_6600; // @[Bitwise.scala 48:55:@4549.4]
  wire [1:0] _GEN_773; // @[Bitwise.scala 48:55:@4550.4]
  wire [2:0] _T_6601; // @[Bitwise.scala 48:55:@4550.4]
  wire [2:0] _GEN_774; // @[Bitwise.scala 48:55:@4551.4]
  wire [3:0] _T_6602; // @[Bitwise.scala 48:55:@4551.4]
  wire [1:0] _T_6603; // @[Bitwise.scala 48:55:@4552.4]
  wire [1:0] _T_6604; // @[Bitwise.scala 48:55:@4553.4]
  wire [1:0] _GEN_775; // @[Bitwise.scala 48:55:@4554.4]
  wire [2:0] _T_6605; // @[Bitwise.scala 48:55:@4554.4]
  wire [2:0] _GEN_776; // @[Bitwise.scala 48:55:@4555.4]
  wire [3:0] _T_6606; // @[Bitwise.scala 48:55:@4555.4]
  wire [4:0] _T_6607; // @[Bitwise.scala 48:55:@4556.4]
  wire [1:0] _T_6608; // @[Bitwise.scala 48:55:@4557.4]
  wire [1:0] _T_6609; // @[Bitwise.scala 48:55:@4558.4]
  wire [1:0] _GEN_777; // @[Bitwise.scala 48:55:@4559.4]
  wire [2:0] _T_6610; // @[Bitwise.scala 48:55:@4559.4]
  wire [2:0] _GEN_778; // @[Bitwise.scala 48:55:@4560.4]
  wire [3:0] _T_6611; // @[Bitwise.scala 48:55:@4560.4]
  wire [1:0] _T_6612; // @[Bitwise.scala 48:55:@4561.4]
  wire [1:0] _GEN_779; // @[Bitwise.scala 48:55:@4562.4]
  wire [2:0] _T_6613; // @[Bitwise.scala 48:55:@4562.4]
  wire [1:0] _T_6614; // @[Bitwise.scala 48:55:@4563.4]
  wire [1:0] _GEN_780; // @[Bitwise.scala 48:55:@4564.4]
  wire [2:0] _T_6615; // @[Bitwise.scala 48:55:@4564.4]
  wire [3:0] _T_6616; // @[Bitwise.scala 48:55:@4565.4]
  wire [4:0] _T_6617; // @[Bitwise.scala 48:55:@4566.4]
  wire [5:0] _T_6618; // @[Bitwise.scala 48:55:@4567.4]
  wire [6:0] _T_6619; // @[Bitwise.scala 48:55:@4568.4]
  wire [42:0] _T_6683; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4633.4]
  wire  _T_6684; // @[Bitwise.scala 50:65:@4634.4]
  wire  _T_6685; // @[Bitwise.scala 50:65:@4635.4]
  wire  _T_6686; // @[Bitwise.scala 50:65:@4636.4]
  wire  _T_6687; // @[Bitwise.scala 50:65:@4637.4]
  wire  _T_6688; // @[Bitwise.scala 50:65:@4638.4]
  wire  _T_6689; // @[Bitwise.scala 50:65:@4639.4]
  wire  _T_6690; // @[Bitwise.scala 50:65:@4640.4]
  wire  _T_6691; // @[Bitwise.scala 50:65:@4641.4]
  wire  _T_6692; // @[Bitwise.scala 50:65:@4642.4]
  wire  _T_6693; // @[Bitwise.scala 50:65:@4643.4]
  wire  _T_6694; // @[Bitwise.scala 50:65:@4644.4]
  wire  _T_6695; // @[Bitwise.scala 50:65:@4645.4]
  wire  _T_6696; // @[Bitwise.scala 50:65:@4646.4]
  wire  _T_6697; // @[Bitwise.scala 50:65:@4647.4]
  wire  _T_6698; // @[Bitwise.scala 50:65:@4648.4]
  wire  _T_6699; // @[Bitwise.scala 50:65:@4649.4]
  wire  _T_6700; // @[Bitwise.scala 50:65:@4650.4]
  wire  _T_6701; // @[Bitwise.scala 50:65:@4651.4]
  wire  _T_6702; // @[Bitwise.scala 50:65:@4652.4]
  wire  _T_6703; // @[Bitwise.scala 50:65:@4653.4]
  wire  _T_6704; // @[Bitwise.scala 50:65:@4654.4]
  wire  _T_6705; // @[Bitwise.scala 50:65:@4655.4]
  wire  _T_6706; // @[Bitwise.scala 50:65:@4656.4]
  wire  _T_6707; // @[Bitwise.scala 50:65:@4657.4]
  wire  _T_6708; // @[Bitwise.scala 50:65:@4658.4]
  wire  _T_6709; // @[Bitwise.scala 50:65:@4659.4]
  wire  _T_6710; // @[Bitwise.scala 50:65:@4660.4]
  wire  _T_6711; // @[Bitwise.scala 50:65:@4661.4]
  wire  _T_6712; // @[Bitwise.scala 50:65:@4662.4]
  wire  _T_6713; // @[Bitwise.scala 50:65:@4663.4]
  wire  _T_6714; // @[Bitwise.scala 50:65:@4664.4]
  wire  _T_6715; // @[Bitwise.scala 50:65:@4665.4]
  wire  _T_6716; // @[Bitwise.scala 50:65:@4666.4]
  wire  _T_6717; // @[Bitwise.scala 50:65:@4667.4]
  wire  _T_6718; // @[Bitwise.scala 50:65:@4668.4]
  wire  _T_6719; // @[Bitwise.scala 50:65:@4669.4]
  wire  _T_6720; // @[Bitwise.scala 50:65:@4670.4]
  wire  _T_6721; // @[Bitwise.scala 50:65:@4671.4]
  wire  _T_6722; // @[Bitwise.scala 50:65:@4672.4]
  wire  _T_6723; // @[Bitwise.scala 50:65:@4673.4]
  wire  _T_6724; // @[Bitwise.scala 50:65:@4674.4]
  wire  _T_6725; // @[Bitwise.scala 50:65:@4675.4]
  wire  _T_6726; // @[Bitwise.scala 50:65:@4676.4]
  wire [1:0] _T_6727; // @[Bitwise.scala 48:55:@4677.4]
  wire [1:0] _T_6728; // @[Bitwise.scala 48:55:@4678.4]
  wire [1:0] _GEN_781; // @[Bitwise.scala 48:55:@4679.4]
  wire [2:0] _T_6729; // @[Bitwise.scala 48:55:@4679.4]
  wire [2:0] _GEN_782; // @[Bitwise.scala 48:55:@4680.4]
  wire [3:0] _T_6730; // @[Bitwise.scala 48:55:@4680.4]
  wire [1:0] _T_6731; // @[Bitwise.scala 48:55:@4681.4]
  wire [1:0] _T_6732; // @[Bitwise.scala 48:55:@4682.4]
  wire [1:0] _GEN_783; // @[Bitwise.scala 48:55:@4683.4]
  wire [2:0] _T_6733; // @[Bitwise.scala 48:55:@4683.4]
  wire [2:0] _GEN_784; // @[Bitwise.scala 48:55:@4684.4]
  wire [3:0] _T_6734; // @[Bitwise.scala 48:55:@4684.4]
  wire [4:0] _T_6735; // @[Bitwise.scala 48:55:@4685.4]
  wire [1:0] _T_6736; // @[Bitwise.scala 48:55:@4686.4]
  wire [1:0] _T_6737; // @[Bitwise.scala 48:55:@4687.4]
  wire [1:0] _GEN_785; // @[Bitwise.scala 48:55:@4688.4]
  wire [2:0] _T_6738; // @[Bitwise.scala 48:55:@4688.4]
  wire [2:0] _GEN_786; // @[Bitwise.scala 48:55:@4689.4]
  wire [3:0] _T_6739; // @[Bitwise.scala 48:55:@4689.4]
  wire [1:0] _T_6740; // @[Bitwise.scala 48:55:@4690.4]
  wire [1:0] _GEN_787; // @[Bitwise.scala 48:55:@4691.4]
  wire [2:0] _T_6741; // @[Bitwise.scala 48:55:@4691.4]
  wire [1:0] _T_6742; // @[Bitwise.scala 48:55:@4692.4]
  wire [1:0] _GEN_788; // @[Bitwise.scala 48:55:@4693.4]
  wire [2:0] _T_6743; // @[Bitwise.scala 48:55:@4693.4]
  wire [3:0] _T_6744; // @[Bitwise.scala 48:55:@4694.4]
  wire [4:0] _T_6745; // @[Bitwise.scala 48:55:@4695.4]
  wire [5:0] _T_6746; // @[Bitwise.scala 48:55:@4696.4]
  wire [1:0] _T_6747; // @[Bitwise.scala 48:55:@4697.4]
  wire [1:0] _T_6748; // @[Bitwise.scala 48:55:@4698.4]
  wire [1:0] _GEN_789; // @[Bitwise.scala 48:55:@4699.4]
  wire [2:0] _T_6749; // @[Bitwise.scala 48:55:@4699.4]
  wire [2:0] _GEN_790; // @[Bitwise.scala 48:55:@4700.4]
  wire [3:0] _T_6750; // @[Bitwise.scala 48:55:@4700.4]
  wire [1:0] _T_6751; // @[Bitwise.scala 48:55:@4701.4]
  wire [1:0] _GEN_791; // @[Bitwise.scala 48:55:@4702.4]
  wire [2:0] _T_6752; // @[Bitwise.scala 48:55:@4702.4]
  wire [1:0] _T_6753; // @[Bitwise.scala 48:55:@4703.4]
  wire [1:0] _GEN_792; // @[Bitwise.scala 48:55:@4704.4]
  wire [2:0] _T_6754; // @[Bitwise.scala 48:55:@4704.4]
  wire [3:0] _T_6755; // @[Bitwise.scala 48:55:@4705.4]
  wire [4:0] _T_6756; // @[Bitwise.scala 48:55:@4706.4]
  wire [1:0] _T_6757; // @[Bitwise.scala 48:55:@4707.4]
  wire [1:0] _T_6758; // @[Bitwise.scala 48:55:@4708.4]
  wire [1:0] _GEN_793; // @[Bitwise.scala 48:55:@4709.4]
  wire [2:0] _T_6759; // @[Bitwise.scala 48:55:@4709.4]
  wire [2:0] _GEN_794; // @[Bitwise.scala 48:55:@4710.4]
  wire [3:0] _T_6760; // @[Bitwise.scala 48:55:@4710.4]
  wire [1:0] _T_6761; // @[Bitwise.scala 48:55:@4711.4]
  wire [1:0] _GEN_795; // @[Bitwise.scala 48:55:@4712.4]
  wire [2:0] _T_6762; // @[Bitwise.scala 48:55:@4712.4]
  wire [1:0] _T_6763; // @[Bitwise.scala 48:55:@4713.4]
  wire [1:0] _GEN_796; // @[Bitwise.scala 48:55:@4714.4]
  wire [2:0] _T_6764; // @[Bitwise.scala 48:55:@4714.4]
  wire [3:0] _T_6765; // @[Bitwise.scala 48:55:@4715.4]
  wire [4:0] _T_6766; // @[Bitwise.scala 48:55:@4716.4]
  wire [5:0] _T_6767; // @[Bitwise.scala 48:55:@4717.4]
  wire [6:0] _T_6768; // @[Bitwise.scala 48:55:@4718.4]
  wire [43:0] _T_6832; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4783.4]
  wire  _T_6833; // @[Bitwise.scala 50:65:@4784.4]
  wire  _T_6834; // @[Bitwise.scala 50:65:@4785.4]
  wire  _T_6835; // @[Bitwise.scala 50:65:@4786.4]
  wire  _T_6836; // @[Bitwise.scala 50:65:@4787.4]
  wire  _T_6837; // @[Bitwise.scala 50:65:@4788.4]
  wire  _T_6838; // @[Bitwise.scala 50:65:@4789.4]
  wire  _T_6839; // @[Bitwise.scala 50:65:@4790.4]
  wire  _T_6840; // @[Bitwise.scala 50:65:@4791.4]
  wire  _T_6841; // @[Bitwise.scala 50:65:@4792.4]
  wire  _T_6842; // @[Bitwise.scala 50:65:@4793.4]
  wire  _T_6843; // @[Bitwise.scala 50:65:@4794.4]
  wire  _T_6844; // @[Bitwise.scala 50:65:@4795.4]
  wire  _T_6845; // @[Bitwise.scala 50:65:@4796.4]
  wire  _T_6846; // @[Bitwise.scala 50:65:@4797.4]
  wire  _T_6847; // @[Bitwise.scala 50:65:@4798.4]
  wire  _T_6848; // @[Bitwise.scala 50:65:@4799.4]
  wire  _T_6849; // @[Bitwise.scala 50:65:@4800.4]
  wire  _T_6850; // @[Bitwise.scala 50:65:@4801.4]
  wire  _T_6851; // @[Bitwise.scala 50:65:@4802.4]
  wire  _T_6852; // @[Bitwise.scala 50:65:@4803.4]
  wire  _T_6853; // @[Bitwise.scala 50:65:@4804.4]
  wire  _T_6854; // @[Bitwise.scala 50:65:@4805.4]
  wire  _T_6855; // @[Bitwise.scala 50:65:@4806.4]
  wire  _T_6856; // @[Bitwise.scala 50:65:@4807.4]
  wire  _T_6857; // @[Bitwise.scala 50:65:@4808.4]
  wire  _T_6858; // @[Bitwise.scala 50:65:@4809.4]
  wire  _T_6859; // @[Bitwise.scala 50:65:@4810.4]
  wire  _T_6860; // @[Bitwise.scala 50:65:@4811.4]
  wire  _T_6861; // @[Bitwise.scala 50:65:@4812.4]
  wire  _T_6862; // @[Bitwise.scala 50:65:@4813.4]
  wire  _T_6863; // @[Bitwise.scala 50:65:@4814.4]
  wire  _T_6864; // @[Bitwise.scala 50:65:@4815.4]
  wire  _T_6865; // @[Bitwise.scala 50:65:@4816.4]
  wire  _T_6866; // @[Bitwise.scala 50:65:@4817.4]
  wire  _T_6867; // @[Bitwise.scala 50:65:@4818.4]
  wire  _T_6868; // @[Bitwise.scala 50:65:@4819.4]
  wire  _T_6869; // @[Bitwise.scala 50:65:@4820.4]
  wire  _T_6870; // @[Bitwise.scala 50:65:@4821.4]
  wire  _T_6871; // @[Bitwise.scala 50:65:@4822.4]
  wire  _T_6872; // @[Bitwise.scala 50:65:@4823.4]
  wire  _T_6873; // @[Bitwise.scala 50:65:@4824.4]
  wire  _T_6874; // @[Bitwise.scala 50:65:@4825.4]
  wire  _T_6875; // @[Bitwise.scala 50:65:@4826.4]
  wire  _T_6876; // @[Bitwise.scala 50:65:@4827.4]
  wire [1:0] _T_6877; // @[Bitwise.scala 48:55:@4828.4]
  wire [1:0] _T_6878; // @[Bitwise.scala 48:55:@4829.4]
  wire [1:0] _GEN_797; // @[Bitwise.scala 48:55:@4830.4]
  wire [2:0] _T_6879; // @[Bitwise.scala 48:55:@4830.4]
  wire [2:0] _GEN_798; // @[Bitwise.scala 48:55:@4831.4]
  wire [3:0] _T_6880; // @[Bitwise.scala 48:55:@4831.4]
  wire [1:0] _T_6881; // @[Bitwise.scala 48:55:@4832.4]
  wire [1:0] _GEN_799; // @[Bitwise.scala 48:55:@4833.4]
  wire [2:0] _T_6882; // @[Bitwise.scala 48:55:@4833.4]
  wire [1:0] _T_6883; // @[Bitwise.scala 48:55:@4834.4]
  wire [1:0] _GEN_800; // @[Bitwise.scala 48:55:@4835.4]
  wire [2:0] _T_6884; // @[Bitwise.scala 48:55:@4835.4]
  wire [3:0] _T_6885; // @[Bitwise.scala 48:55:@4836.4]
  wire [4:0] _T_6886; // @[Bitwise.scala 48:55:@4837.4]
  wire [1:0] _T_6887; // @[Bitwise.scala 48:55:@4838.4]
  wire [1:0] _T_6888; // @[Bitwise.scala 48:55:@4839.4]
  wire [1:0] _GEN_801; // @[Bitwise.scala 48:55:@4840.4]
  wire [2:0] _T_6889; // @[Bitwise.scala 48:55:@4840.4]
  wire [2:0] _GEN_802; // @[Bitwise.scala 48:55:@4841.4]
  wire [3:0] _T_6890; // @[Bitwise.scala 48:55:@4841.4]
  wire [1:0] _T_6891; // @[Bitwise.scala 48:55:@4842.4]
  wire [1:0] _GEN_803; // @[Bitwise.scala 48:55:@4843.4]
  wire [2:0] _T_6892; // @[Bitwise.scala 48:55:@4843.4]
  wire [1:0] _T_6893; // @[Bitwise.scala 48:55:@4844.4]
  wire [1:0] _GEN_804; // @[Bitwise.scala 48:55:@4845.4]
  wire [2:0] _T_6894; // @[Bitwise.scala 48:55:@4845.4]
  wire [3:0] _T_6895; // @[Bitwise.scala 48:55:@4846.4]
  wire [4:0] _T_6896; // @[Bitwise.scala 48:55:@4847.4]
  wire [5:0] _T_6897; // @[Bitwise.scala 48:55:@4848.4]
  wire [1:0] _T_6898; // @[Bitwise.scala 48:55:@4849.4]
  wire [1:0] _T_6899; // @[Bitwise.scala 48:55:@4850.4]
  wire [1:0] _GEN_805; // @[Bitwise.scala 48:55:@4851.4]
  wire [2:0] _T_6900; // @[Bitwise.scala 48:55:@4851.4]
  wire [2:0] _GEN_806; // @[Bitwise.scala 48:55:@4852.4]
  wire [3:0] _T_6901; // @[Bitwise.scala 48:55:@4852.4]
  wire [1:0] _T_6902; // @[Bitwise.scala 48:55:@4853.4]
  wire [1:0] _GEN_807; // @[Bitwise.scala 48:55:@4854.4]
  wire [2:0] _T_6903; // @[Bitwise.scala 48:55:@4854.4]
  wire [1:0] _T_6904; // @[Bitwise.scala 48:55:@4855.4]
  wire [1:0] _GEN_808; // @[Bitwise.scala 48:55:@4856.4]
  wire [2:0] _T_6905; // @[Bitwise.scala 48:55:@4856.4]
  wire [3:0] _T_6906; // @[Bitwise.scala 48:55:@4857.4]
  wire [4:0] _T_6907; // @[Bitwise.scala 48:55:@4858.4]
  wire [1:0] _T_6908; // @[Bitwise.scala 48:55:@4859.4]
  wire [1:0] _T_6909; // @[Bitwise.scala 48:55:@4860.4]
  wire [1:0] _GEN_809; // @[Bitwise.scala 48:55:@4861.4]
  wire [2:0] _T_6910; // @[Bitwise.scala 48:55:@4861.4]
  wire [2:0] _GEN_810; // @[Bitwise.scala 48:55:@4862.4]
  wire [3:0] _T_6911; // @[Bitwise.scala 48:55:@4862.4]
  wire [1:0] _T_6912; // @[Bitwise.scala 48:55:@4863.4]
  wire [1:0] _GEN_811; // @[Bitwise.scala 48:55:@4864.4]
  wire [2:0] _T_6913; // @[Bitwise.scala 48:55:@4864.4]
  wire [1:0] _T_6914; // @[Bitwise.scala 48:55:@4865.4]
  wire [1:0] _GEN_812; // @[Bitwise.scala 48:55:@4866.4]
  wire [2:0] _T_6915; // @[Bitwise.scala 48:55:@4866.4]
  wire [3:0] _T_6916; // @[Bitwise.scala 48:55:@4867.4]
  wire [4:0] _T_6917; // @[Bitwise.scala 48:55:@4868.4]
  wire [5:0] _T_6918; // @[Bitwise.scala 48:55:@4869.4]
  wire [6:0] _T_6919; // @[Bitwise.scala 48:55:@4870.4]
  wire [44:0] _T_6983; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4935.4]
  wire  _T_6984; // @[Bitwise.scala 50:65:@4936.4]
  wire  _T_6985; // @[Bitwise.scala 50:65:@4937.4]
  wire  _T_6986; // @[Bitwise.scala 50:65:@4938.4]
  wire  _T_6987; // @[Bitwise.scala 50:65:@4939.4]
  wire  _T_6988; // @[Bitwise.scala 50:65:@4940.4]
  wire  _T_6989; // @[Bitwise.scala 50:65:@4941.4]
  wire  _T_6990; // @[Bitwise.scala 50:65:@4942.4]
  wire  _T_6991; // @[Bitwise.scala 50:65:@4943.4]
  wire  _T_6992; // @[Bitwise.scala 50:65:@4944.4]
  wire  _T_6993; // @[Bitwise.scala 50:65:@4945.4]
  wire  _T_6994; // @[Bitwise.scala 50:65:@4946.4]
  wire  _T_6995; // @[Bitwise.scala 50:65:@4947.4]
  wire  _T_6996; // @[Bitwise.scala 50:65:@4948.4]
  wire  _T_6997; // @[Bitwise.scala 50:65:@4949.4]
  wire  _T_6998; // @[Bitwise.scala 50:65:@4950.4]
  wire  _T_6999; // @[Bitwise.scala 50:65:@4951.4]
  wire  _T_7000; // @[Bitwise.scala 50:65:@4952.4]
  wire  _T_7001; // @[Bitwise.scala 50:65:@4953.4]
  wire  _T_7002; // @[Bitwise.scala 50:65:@4954.4]
  wire  _T_7003; // @[Bitwise.scala 50:65:@4955.4]
  wire  _T_7004; // @[Bitwise.scala 50:65:@4956.4]
  wire  _T_7005; // @[Bitwise.scala 50:65:@4957.4]
  wire  _T_7006; // @[Bitwise.scala 50:65:@4958.4]
  wire  _T_7007; // @[Bitwise.scala 50:65:@4959.4]
  wire  _T_7008; // @[Bitwise.scala 50:65:@4960.4]
  wire  _T_7009; // @[Bitwise.scala 50:65:@4961.4]
  wire  _T_7010; // @[Bitwise.scala 50:65:@4962.4]
  wire  _T_7011; // @[Bitwise.scala 50:65:@4963.4]
  wire  _T_7012; // @[Bitwise.scala 50:65:@4964.4]
  wire  _T_7013; // @[Bitwise.scala 50:65:@4965.4]
  wire  _T_7014; // @[Bitwise.scala 50:65:@4966.4]
  wire  _T_7015; // @[Bitwise.scala 50:65:@4967.4]
  wire  _T_7016; // @[Bitwise.scala 50:65:@4968.4]
  wire  _T_7017; // @[Bitwise.scala 50:65:@4969.4]
  wire  _T_7018; // @[Bitwise.scala 50:65:@4970.4]
  wire  _T_7019; // @[Bitwise.scala 50:65:@4971.4]
  wire  _T_7020; // @[Bitwise.scala 50:65:@4972.4]
  wire  _T_7021; // @[Bitwise.scala 50:65:@4973.4]
  wire  _T_7022; // @[Bitwise.scala 50:65:@4974.4]
  wire  _T_7023; // @[Bitwise.scala 50:65:@4975.4]
  wire  _T_7024; // @[Bitwise.scala 50:65:@4976.4]
  wire  _T_7025; // @[Bitwise.scala 50:65:@4977.4]
  wire  _T_7026; // @[Bitwise.scala 50:65:@4978.4]
  wire  _T_7027; // @[Bitwise.scala 50:65:@4979.4]
  wire  _T_7028; // @[Bitwise.scala 50:65:@4980.4]
  wire [1:0] _T_7029; // @[Bitwise.scala 48:55:@4981.4]
  wire [1:0] _T_7030; // @[Bitwise.scala 48:55:@4982.4]
  wire [1:0] _GEN_813; // @[Bitwise.scala 48:55:@4983.4]
  wire [2:0] _T_7031; // @[Bitwise.scala 48:55:@4983.4]
  wire [2:0] _GEN_814; // @[Bitwise.scala 48:55:@4984.4]
  wire [3:0] _T_7032; // @[Bitwise.scala 48:55:@4984.4]
  wire [1:0] _T_7033; // @[Bitwise.scala 48:55:@4985.4]
  wire [1:0] _GEN_815; // @[Bitwise.scala 48:55:@4986.4]
  wire [2:0] _T_7034; // @[Bitwise.scala 48:55:@4986.4]
  wire [1:0] _T_7035; // @[Bitwise.scala 48:55:@4987.4]
  wire [1:0] _GEN_816; // @[Bitwise.scala 48:55:@4988.4]
  wire [2:0] _T_7036; // @[Bitwise.scala 48:55:@4988.4]
  wire [3:0] _T_7037; // @[Bitwise.scala 48:55:@4989.4]
  wire [4:0] _T_7038; // @[Bitwise.scala 48:55:@4990.4]
  wire [1:0] _T_7039; // @[Bitwise.scala 48:55:@4991.4]
  wire [1:0] _T_7040; // @[Bitwise.scala 48:55:@4992.4]
  wire [1:0] _GEN_817; // @[Bitwise.scala 48:55:@4993.4]
  wire [2:0] _T_7041; // @[Bitwise.scala 48:55:@4993.4]
  wire [2:0] _GEN_818; // @[Bitwise.scala 48:55:@4994.4]
  wire [3:0] _T_7042; // @[Bitwise.scala 48:55:@4994.4]
  wire [1:0] _T_7043; // @[Bitwise.scala 48:55:@4995.4]
  wire [1:0] _GEN_819; // @[Bitwise.scala 48:55:@4996.4]
  wire [2:0] _T_7044; // @[Bitwise.scala 48:55:@4996.4]
  wire [1:0] _T_7045; // @[Bitwise.scala 48:55:@4997.4]
  wire [1:0] _GEN_820; // @[Bitwise.scala 48:55:@4998.4]
  wire [2:0] _T_7046; // @[Bitwise.scala 48:55:@4998.4]
  wire [3:0] _T_7047; // @[Bitwise.scala 48:55:@4999.4]
  wire [4:0] _T_7048; // @[Bitwise.scala 48:55:@5000.4]
  wire [5:0] _T_7049; // @[Bitwise.scala 48:55:@5001.4]
  wire [1:0] _T_7050; // @[Bitwise.scala 48:55:@5002.4]
  wire [1:0] _T_7051; // @[Bitwise.scala 48:55:@5003.4]
  wire [1:0] _GEN_821; // @[Bitwise.scala 48:55:@5004.4]
  wire [2:0] _T_7052; // @[Bitwise.scala 48:55:@5004.4]
  wire [2:0] _GEN_822; // @[Bitwise.scala 48:55:@5005.4]
  wire [3:0] _T_7053; // @[Bitwise.scala 48:55:@5005.4]
  wire [1:0] _T_7054; // @[Bitwise.scala 48:55:@5006.4]
  wire [1:0] _GEN_823; // @[Bitwise.scala 48:55:@5007.4]
  wire [2:0] _T_7055; // @[Bitwise.scala 48:55:@5007.4]
  wire [1:0] _T_7056; // @[Bitwise.scala 48:55:@5008.4]
  wire [1:0] _GEN_824; // @[Bitwise.scala 48:55:@5009.4]
  wire [2:0] _T_7057; // @[Bitwise.scala 48:55:@5009.4]
  wire [3:0] _T_7058; // @[Bitwise.scala 48:55:@5010.4]
  wire [4:0] _T_7059; // @[Bitwise.scala 48:55:@5011.4]
  wire [1:0] _T_7060; // @[Bitwise.scala 48:55:@5012.4]
  wire [1:0] _GEN_825; // @[Bitwise.scala 48:55:@5013.4]
  wire [2:0] _T_7061; // @[Bitwise.scala 48:55:@5013.4]
  wire [1:0] _T_7062; // @[Bitwise.scala 48:55:@5014.4]
  wire [1:0] _GEN_826; // @[Bitwise.scala 48:55:@5015.4]
  wire [2:0] _T_7063; // @[Bitwise.scala 48:55:@5015.4]
  wire [3:0] _T_7064; // @[Bitwise.scala 48:55:@5016.4]
  wire [1:0] _T_7065; // @[Bitwise.scala 48:55:@5017.4]
  wire [1:0] _GEN_827; // @[Bitwise.scala 48:55:@5018.4]
  wire [2:0] _T_7066; // @[Bitwise.scala 48:55:@5018.4]
  wire [1:0] _T_7067; // @[Bitwise.scala 48:55:@5019.4]
  wire [1:0] _GEN_828; // @[Bitwise.scala 48:55:@5020.4]
  wire [2:0] _T_7068; // @[Bitwise.scala 48:55:@5020.4]
  wire [3:0] _T_7069; // @[Bitwise.scala 48:55:@5021.4]
  wire [4:0] _T_7070; // @[Bitwise.scala 48:55:@5022.4]
  wire [5:0] _T_7071; // @[Bitwise.scala 48:55:@5023.4]
  wire [6:0] _T_7072; // @[Bitwise.scala 48:55:@5024.4]
  wire [45:0] _T_7136; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5089.4]
  wire  _T_7137; // @[Bitwise.scala 50:65:@5090.4]
  wire  _T_7138; // @[Bitwise.scala 50:65:@5091.4]
  wire  _T_7139; // @[Bitwise.scala 50:65:@5092.4]
  wire  _T_7140; // @[Bitwise.scala 50:65:@5093.4]
  wire  _T_7141; // @[Bitwise.scala 50:65:@5094.4]
  wire  _T_7142; // @[Bitwise.scala 50:65:@5095.4]
  wire  _T_7143; // @[Bitwise.scala 50:65:@5096.4]
  wire  _T_7144; // @[Bitwise.scala 50:65:@5097.4]
  wire  _T_7145; // @[Bitwise.scala 50:65:@5098.4]
  wire  _T_7146; // @[Bitwise.scala 50:65:@5099.4]
  wire  _T_7147; // @[Bitwise.scala 50:65:@5100.4]
  wire  _T_7148; // @[Bitwise.scala 50:65:@5101.4]
  wire  _T_7149; // @[Bitwise.scala 50:65:@5102.4]
  wire  _T_7150; // @[Bitwise.scala 50:65:@5103.4]
  wire  _T_7151; // @[Bitwise.scala 50:65:@5104.4]
  wire  _T_7152; // @[Bitwise.scala 50:65:@5105.4]
  wire  _T_7153; // @[Bitwise.scala 50:65:@5106.4]
  wire  _T_7154; // @[Bitwise.scala 50:65:@5107.4]
  wire  _T_7155; // @[Bitwise.scala 50:65:@5108.4]
  wire  _T_7156; // @[Bitwise.scala 50:65:@5109.4]
  wire  _T_7157; // @[Bitwise.scala 50:65:@5110.4]
  wire  _T_7158; // @[Bitwise.scala 50:65:@5111.4]
  wire  _T_7159; // @[Bitwise.scala 50:65:@5112.4]
  wire  _T_7160; // @[Bitwise.scala 50:65:@5113.4]
  wire  _T_7161; // @[Bitwise.scala 50:65:@5114.4]
  wire  _T_7162; // @[Bitwise.scala 50:65:@5115.4]
  wire  _T_7163; // @[Bitwise.scala 50:65:@5116.4]
  wire  _T_7164; // @[Bitwise.scala 50:65:@5117.4]
  wire  _T_7165; // @[Bitwise.scala 50:65:@5118.4]
  wire  _T_7166; // @[Bitwise.scala 50:65:@5119.4]
  wire  _T_7167; // @[Bitwise.scala 50:65:@5120.4]
  wire  _T_7168; // @[Bitwise.scala 50:65:@5121.4]
  wire  _T_7169; // @[Bitwise.scala 50:65:@5122.4]
  wire  _T_7170; // @[Bitwise.scala 50:65:@5123.4]
  wire  _T_7171; // @[Bitwise.scala 50:65:@5124.4]
  wire  _T_7172; // @[Bitwise.scala 50:65:@5125.4]
  wire  _T_7173; // @[Bitwise.scala 50:65:@5126.4]
  wire  _T_7174; // @[Bitwise.scala 50:65:@5127.4]
  wire  _T_7175; // @[Bitwise.scala 50:65:@5128.4]
  wire  _T_7176; // @[Bitwise.scala 50:65:@5129.4]
  wire  _T_7177; // @[Bitwise.scala 50:65:@5130.4]
  wire  _T_7178; // @[Bitwise.scala 50:65:@5131.4]
  wire  _T_7179; // @[Bitwise.scala 50:65:@5132.4]
  wire  _T_7180; // @[Bitwise.scala 50:65:@5133.4]
  wire  _T_7181; // @[Bitwise.scala 50:65:@5134.4]
  wire  _T_7182; // @[Bitwise.scala 50:65:@5135.4]
  wire [1:0] _T_7183; // @[Bitwise.scala 48:55:@5136.4]
  wire [1:0] _T_7184; // @[Bitwise.scala 48:55:@5137.4]
  wire [1:0] _GEN_829; // @[Bitwise.scala 48:55:@5138.4]
  wire [2:0] _T_7185; // @[Bitwise.scala 48:55:@5138.4]
  wire [2:0] _GEN_830; // @[Bitwise.scala 48:55:@5139.4]
  wire [3:0] _T_7186; // @[Bitwise.scala 48:55:@5139.4]
  wire [1:0] _T_7187; // @[Bitwise.scala 48:55:@5140.4]
  wire [1:0] _GEN_831; // @[Bitwise.scala 48:55:@5141.4]
  wire [2:0] _T_7188; // @[Bitwise.scala 48:55:@5141.4]
  wire [1:0] _T_7189; // @[Bitwise.scala 48:55:@5142.4]
  wire [1:0] _GEN_832; // @[Bitwise.scala 48:55:@5143.4]
  wire [2:0] _T_7190; // @[Bitwise.scala 48:55:@5143.4]
  wire [3:0] _T_7191; // @[Bitwise.scala 48:55:@5144.4]
  wire [4:0] _T_7192; // @[Bitwise.scala 48:55:@5145.4]
  wire [1:0] _T_7193; // @[Bitwise.scala 48:55:@5146.4]
  wire [1:0] _GEN_833; // @[Bitwise.scala 48:55:@5147.4]
  wire [2:0] _T_7194; // @[Bitwise.scala 48:55:@5147.4]
  wire [1:0] _T_7195; // @[Bitwise.scala 48:55:@5148.4]
  wire [1:0] _GEN_834; // @[Bitwise.scala 48:55:@5149.4]
  wire [2:0] _T_7196; // @[Bitwise.scala 48:55:@5149.4]
  wire [3:0] _T_7197; // @[Bitwise.scala 48:55:@5150.4]
  wire [1:0] _T_7198; // @[Bitwise.scala 48:55:@5151.4]
  wire [1:0] _GEN_835; // @[Bitwise.scala 48:55:@5152.4]
  wire [2:0] _T_7199; // @[Bitwise.scala 48:55:@5152.4]
  wire [1:0] _T_7200; // @[Bitwise.scala 48:55:@5153.4]
  wire [1:0] _GEN_836; // @[Bitwise.scala 48:55:@5154.4]
  wire [2:0] _T_7201; // @[Bitwise.scala 48:55:@5154.4]
  wire [3:0] _T_7202; // @[Bitwise.scala 48:55:@5155.4]
  wire [4:0] _T_7203; // @[Bitwise.scala 48:55:@5156.4]
  wire [5:0] _T_7204; // @[Bitwise.scala 48:55:@5157.4]
  wire [1:0] _T_7205; // @[Bitwise.scala 48:55:@5158.4]
  wire [1:0] _T_7206; // @[Bitwise.scala 48:55:@5159.4]
  wire [1:0] _GEN_837; // @[Bitwise.scala 48:55:@5160.4]
  wire [2:0] _T_7207; // @[Bitwise.scala 48:55:@5160.4]
  wire [2:0] _GEN_838; // @[Bitwise.scala 48:55:@5161.4]
  wire [3:0] _T_7208; // @[Bitwise.scala 48:55:@5161.4]
  wire [1:0] _T_7209; // @[Bitwise.scala 48:55:@5162.4]
  wire [1:0] _GEN_839; // @[Bitwise.scala 48:55:@5163.4]
  wire [2:0] _T_7210; // @[Bitwise.scala 48:55:@5163.4]
  wire [1:0] _T_7211; // @[Bitwise.scala 48:55:@5164.4]
  wire [1:0] _GEN_840; // @[Bitwise.scala 48:55:@5165.4]
  wire [2:0] _T_7212; // @[Bitwise.scala 48:55:@5165.4]
  wire [3:0] _T_7213; // @[Bitwise.scala 48:55:@5166.4]
  wire [4:0] _T_7214; // @[Bitwise.scala 48:55:@5167.4]
  wire [1:0] _T_7215; // @[Bitwise.scala 48:55:@5168.4]
  wire [1:0] _GEN_841; // @[Bitwise.scala 48:55:@5169.4]
  wire [2:0] _T_7216; // @[Bitwise.scala 48:55:@5169.4]
  wire [1:0] _T_7217; // @[Bitwise.scala 48:55:@5170.4]
  wire [1:0] _GEN_842; // @[Bitwise.scala 48:55:@5171.4]
  wire [2:0] _T_7218; // @[Bitwise.scala 48:55:@5171.4]
  wire [3:0] _T_7219; // @[Bitwise.scala 48:55:@5172.4]
  wire [1:0] _T_7220; // @[Bitwise.scala 48:55:@5173.4]
  wire [1:0] _GEN_843; // @[Bitwise.scala 48:55:@5174.4]
  wire [2:0] _T_7221; // @[Bitwise.scala 48:55:@5174.4]
  wire [1:0] _T_7222; // @[Bitwise.scala 48:55:@5175.4]
  wire [1:0] _GEN_844; // @[Bitwise.scala 48:55:@5176.4]
  wire [2:0] _T_7223; // @[Bitwise.scala 48:55:@5176.4]
  wire [3:0] _T_7224; // @[Bitwise.scala 48:55:@5177.4]
  wire [4:0] _T_7225; // @[Bitwise.scala 48:55:@5178.4]
  wire [5:0] _T_7226; // @[Bitwise.scala 48:55:@5179.4]
  wire [6:0] _T_7227; // @[Bitwise.scala 48:55:@5180.4]
  wire [46:0] _T_7291; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5245.4]
  wire  _T_7292; // @[Bitwise.scala 50:65:@5246.4]
  wire  _T_7293; // @[Bitwise.scala 50:65:@5247.4]
  wire  _T_7294; // @[Bitwise.scala 50:65:@5248.4]
  wire  _T_7295; // @[Bitwise.scala 50:65:@5249.4]
  wire  _T_7296; // @[Bitwise.scala 50:65:@5250.4]
  wire  _T_7297; // @[Bitwise.scala 50:65:@5251.4]
  wire  _T_7298; // @[Bitwise.scala 50:65:@5252.4]
  wire  _T_7299; // @[Bitwise.scala 50:65:@5253.4]
  wire  _T_7300; // @[Bitwise.scala 50:65:@5254.4]
  wire  _T_7301; // @[Bitwise.scala 50:65:@5255.4]
  wire  _T_7302; // @[Bitwise.scala 50:65:@5256.4]
  wire  _T_7303; // @[Bitwise.scala 50:65:@5257.4]
  wire  _T_7304; // @[Bitwise.scala 50:65:@5258.4]
  wire  _T_7305; // @[Bitwise.scala 50:65:@5259.4]
  wire  _T_7306; // @[Bitwise.scala 50:65:@5260.4]
  wire  _T_7307; // @[Bitwise.scala 50:65:@5261.4]
  wire  _T_7308; // @[Bitwise.scala 50:65:@5262.4]
  wire  _T_7309; // @[Bitwise.scala 50:65:@5263.4]
  wire  _T_7310; // @[Bitwise.scala 50:65:@5264.4]
  wire  _T_7311; // @[Bitwise.scala 50:65:@5265.4]
  wire  _T_7312; // @[Bitwise.scala 50:65:@5266.4]
  wire  _T_7313; // @[Bitwise.scala 50:65:@5267.4]
  wire  _T_7314; // @[Bitwise.scala 50:65:@5268.4]
  wire  _T_7315; // @[Bitwise.scala 50:65:@5269.4]
  wire  _T_7316; // @[Bitwise.scala 50:65:@5270.4]
  wire  _T_7317; // @[Bitwise.scala 50:65:@5271.4]
  wire  _T_7318; // @[Bitwise.scala 50:65:@5272.4]
  wire  _T_7319; // @[Bitwise.scala 50:65:@5273.4]
  wire  _T_7320; // @[Bitwise.scala 50:65:@5274.4]
  wire  _T_7321; // @[Bitwise.scala 50:65:@5275.4]
  wire  _T_7322; // @[Bitwise.scala 50:65:@5276.4]
  wire  _T_7323; // @[Bitwise.scala 50:65:@5277.4]
  wire  _T_7324; // @[Bitwise.scala 50:65:@5278.4]
  wire  _T_7325; // @[Bitwise.scala 50:65:@5279.4]
  wire  _T_7326; // @[Bitwise.scala 50:65:@5280.4]
  wire  _T_7327; // @[Bitwise.scala 50:65:@5281.4]
  wire  _T_7328; // @[Bitwise.scala 50:65:@5282.4]
  wire  _T_7329; // @[Bitwise.scala 50:65:@5283.4]
  wire  _T_7330; // @[Bitwise.scala 50:65:@5284.4]
  wire  _T_7331; // @[Bitwise.scala 50:65:@5285.4]
  wire  _T_7332; // @[Bitwise.scala 50:65:@5286.4]
  wire  _T_7333; // @[Bitwise.scala 50:65:@5287.4]
  wire  _T_7334; // @[Bitwise.scala 50:65:@5288.4]
  wire  _T_7335; // @[Bitwise.scala 50:65:@5289.4]
  wire  _T_7336; // @[Bitwise.scala 50:65:@5290.4]
  wire  _T_7337; // @[Bitwise.scala 50:65:@5291.4]
  wire  _T_7338; // @[Bitwise.scala 50:65:@5292.4]
  wire [1:0] _T_7339; // @[Bitwise.scala 48:55:@5293.4]
  wire [1:0] _T_7340; // @[Bitwise.scala 48:55:@5294.4]
  wire [1:0] _GEN_845; // @[Bitwise.scala 48:55:@5295.4]
  wire [2:0] _T_7341; // @[Bitwise.scala 48:55:@5295.4]
  wire [2:0] _GEN_846; // @[Bitwise.scala 48:55:@5296.4]
  wire [3:0] _T_7342; // @[Bitwise.scala 48:55:@5296.4]
  wire [1:0] _T_7343; // @[Bitwise.scala 48:55:@5297.4]
  wire [1:0] _GEN_847; // @[Bitwise.scala 48:55:@5298.4]
  wire [2:0] _T_7344; // @[Bitwise.scala 48:55:@5298.4]
  wire [1:0] _T_7345; // @[Bitwise.scala 48:55:@5299.4]
  wire [1:0] _GEN_848; // @[Bitwise.scala 48:55:@5300.4]
  wire [2:0] _T_7346; // @[Bitwise.scala 48:55:@5300.4]
  wire [3:0] _T_7347; // @[Bitwise.scala 48:55:@5301.4]
  wire [4:0] _T_7348; // @[Bitwise.scala 48:55:@5302.4]
  wire [1:0] _T_7349; // @[Bitwise.scala 48:55:@5303.4]
  wire [1:0] _GEN_849; // @[Bitwise.scala 48:55:@5304.4]
  wire [2:0] _T_7350; // @[Bitwise.scala 48:55:@5304.4]
  wire [1:0] _T_7351; // @[Bitwise.scala 48:55:@5305.4]
  wire [1:0] _GEN_850; // @[Bitwise.scala 48:55:@5306.4]
  wire [2:0] _T_7352; // @[Bitwise.scala 48:55:@5306.4]
  wire [3:0] _T_7353; // @[Bitwise.scala 48:55:@5307.4]
  wire [1:0] _T_7354; // @[Bitwise.scala 48:55:@5308.4]
  wire [1:0] _GEN_851; // @[Bitwise.scala 48:55:@5309.4]
  wire [2:0] _T_7355; // @[Bitwise.scala 48:55:@5309.4]
  wire [1:0] _T_7356; // @[Bitwise.scala 48:55:@5310.4]
  wire [1:0] _GEN_852; // @[Bitwise.scala 48:55:@5311.4]
  wire [2:0] _T_7357; // @[Bitwise.scala 48:55:@5311.4]
  wire [3:0] _T_7358; // @[Bitwise.scala 48:55:@5312.4]
  wire [4:0] _T_7359; // @[Bitwise.scala 48:55:@5313.4]
  wire [5:0] _T_7360; // @[Bitwise.scala 48:55:@5314.4]
  wire [1:0] _T_7361; // @[Bitwise.scala 48:55:@5315.4]
  wire [1:0] _GEN_853; // @[Bitwise.scala 48:55:@5316.4]
  wire [2:0] _T_7362; // @[Bitwise.scala 48:55:@5316.4]
  wire [1:0] _T_7363; // @[Bitwise.scala 48:55:@5317.4]
  wire [1:0] _GEN_854; // @[Bitwise.scala 48:55:@5318.4]
  wire [2:0] _T_7364; // @[Bitwise.scala 48:55:@5318.4]
  wire [3:0] _T_7365; // @[Bitwise.scala 48:55:@5319.4]
  wire [1:0] _T_7366; // @[Bitwise.scala 48:55:@5320.4]
  wire [1:0] _GEN_855; // @[Bitwise.scala 48:55:@5321.4]
  wire [2:0] _T_7367; // @[Bitwise.scala 48:55:@5321.4]
  wire [1:0] _T_7368; // @[Bitwise.scala 48:55:@5322.4]
  wire [1:0] _GEN_856; // @[Bitwise.scala 48:55:@5323.4]
  wire [2:0] _T_7369; // @[Bitwise.scala 48:55:@5323.4]
  wire [3:0] _T_7370; // @[Bitwise.scala 48:55:@5324.4]
  wire [4:0] _T_7371; // @[Bitwise.scala 48:55:@5325.4]
  wire [1:0] _T_7372; // @[Bitwise.scala 48:55:@5326.4]
  wire [1:0] _GEN_857; // @[Bitwise.scala 48:55:@5327.4]
  wire [2:0] _T_7373; // @[Bitwise.scala 48:55:@5327.4]
  wire [1:0] _T_7374; // @[Bitwise.scala 48:55:@5328.4]
  wire [1:0] _GEN_858; // @[Bitwise.scala 48:55:@5329.4]
  wire [2:0] _T_7375; // @[Bitwise.scala 48:55:@5329.4]
  wire [3:0] _T_7376; // @[Bitwise.scala 48:55:@5330.4]
  wire [1:0] _T_7377; // @[Bitwise.scala 48:55:@5331.4]
  wire [1:0] _GEN_859; // @[Bitwise.scala 48:55:@5332.4]
  wire [2:0] _T_7378; // @[Bitwise.scala 48:55:@5332.4]
  wire [1:0] _T_7379; // @[Bitwise.scala 48:55:@5333.4]
  wire [1:0] _GEN_860; // @[Bitwise.scala 48:55:@5334.4]
  wire [2:0] _T_7380; // @[Bitwise.scala 48:55:@5334.4]
  wire [3:0] _T_7381; // @[Bitwise.scala 48:55:@5335.4]
  wire [4:0] _T_7382; // @[Bitwise.scala 48:55:@5336.4]
  wire [5:0] _T_7383; // @[Bitwise.scala 48:55:@5337.4]
  wire [6:0] _T_7384; // @[Bitwise.scala 48:55:@5338.4]
  wire [47:0] _T_7448; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5403.4]
  wire  _T_7449; // @[Bitwise.scala 50:65:@5404.4]
  wire  _T_7450; // @[Bitwise.scala 50:65:@5405.4]
  wire  _T_7451; // @[Bitwise.scala 50:65:@5406.4]
  wire  _T_7452; // @[Bitwise.scala 50:65:@5407.4]
  wire  _T_7453; // @[Bitwise.scala 50:65:@5408.4]
  wire  _T_7454; // @[Bitwise.scala 50:65:@5409.4]
  wire  _T_7455; // @[Bitwise.scala 50:65:@5410.4]
  wire  _T_7456; // @[Bitwise.scala 50:65:@5411.4]
  wire  _T_7457; // @[Bitwise.scala 50:65:@5412.4]
  wire  _T_7458; // @[Bitwise.scala 50:65:@5413.4]
  wire  _T_7459; // @[Bitwise.scala 50:65:@5414.4]
  wire  _T_7460; // @[Bitwise.scala 50:65:@5415.4]
  wire  _T_7461; // @[Bitwise.scala 50:65:@5416.4]
  wire  _T_7462; // @[Bitwise.scala 50:65:@5417.4]
  wire  _T_7463; // @[Bitwise.scala 50:65:@5418.4]
  wire  _T_7464; // @[Bitwise.scala 50:65:@5419.4]
  wire  _T_7465; // @[Bitwise.scala 50:65:@5420.4]
  wire  _T_7466; // @[Bitwise.scala 50:65:@5421.4]
  wire  _T_7467; // @[Bitwise.scala 50:65:@5422.4]
  wire  _T_7468; // @[Bitwise.scala 50:65:@5423.4]
  wire  _T_7469; // @[Bitwise.scala 50:65:@5424.4]
  wire  _T_7470; // @[Bitwise.scala 50:65:@5425.4]
  wire  _T_7471; // @[Bitwise.scala 50:65:@5426.4]
  wire  _T_7472; // @[Bitwise.scala 50:65:@5427.4]
  wire  _T_7473; // @[Bitwise.scala 50:65:@5428.4]
  wire  _T_7474; // @[Bitwise.scala 50:65:@5429.4]
  wire  _T_7475; // @[Bitwise.scala 50:65:@5430.4]
  wire  _T_7476; // @[Bitwise.scala 50:65:@5431.4]
  wire  _T_7477; // @[Bitwise.scala 50:65:@5432.4]
  wire  _T_7478; // @[Bitwise.scala 50:65:@5433.4]
  wire  _T_7479; // @[Bitwise.scala 50:65:@5434.4]
  wire  _T_7480; // @[Bitwise.scala 50:65:@5435.4]
  wire  _T_7481; // @[Bitwise.scala 50:65:@5436.4]
  wire  _T_7482; // @[Bitwise.scala 50:65:@5437.4]
  wire  _T_7483; // @[Bitwise.scala 50:65:@5438.4]
  wire  _T_7484; // @[Bitwise.scala 50:65:@5439.4]
  wire  _T_7485; // @[Bitwise.scala 50:65:@5440.4]
  wire  _T_7486; // @[Bitwise.scala 50:65:@5441.4]
  wire  _T_7487; // @[Bitwise.scala 50:65:@5442.4]
  wire  _T_7488; // @[Bitwise.scala 50:65:@5443.4]
  wire  _T_7489; // @[Bitwise.scala 50:65:@5444.4]
  wire  _T_7490; // @[Bitwise.scala 50:65:@5445.4]
  wire  _T_7491; // @[Bitwise.scala 50:65:@5446.4]
  wire  _T_7492; // @[Bitwise.scala 50:65:@5447.4]
  wire  _T_7493; // @[Bitwise.scala 50:65:@5448.4]
  wire  _T_7494; // @[Bitwise.scala 50:65:@5449.4]
  wire  _T_7495; // @[Bitwise.scala 50:65:@5450.4]
  wire  _T_7496; // @[Bitwise.scala 50:65:@5451.4]
  wire [1:0] _T_7497; // @[Bitwise.scala 48:55:@5452.4]
  wire [1:0] _GEN_861; // @[Bitwise.scala 48:55:@5453.4]
  wire [2:0] _T_7498; // @[Bitwise.scala 48:55:@5453.4]
  wire [1:0] _T_7499; // @[Bitwise.scala 48:55:@5454.4]
  wire [1:0] _GEN_862; // @[Bitwise.scala 48:55:@5455.4]
  wire [2:0] _T_7500; // @[Bitwise.scala 48:55:@5455.4]
  wire [3:0] _T_7501; // @[Bitwise.scala 48:55:@5456.4]
  wire [1:0] _T_7502; // @[Bitwise.scala 48:55:@5457.4]
  wire [1:0] _GEN_863; // @[Bitwise.scala 48:55:@5458.4]
  wire [2:0] _T_7503; // @[Bitwise.scala 48:55:@5458.4]
  wire [1:0] _T_7504; // @[Bitwise.scala 48:55:@5459.4]
  wire [1:0] _GEN_864; // @[Bitwise.scala 48:55:@5460.4]
  wire [2:0] _T_7505; // @[Bitwise.scala 48:55:@5460.4]
  wire [3:0] _T_7506; // @[Bitwise.scala 48:55:@5461.4]
  wire [4:0] _T_7507; // @[Bitwise.scala 48:55:@5462.4]
  wire [1:0] _T_7508; // @[Bitwise.scala 48:55:@5463.4]
  wire [1:0] _GEN_865; // @[Bitwise.scala 48:55:@5464.4]
  wire [2:0] _T_7509; // @[Bitwise.scala 48:55:@5464.4]
  wire [1:0] _T_7510; // @[Bitwise.scala 48:55:@5465.4]
  wire [1:0] _GEN_866; // @[Bitwise.scala 48:55:@5466.4]
  wire [2:0] _T_7511; // @[Bitwise.scala 48:55:@5466.4]
  wire [3:0] _T_7512; // @[Bitwise.scala 48:55:@5467.4]
  wire [1:0] _T_7513; // @[Bitwise.scala 48:55:@5468.4]
  wire [1:0] _GEN_867; // @[Bitwise.scala 48:55:@5469.4]
  wire [2:0] _T_7514; // @[Bitwise.scala 48:55:@5469.4]
  wire [1:0] _T_7515; // @[Bitwise.scala 48:55:@5470.4]
  wire [1:0] _GEN_868; // @[Bitwise.scala 48:55:@5471.4]
  wire [2:0] _T_7516; // @[Bitwise.scala 48:55:@5471.4]
  wire [3:0] _T_7517; // @[Bitwise.scala 48:55:@5472.4]
  wire [4:0] _T_7518; // @[Bitwise.scala 48:55:@5473.4]
  wire [5:0] _T_7519; // @[Bitwise.scala 48:55:@5474.4]
  wire [1:0] _T_7520; // @[Bitwise.scala 48:55:@5475.4]
  wire [1:0] _GEN_869; // @[Bitwise.scala 48:55:@5476.4]
  wire [2:0] _T_7521; // @[Bitwise.scala 48:55:@5476.4]
  wire [1:0] _T_7522; // @[Bitwise.scala 48:55:@5477.4]
  wire [1:0] _GEN_870; // @[Bitwise.scala 48:55:@5478.4]
  wire [2:0] _T_7523; // @[Bitwise.scala 48:55:@5478.4]
  wire [3:0] _T_7524; // @[Bitwise.scala 48:55:@5479.4]
  wire [1:0] _T_7525; // @[Bitwise.scala 48:55:@5480.4]
  wire [1:0] _GEN_871; // @[Bitwise.scala 48:55:@5481.4]
  wire [2:0] _T_7526; // @[Bitwise.scala 48:55:@5481.4]
  wire [1:0] _T_7527; // @[Bitwise.scala 48:55:@5482.4]
  wire [1:0] _GEN_872; // @[Bitwise.scala 48:55:@5483.4]
  wire [2:0] _T_7528; // @[Bitwise.scala 48:55:@5483.4]
  wire [3:0] _T_7529; // @[Bitwise.scala 48:55:@5484.4]
  wire [4:0] _T_7530; // @[Bitwise.scala 48:55:@5485.4]
  wire [1:0] _T_7531; // @[Bitwise.scala 48:55:@5486.4]
  wire [1:0] _GEN_873; // @[Bitwise.scala 48:55:@5487.4]
  wire [2:0] _T_7532; // @[Bitwise.scala 48:55:@5487.4]
  wire [1:0] _T_7533; // @[Bitwise.scala 48:55:@5488.4]
  wire [1:0] _GEN_874; // @[Bitwise.scala 48:55:@5489.4]
  wire [2:0] _T_7534; // @[Bitwise.scala 48:55:@5489.4]
  wire [3:0] _T_7535; // @[Bitwise.scala 48:55:@5490.4]
  wire [1:0] _T_7536; // @[Bitwise.scala 48:55:@5491.4]
  wire [1:0] _GEN_875; // @[Bitwise.scala 48:55:@5492.4]
  wire [2:0] _T_7537; // @[Bitwise.scala 48:55:@5492.4]
  wire [1:0] _T_7538; // @[Bitwise.scala 48:55:@5493.4]
  wire [1:0] _GEN_876; // @[Bitwise.scala 48:55:@5494.4]
  wire [2:0] _T_7539; // @[Bitwise.scala 48:55:@5494.4]
  wire [3:0] _T_7540; // @[Bitwise.scala 48:55:@5495.4]
  wire [4:0] _T_7541; // @[Bitwise.scala 48:55:@5496.4]
  wire [5:0] _T_7542; // @[Bitwise.scala 48:55:@5497.4]
  wire [6:0] _T_7543; // @[Bitwise.scala 48:55:@5498.4]
  wire [48:0] _T_7607; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5563.4]
  wire  _T_7608; // @[Bitwise.scala 50:65:@5564.4]
  wire  _T_7609; // @[Bitwise.scala 50:65:@5565.4]
  wire  _T_7610; // @[Bitwise.scala 50:65:@5566.4]
  wire  _T_7611; // @[Bitwise.scala 50:65:@5567.4]
  wire  _T_7612; // @[Bitwise.scala 50:65:@5568.4]
  wire  _T_7613; // @[Bitwise.scala 50:65:@5569.4]
  wire  _T_7614; // @[Bitwise.scala 50:65:@5570.4]
  wire  _T_7615; // @[Bitwise.scala 50:65:@5571.4]
  wire  _T_7616; // @[Bitwise.scala 50:65:@5572.4]
  wire  _T_7617; // @[Bitwise.scala 50:65:@5573.4]
  wire  _T_7618; // @[Bitwise.scala 50:65:@5574.4]
  wire  _T_7619; // @[Bitwise.scala 50:65:@5575.4]
  wire  _T_7620; // @[Bitwise.scala 50:65:@5576.4]
  wire  _T_7621; // @[Bitwise.scala 50:65:@5577.4]
  wire  _T_7622; // @[Bitwise.scala 50:65:@5578.4]
  wire  _T_7623; // @[Bitwise.scala 50:65:@5579.4]
  wire  _T_7624; // @[Bitwise.scala 50:65:@5580.4]
  wire  _T_7625; // @[Bitwise.scala 50:65:@5581.4]
  wire  _T_7626; // @[Bitwise.scala 50:65:@5582.4]
  wire  _T_7627; // @[Bitwise.scala 50:65:@5583.4]
  wire  _T_7628; // @[Bitwise.scala 50:65:@5584.4]
  wire  _T_7629; // @[Bitwise.scala 50:65:@5585.4]
  wire  _T_7630; // @[Bitwise.scala 50:65:@5586.4]
  wire  _T_7631; // @[Bitwise.scala 50:65:@5587.4]
  wire  _T_7632; // @[Bitwise.scala 50:65:@5588.4]
  wire  _T_7633; // @[Bitwise.scala 50:65:@5589.4]
  wire  _T_7634; // @[Bitwise.scala 50:65:@5590.4]
  wire  _T_7635; // @[Bitwise.scala 50:65:@5591.4]
  wire  _T_7636; // @[Bitwise.scala 50:65:@5592.4]
  wire  _T_7637; // @[Bitwise.scala 50:65:@5593.4]
  wire  _T_7638; // @[Bitwise.scala 50:65:@5594.4]
  wire  _T_7639; // @[Bitwise.scala 50:65:@5595.4]
  wire  _T_7640; // @[Bitwise.scala 50:65:@5596.4]
  wire  _T_7641; // @[Bitwise.scala 50:65:@5597.4]
  wire  _T_7642; // @[Bitwise.scala 50:65:@5598.4]
  wire  _T_7643; // @[Bitwise.scala 50:65:@5599.4]
  wire  _T_7644; // @[Bitwise.scala 50:65:@5600.4]
  wire  _T_7645; // @[Bitwise.scala 50:65:@5601.4]
  wire  _T_7646; // @[Bitwise.scala 50:65:@5602.4]
  wire  _T_7647; // @[Bitwise.scala 50:65:@5603.4]
  wire  _T_7648; // @[Bitwise.scala 50:65:@5604.4]
  wire  _T_7649; // @[Bitwise.scala 50:65:@5605.4]
  wire  _T_7650; // @[Bitwise.scala 50:65:@5606.4]
  wire  _T_7651; // @[Bitwise.scala 50:65:@5607.4]
  wire  _T_7652; // @[Bitwise.scala 50:65:@5608.4]
  wire  _T_7653; // @[Bitwise.scala 50:65:@5609.4]
  wire  _T_7654; // @[Bitwise.scala 50:65:@5610.4]
  wire  _T_7655; // @[Bitwise.scala 50:65:@5611.4]
  wire  _T_7656; // @[Bitwise.scala 50:65:@5612.4]
  wire [1:0] _T_7657; // @[Bitwise.scala 48:55:@5613.4]
  wire [1:0] _GEN_877; // @[Bitwise.scala 48:55:@5614.4]
  wire [2:0] _T_7658; // @[Bitwise.scala 48:55:@5614.4]
  wire [1:0] _T_7659; // @[Bitwise.scala 48:55:@5615.4]
  wire [1:0] _GEN_878; // @[Bitwise.scala 48:55:@5616.4]
  wire [2:0] _T_7660; // @[Bitwise.scala 48:55:@5616.4]
  wire [3:0] _T_7661; // @[Bitwise.scala 48:55:@5617.4]
  wire [1:0] _T_7662; // @[Bitwise.scala 48:55:@5618.4]
  wire [1:0] _GEN_879; // @[Bitwise.scala 48:55:@5619.4]
  wire [2:0] _T_7663; // @[Bitwise.scala 48:55:@5619.4]
  wire [1:0] _T_7664; // @[Bitwise.scala 48:55:@5620.4]
  wire [1:0] _GEN_880; // @[Bitwise.scala 48:55:@5621.4]
  wire [2:0] _T_7665; // @[Bitwise.scala 48:55:@5621.4]
  wire [3:0] _T_7666; // @[Bitwise.scala 48:55:@5622.4]
  wire [4:0] _T_7667; // @[Bitwise.scala 48:55:@5623.4]
  wire [1:0] _T_7668; // @[Bitwise.scala 48:55:@5624.4]
  wire [1:0] _GEN_881; // @[Bitwise.scala 48:55:@5625.4]
  wire [2:0] _T_7669; // @[Bitwise.scala 48:55:@5625.4]
  wire [1:0] _T_7670; // @[Bitwise.scala 48:55:@5626.4]
  wire [1:0] _GEN_882; // @[Bitwise.scala 48:55:@5627.4]
  wire [2:0] _T_7671; // @[Bitwise.scala 48:55:@5627.4]
  wire [3:0] _T_7672; // @[Bitwise.scala 48:55:@5628.4]
  wire [1:0] _T_7673; // @[Bitwise.scala 48:55:@5629.4]
  wire [1:0] _GEN_883; // @[Bitwise.scala 48:55:@5630.4]
  wire [2:0] _T_7674; // @[Bitwise.scala 48:55:@5630.4]
  wire [1:0] _T_7675; // @[Bitwise.scala 48:55:@5631.4]
  wire [1:0] _GEN_884; // @[Bitwise.scala 48:55:@5632.4]
  wire [2:0] _T_7676; // @[Bitwise.scala 48:55:@5632.4]
  wire [3:0] _T_7677; // @[Bitwise.scala 48:55:@5633.4]
  wire [4:0] _T_7678; // @[Bitwise.scala 48:55:@5634.4]
  wire [5:0] _T_7679; // @[Bitwise.scala 48:55:@5635.4]
  wire [1:0] _T_7680; // @[Bitwise.scala 48:55:@5636.4]
  wire [1:0] _GEN_885; // @[Bitwise.scala 48:55:@5637.4]
  wire [2:0] _T_7681; // @[Bitwise.scala 48:55:@5637.4]
  wire [1:0] _T_7682; // @[Bitwise.scala 48:55:@5638.4]
  wire [1:0] _GEN_886; // @[Bitwise.scala 48:55:@5639.4]
  wire [2:0] _T_7683; // @[Bitwise.scala 48:55:@5639.4]
  wire [3:0] _T_7684; // @[Bitwise.scala 48:55:@5640.4]
  wire [1:0] _T_7685; // @[Bitwise.scala 48:55:@5641.4]
  wire [1:0] _GEN_887; // @[Bitwise.scala 48:55:@5642.4]
  wire [2:0] _T_7686; // @[Bitwise.scala 48:55:@5642.4]
  wire [1:0] _T_7687; // @[Bitwise.scala 48:55:@5643.4]
  wire [1:0] _GEN_888; // @[Bitwise.scala 48:55:@5644.4]
  wire [2:0] _T_7688; // @[Bitwise.scala 48:55:@5644.4]
  wire [3:0] _T_7689; // @[Bitwise.scala 48:55:@5645.4]
  wire [4:0] _T_7690; // @[Bitwise.scala 48:55:@5646.4]
  wire [1:0] _T_7691; // @[Bitwise.scala 48:55:@5647.4]
  wire [1:0] _GEN_889; // @[Bitwise.scala 48:55:@5648.4]
  wire [2:0] _T_7692; // @[Bitwise.scala 48:55:@5648.4]
  wire [1:0] _T_7693; // @[Bitwise.scala 48:55:@5649.4]
  wire [1:0] _GEN_890; // @[Bitwise.scala 48:55:@5650.4]
  wire [2:0] _T_7694; // @[Bitwise.scala 48:55:@5650.4]
  wire [3:0] _T_7695; // @[Bitwise.scala 48:55:@5651.4]
  wire [1:0] _T_7696; // @[Bitwise.scala 48:55:@5652.4]
  wire [1:0] _GEN_891; // @[Bitwise.scala 48:55:@5653.4]
  wire [2:0] _T_7697; // @[Bitwise.scala 48:55:@5653.4]
  wire [1:0] _T_7698; // @[Bitwise.scala 48:55:@5654.4]
  wire [1:0] _T_7699; // @[Bitwise.scala 48:55:@5655.4]
  wire [2:0] _T_7700; // @[Bitwise.scala 48:55:@5656.4]
  wire [3:0] _T_7701; // @[Bitwise.scala 48:55:@5657.4]
  wire [4:0] _T_7702; // @[Bitwise.scala 48:55:@5658.4]
  wire [5:0] _T_7703; // @[Bitwise.scala 48:55:@5659.4]
  wire [6:0] _T_7704; // @[Bitwise.scala 48:55:@5660.4]
  wire [49:0] _T_7768; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5725.4]
  wire  _T_7769; // @[Bitwise.scala 50:65:@5726.4]
  wire  _T_7770; // @[Bitwise.scala 50:65:@5727.4]
  wire  _T_7771; // @[Bitwise.scala 50:65:@5728.4]
  wire  _T_7772; // @[Bitwise.scala 50:65:@5729.4]
  wire  _T_7773; // @[Bitwise.scala 50:65:@5730.4]
  wire  _T_7774; // @[Bitwise.scala 50:65:@5731.4]
  wire  _T_7775; // @[Bitwise.scala 50:65:@5732.4]
  wire  _T_7776; // @[Bitwise.scala 50:65:@5733.4]
  wire  _T_7777; // @[Bitwise.scala 50:65:@5734.4]
  wire  _T_7778; // @[Bitwise.scala 50:65:@5735.4]
  wire  _T_7779; // @[Bitwise.scala 50:65:@5736.4]
  wire  _T_7780; // @[Bitwise.scala 50:65:@5737.4]
  wire  _T_7781; // @[Bitwise.scala 50:65:@5738.4]
  wire  _T_7782; // @[Bitwise.scala 50:65:@5739.4]
  wire  _T_7783; // @[Bitwise.scala 50:65:@5740.4]
  wire  _T_7784; // @[Bitwise.scala 50:65:@5741.4]
  wire  _T_7785; // @[Bitwise.scala 50:65:@5742.4]
  wire  _T_7786; // @[Bitwise.scala 50:65:@5743.4]
  wire  _T_7787; // @[Bitwise.scala 50:65:@5744.4]
  wire  _T_7788; // @[Bitwise.scala 50:65:@5745.4]
  wire  _T_7789; // @[Bitwise.scala 50:65:@5746.4]
  wire  _T_7790; // @[Bitwise.scala 50:65:@5747.4]
  wire  _T_7791; // @[Bitwise.scala 50:65:@5748.4]
  wire  _T_7792; // @[Bitwise.scala 50:65:@5749.4]
  wire  _T_7793; // @[Bitwise.scala 50:65:@5750.4]
  wire  _T_7794; // @[Bitwise.scala 50:65:@5751.4]
  wire  _T_7795; // @[Bitwise.scala 50:65:@5752.4]
  wire  _T_7796; // @[Bitwise.scala 50:65:@5753.4]
  wire  _T_7797; // @[Bitwise.scala 50:65:@5754.4]
  wire  _T_7798; // @[Bitwise.scala 50:65:@5755.4]
  wire  _T_7799; // @[Bitwise.scala 50:65:@5756.4]
  wire  _T_7800; // @[Bitwise.scala 50:65:@5757.4]
  wire  _T_7801; // @[Bitwise.scala 50:65:@5758.4]
  wire  _T_7802; // @[Bitwise.scala 50:65:@5759.4]
  wire  _T_7803; // @[Bitwise.scala 50:65:@5760.4]
  wire  _T_7804; // @[Bitwise.scala 50:65:@5761.4]
  wire  _T_7805; // @[Bitwise.scala 50:65:@5762.4]
  wire  _T_7806; // @[Bitwise.scala 50:65:@5763.4]
  wire  _T_7807; // @[Bitwise.scala 50:65:@5764.4]
  wire  _T_7808; // @[Bitwise.scala 50:65:@5765.4]
  wire  _T_7809; // @[Bitwise.scala 50:65:@5766.4]
  wire  _T_7810; // @[Bitwise.scala 50:65:@5767.4]
  wire  _T_7811; // @[Bitwise.scala 50:65:@5768.4]
  wire  _T_7812; // @[Bitwise.scala 50:65:@5769.4]
  wire  _T_7813; // @[Bitwise.scala 50:65:@5770.4]
  wire  _T_7814; // @[Bitwise.scala 50:65:@5771.4]
  wire  _T_7815; // @[Bitwise.scala 50:65:@5772.4]
  wire  _T_7816; // @[Bitwise.scala 50:65:@5773.4]
  wire  _T_7817; // @[Bitwise.scala 50:65:@5774.4]
  wire  _T_7818; // @[Bitwise.scala 50:65:@5775.4]
  wire [1:0] _T_7819; // @[Bitwise.scala 48:55:@5776.4]
  wire [1:0] _GEN_892; // @[Bitwise.scala 48:55:@5777.4]
  wire [2:0] _T_7820; // @[Bitwise.scala 48:55:@5777.4]
  wire [1:0] _T_7821; // @[Bitwise.scala 48:55:@5778.4]
  wire [1:0] _GEN_893; // @[Bitwise.scala 48:55:@5779.4]
  wire [2:0] _T_7822; // @[Bitwise.scala 48:55:@5779.4]
  wire [3:0] _T_7823; // @[Bitwise.scala 48:55:@5780.4]
  wire [1:0] _T_7824; // @[Bitwise.scala 48:55:@5781.4]
  wire [1:0] _GEN_894; // @[Bitwise.scala 48:55:@5782.4]
  wire [2:0] _T_7825; // @[Bitwise.scala 48:55:@5782.4]
  wire [1:0] _T_7826; // @[Bitwise.scala 48:55:@5783.4]
  wire [1:0] _GEN_895; // @[Bitwise.scala 48:55:@5784.4]
  wire [2:0] _T_7827; // @[Bitwise.scala 48:55:@5784.4]
  wire [3:0] _T_7828; // @[Bitwise.scala 48:55:@5785.4]
  wire [4:0] _T_7829; // @[Bitwise.scala 48:55:@5786.4]
  wire [1:0] _T_7830; // @[Bitwise.scala 48:55:@5787.4]
  wire [1:0] _GEN_896; // @[Bitwise.scala 48:55:@5788.4]
  wire [2:0] _T_7831; // @[Bitwise.scala 48:55:@5788.4]
  wire [1:0] _T_7832; // @[Bitwise.scala 48:55:@5789.4]
  wire [1:0] _GEN_897; // @[Bitwise.scala 48:55:@5790.4]
  wire [2:0] _T_7833; // @[Bitwise.scala 48:55:@5790.4]
  wire [3:0] _T_7834; // @[Bitwise.scala 48:55:@5791.4]
  wire [1:0] _T_7835; // @[Bitwise.scala 48:55:@5792.4]
  wire [1:0] _GEN_898; // @[Bitwise.scala 48:55:@5793.4]
  wire [2:0] _T_7836; // @[Bitwise.scala 48:55:@5793.4]
  wire [1:0] _T_7837; // @[Bitwise.scala 48:55:@5794.4]
  wire [1:0] _T_7838; // @[Bitwise.scala 48:55:@5795.4]
  wire [2:0] _T_7839; // @[Bitwise.scala 48:55:@5796.4]
  wire [3:0] _T_7840; // @[Bitwise.scala 48:55:@5797.4]
  wire [4:0] _T_7841; // @[Bitwise.scala 48:55:@5798.4]
  wire [5:0] _T_7842; // @[Bitwise.scala 48:55:@5799.4]
  wire [1:0] _T_7843; // @[Bitwise.scala 48:55:@5800.4]
  wire [1:0] _GEN_899; // @[Bitwise.scala 48:55:@5801.4]
  wire [2:0] _T_7844; // @[Bitwise.scala 48:55:@5801.4]
  wire [1:0] _T_7845; // @[Bitwise.scala 48:55:@5802.4]
  wire [1:0] _GEN_900; // @[Bitwise.scala 48:55:@5803.4]
  wire [2:0] _T_7846; // @[Bitwise.scala 48:55:@5803.4]
  wire [3:0] _T_7847; // @[Bitwise.scala 48:55:@5804.4]
  wire [1:0] _T_7848; // @[Bitwise.scala 48:55:@5805.4]
  wire [1:0] _GEN_901; // @[Bitwise.scala 48:55:@5806.4]
  wire [2:0] _T_7849; // @[Bitwise.scala 48:55:@5806.4]
  wire [1:0] _T_7850; // @[Bitwise.scala 48:55:@5807.4]
  wire [1:0] _GEN_902; // @[Bitwise.scala 48:55:@5808.4]
  wire [2:0] _T_7851; // @[Bitwise.scala 48:55:@5808.4]
  wire [3:0] _T_7852; // @[Bitwise.scala 48:55:@5809.4]
  wire [4:0] _T_7853; // @[Bitwise.scala 48:55:@5810.4]
  wire [1:0] _T_7854; // @[Bitwise.scala 48:55:@5811.4]
  wire [1:0] _GEN_903; // @[Bitwise.scala 48:55:@5812.4]
  wire [2:0] _T_7855; // @[Bitwise.scala 48:55:@5812.4]
  wire [1:0] _T_7856; // @[Bitwise.scala 48:55:@5813.4]
  wire [1:0] _GEN_904; // @[Bitwise.scala 48:55:@5814.4]
  wire [2:0] _T_7857; // @[Bitwise.scala 48:55:@5814.4]
  wire [3:0] _T_7858; // @[Bitwise.scala 48:55:@5815.4]
  wire [1:0] _T_7859; // @[Bitwise.scala 48:55:@5816.4]
  wire [1:0] _GEN_905; // @[Bitwise.scala 48:55:@5817.4]
  wire [2:0] _T_7860; // @[Bitwise.scala 48:55:@5817.4]
  wire [1:0] _T_7861; // @[Bitwise.scala 48:55:@5818.4]
  wire [1:0] _T_7862; // @[Bitwise.scala 48:55:@5819.4]
  wire [2:0] _T_7863; // @[Bitwise.scala 48:55:@5820.4]
  wire [3:0] _T_7864; // @[Bitwise.scala 48:55:@5821.4]
  wire [4:0] _T_7865; // @[Bitwise.scala 48:55:@5822.4]
  wire [5:0] _T_7866; // @[Bitwise.scala 48:55:@5823.4]
  wire [6:0] _T_7867; // @[Bitwise.scala 48:55:@5824.4]
  wire [50:0] _T_7931; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5889.4]
  wire  _T_7932; // @[Bitwise.scala 50:65:@5890.4]
  wire  _T_7933; // @[Bitwise.scala 50:65:@5891.4]
  wire  _T_7934; // @[Bitwise.scala 50:65:@5892.4]
  wire  _T_7935; // @[Bitwise.scala 50:65:@5893.4]
  wire  _T_7936; // @[Bitwise.scala 50:65:@5894.4]
  wire  _T_7937; // @[Bitwise.scala 50:65:@5895.4]
  wire  _T_7938; // @[Bitwise.scala 50:65:@5896.4]
  wire  _T_7939; // @[Bitwise.scala 50:65:@5897.4]
  wire  _T_7940; // @[Bitwise.scala 50:65:@5898.4]
  wire  _T_7941; // @[Bitwise.scala 50:65:@5899.4]
  wire  _T_7942; // @[Bitwise.scala 50:65:@5900.4]
  wire  _T_7943; // @[Bitwise.scala 50:65:@5901.4]
  wire  _T_7944; // @[Bitwise.scala 50:65:@5902.4]
  wire  _T_7945; // @[Bitwise.scala 50:65:@5903.4]
  wire  _T_7946; // @[Bitwise.scala 50:65:@5904.4]
  wire  _T_7947; // @[Bitwise.scala 50:65:@5905.4]
  wire  _T_7948; // @[Bitwise.scala 50:65:@5906.4]
  wire  _T_7949; // @[Bitwise.scala 50:65:@5907.4]
  wire  _T_7950; // @[Bitwise.scala 50:65:@5908.4]
  wire  _T_7951; // @[Bitwise.scala 50:65:@5909.4]
  wire  _T_7952; // @[Bitwise.scala 50:65:@5910.4]
  wire  _T_7953; // @[Bitwise.scala 50:65:@5911.4]
  wire  _T_7954; // @[Bitwise.scala 50:65:@5912.4]
  wire  _T_7955; // @[Bitwise.scala 50:65:@5913.4]
  wire  _T_7956; // @[Bitwise.scala 50:65:@5914.4]
  wire  _T_7957; // @[Bitwise.scala 50:65:@5915.4]
  wire  _T_7958; // @[Bitwise.scala 50:65:@5916.4]
  wire  _T_7959; // @[Bitwise.scala 50:65:@5917.4]
  wire  _T_7960; // @[Bitwise.scala 50:65:@5918.4]
  wire  _T_7961; // @[Bitwise.scala 50:65:@5919.4]
  wire  _T_7962; // @[Bitwise.scala 50:65:@5920.4]
  wire  _T_7963; // @[Bitwise.scala 50:65:@5921.4]
  wire  _T_7964; // @[Bitwise.scala 50:65:@5922.4]
  wire  _T_7965; // @[Bitwise.scala 50:65:@5923.4]
  wire  _T_7966; // @[Bitwise.scala 50:65:@5924.4]
  wire  _T_7967; // @[Bitwise.scala 50:65:@5925.4]
  wire  _T_7968; // @[Bitwise.scala 50:65:@5926.4]
  wire  _T_7969; // @[Bitwise.scala 50:65:@5927.4]
  wire  _T_7970; // @[Bitwise.scala 50:65:@5928.4]
  wire  _T_7971; // @[Bitwise.scala 50:65:@5929.4]
  wire  _T_7972; // @[Bitwise.scala 50:65:@5930.4]
  wire  _T_7973; // @[Bitwise.scala 50:65:@5931.4]
  wire  _T_7974; // @[Bitwise.scala 50:65:@5932.4]
  wire  _T_7975; // @[Bitwise.scala 50:65:@5933.4]
  wire  _T_7976; // @[Bitwise.scala 50:65:@5934.4]
  wire  _T_7977; // @[Bitwise.scala 50:65:@5935.4]
  wire  _T_7978; // @[Bitwise.scala 50:65:@5936.4]
  wire  _T_7979; // @[Bitwise.scala 50:65:@5937.4]
  wire  _T_7980; // @[Bitwise.scala 50:65:@5938.4]
  wire  _T_7981; // @[Bitwise.scala 50:65:@5939.4]
  wire  _T_7982; // @[Bitwise.scala 50:65:@5940.4]
  wire [1:0] _T_7983; // @[Bitwise.scala 48:55:@5941.4]
  wire [1:0] _GEN_906; // @[Bitwise.scala 48:55:@5942.4]
  wire [2:0] _T_7984; // @[Bitwise.scala 48:55:@5942.4]
  wire [1:0] _T_7985; // @[Bitwise.scala 48:55:@5943.4]
  wire [1:0] _GEN_907; // @[Bitwise.scala 48:55:@5944.4]
  wire [2:0] _T_7986; // @[Bitwise.scala 48:55:@5944.4]
  wire [3:0] _T_7987; // @[Bitwise.scala 48:55:@5945.4]
  wire [1:0] _T_7988; // @[Bitwise.scala 48:55:@5946.4]
  wire [1:0] _GEN_908; // @[Bitwise.scala 48:55:@5947.4]
  wire [2:0] _T_7989; // @[Bitwise.scala 48:55:@5947.4]
  wire [1:0] _T_7990; // @[Bitwise.scala 48:55:@5948.4]
  wire [1:0] _GEN_909; // @[Bitwise.scala 48:55:@5949.4]
  wire [2:0] _T_7991; // @[Bitwise.scala 48:55:@5949.4]
  wire [3:0] _T_7992; // @[Bitwise.scala 48:55:@5950.4]
  wire [4:0] _T_7993; // @[Bitwise.scala 48:55:@5951.4]
  wire [1:0] _T_7994; // @[Bitwise.scala 48:55:@5952.4]
  wire [1:0] _GEN_910; // @[Bitwise.scala 48:55:@5953.4]
  wire [2:0] _T_7995; // @[Bitwise.scala 48:55:@5953.4]
  wire [1:0] _T_7996; // @[Bitwise.scala 48:55:@5954.4]
  wire [1:0] _GEN_911; // @[Bitwise.scala 48:55:@5955.4]
  wire [2:0] _T_7997; // @[Bitwise.scala 48:55:@5955.4]
  wire [3:0] _T_7998; // @[Bitwise.scala 48:55:@5956.4]
  wire [1:0] _T_7999; // @[Bitwise.scala 48:55:@5957.4]
  wire [1:0] _GEN_912; // @[Bitwise.scala 48:55:@5958.4]
  wire [2:0] _T_8000; // @[Bitwise.scala 48:55:@5958.4]
  wire [1:0] _T_8001; // @[Bitwise.scala 48:55:@5959.4]
  wire [1:0] _T_8002; // @[Bitwise.scala 48:55:@5960.4]
  wire [2:0] _T_8003; // @[Bitwise.scala 48:55:@5961.4]
  wire [3:0] _T_8004; // @[Bitwise.scala 48:55:@5962.4]
  wire [4:0] _T_8005; // @[Bitwise.scala 48:55:@5963.4]
  wire [5:0] _T_8006; // @[Bitwise.scala 48:55:@5964.4]
  wire [1:0] _T_8007; // @[Bitwise.scala 48:55:@5965.4]
  wire [1:0] _GEN_913; // @[Bitwise.scala 48:55:@5966.4]
  wire [2:0] _T_8008; // @[Bitwise.scala 48:55:@5966.4]
  wire [1:0] _T_8009; // @[Bitwise.scala 48:55:@5967.4]
  wire [1:0] _GEN_914; // @[Bitwise.scala 48:55:@5968.4]
  wire [2:0] _T_8010; // @[Bitwise.scala 48:55:@5968.4]
  wire [3:0] _T_8011; // @[Bitwise.scala 48:55:@5969.4]
  wire [1:0] _T_8012; // @[Bitwise.scala 48:55:@5970.4]
  wire [1:0] _GEN_915; // @[Bitwise.scala 48:55:@5971.4]
  wire [2:0] _T_8013; // @[Bitwise.scala 48:55:@5971.4]
  wire [1:0] _T_8014; // @[Bitwise.scala 48:55:@5972.4]
  wire [1:0] _T_8015; // @[Bitwise.scala 48:55:@5973.4]
  wire [2:0] _T_8016; // @[Bitwise.scala 48:55:@5974.4]
  wire [3:0] _T_8017; // @[Bitwise.scala 48:55:@5975.4]
  wire [4:0] _T_8018; // @[Bitwise.scala 48:55:@5976.4]
  wire [1:0] _T_8019; // @[Bitwise.scala 48:55:@5977.4]
  wire [1:0] _GEN_916; // @[Bitwise.scala 48:55:@5978.4]
  wire [2:0] _T_8020; // @[Bitwise.scala 48:55:@5978.4]
  wire [1:0] _T_8021; // @[Bitwise.scala 48:55:@5979.4]
  wire [1:0] _GEN_917; // @[Bitwise.scala 48:55:@5980.4]
  wire [2:0] _T_8022; // @[Bitwise.scala 48:55:@5980.4]
  wire [3:0] _T_8023; // @[Bitwise.scala 48:55:@5981.4]
  wire [1:0] _T_8024; // @[Bitwise.scala 48:55:@5982.4]
  wire [1:0] _GEN_918; // @[Bitwise.scala 48:55:@5983.4]
  wire [2:0] _T_8025; // @[Bitwise.scala 48:55:@5983.4]
  wire [1:0] _T_8026; // @[Bitwise.scala 48:55:@5984.4]
  wire [1:0] _T_8027; // @[Bitwise.scala 48:55:@5985.4]
  wire [2:0] _T_8028; // @[Bitwise.scala 48:55:@5986.4]
  wire [3:0] _T_8029; // @[Bitwise.scala 48:55:@5987.4]
  wire [4:0] _T_8030; // @[Bitwise.scala 48:55:@5988.4]
  wire [5:0] _T_8031; // @[Bitwise.scala 48:55:@5989.4]
  wire [6:0] _T_8032; // @[Bitwise.scala 48:55:@5990.4]
  wire [51:0] _T_8096; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6055.4]
  wire  _T_8097; // @[Bitwise.scala 50:65:@6056.4]
  wire  _T_8098; // @[Bitwise.scala 50:65:@6057.4]
  wire  _T_8099; // @[Bitwise.scala 50:65:@6058.4]
  wire  _T_8100; // @[Bitwise.scala 50:65:@6059.4]
  wire  _T_8101; // @[Bitwise.scala 50:65:@6060.4]
  wire  _T_8102; // @[Bitwise.scala 50:65:@6061.4]
  wire  _T_8103; // @[Bitwise.scala 50:65:@6062.4]
  wire  _T_8104; // @[Bitwise.scala 50:65:@6063.4]
  wire  _T_8105; // @[Bitwise.scala 50:65:@6064.4]
  wire  _T_8106; // @[Bitwise.scala 50:65:@6065.4]
  wire  _T_8107; // @[Bitwise.scala 50:65:@6066.4]
  wire  _T_8108; // @[Bitwise.scala 50:65:@6067.4]
  wire  _T_8109; // @[Bitwise.scala 50:65:@6068.4]
  wire  _T_8110; // @[Bitwise.scala 50:65:@6069.4]
  wire  _T_8111; // @[Bitwise.scala 50:65:@6070.4]
  wire  _T_8112; // @[Bitwise.scala 50:65:@6071.4]
  wire  _T_8113; // @[Bitwise.scala 50:65:@6072.4]
  wire  _T_8114; // @[Bitwise.scala 50:65:@6073.4]
  wire  _T_8115; // @[Bitwise.scala 50:65:@6074.4]
  wire  _T_8116; // @[Bitwise.scala 50:65:@6075.4]
  wire  _T_8117; // @[Bitwise.scala 50:65:@6076.4]
  wire  _T_8118; // @[Bitwise.scala 50:65:@6077.4]
  wire  _T_8119; // @[Bitwise.scala 50:65:@6078.4]
  wire  _T_8120; // @[Bitwise.scala 50:65:@6079.4]
  wire  _T_8121; // @[Bitwise.scala 50:65:@6080.4]
  wire  _T_8122; // @[Bitwise.scala 50:65:@6081.4]
  wire  _T_8123; // @[Bitwise.scala 50:65:@6082.4]
  wire  _T_8124; // @[Bitwise.scala 50:65:@6083.4]
  wire  _T_8125; // @[Bitwise.scala 50:65:@6084.4]
  wire  _T_8126; // @[Bitwise.scala 50:65:@6085.4]
  wire  _T_8127; // @[Bitwise.scala 50:65:@6086.4]
  wire  _T_8128; // @[Bitwise.scala 50:65:@6087.4]
  wire  _T_8129; // @[Bitwise.scala 50:65:@6088.4]
  wire  _T_8130; // @[Bitwise.scala 50:65:@6089.4]
  wire  _T_8131; // @[Bitwise.scala 50:65:@6090.4]
  wire  _T_8132; // @[Bitwise.scala 50:65:@6091.4]
  wire  _T_8133; // @[Bitwise.scala 50:65:@6092.4]
  wire  _T_8134; // @[Bitwise.scala 50:65:@6093.4]
  wire  _T_8135; // @[Bitwise.scala 50:65:@6094.4]
  wire  _T_8136; // @[Bitwise.scala 50:65:@6095.4]
  wire  _T_8137; // @[Bitwise.scala 50:65:@6096.4]
  wire  _T_8138; // @[Bitwise.scala 50:65:@6097.4]
  wire  _T_8139; // @[Bitwise.scala 50:65:@6098.4]
  wire  _T_8140; // @[Bitwise.scala 50:65:@6099.4]
  wire  _T_8141; // @[Bitwise.scala 50:65:@6100.4]
  wire  _T_8142; // @[Bitwise.scala 50:65:@6101.4]
  wire  _T_8143; // @[Bitwise.scala 50:65:@6102.4]
  wire  _T_8144; // @[Bitwise.scala 50:65:@6103.4]
  wire  _T_8145; // @[Bitwise.scala 50:65:@6104.4]
  wire  _T_8146; // @[Bitwise.scala 50:65:@6105.4]
  wire  _T_8147; // @[Bitwise.scala 50:65:@6106.4]
  wire  _T_8148; // @[Bitwise.scala 50:65:@6107.4]
  wire [1:0] _T_8149; // @[Bitwise.scala 48:55:@6108.4]
  wire [1:0] _GEN_919; // @[Bitwise.scala 48:55:@6109.4]
  wire [2:0] _T_8150; // @[Bitwise.scala 48:55:@6109.4]
  wire [1:0] _T_8151; // @[Bitwise.scala 48:55:@6110.4]
  wire [1:0] _GEN_920; // @[Bitwise.scala 48:55:@6111.4]
  wire [2:0] _T_8152; // @[Bitwise.scala 48:55:@6111.4]
  wire [3:0] _T_8153; // @[Bitwise.scala 48:55:@6112.4]
  wire [1:0] _T_8154; // @[Bitwise.scala 48:55:@6113.4]
  wire [1:0] _GEN_921; // @[Bitwise.scala 48:55:@6114.4]
  wire [2:0] _T_8155; // @[Bitwise.scala 48:55:@6114.4]
  wire [1:0] _T_8156; // @[Bitwise.scala 48:55:@6115.4]
  wire [1:0] _T_8157; // @[Bitwise.scala 48:55:@6116.4]
  wire [2:0] _T_8158; // @[Bitwise.scala 48:55:@6117.4]
  wire [3:0] _T_8159; // @[Bitwise.scala 48:55:@6118.4]
  wire [4:0] _T_8160; // @[Bitwise.scala 48:55:@6119.4]
  wire [1:0] _T_8161; // @[Bitwise.scala 48:55:@6120.4]
  wire [1:0] _GEN_922; // @[Bitwise.scala 48:55:@6121.4]
  wire [2:0] _T_8162; // @[Bitwise.scala 48:55:@6121.4]
  wire [1:0] _T_8163; // @[Bitwise.scala 48:55:@6122.4]
  wire [1:0] _GEN_923; // @[Bitwise.scala 48:55:@6123.4]
  wire [2:0] _T_8164; // @[Bitwise.scala 48:55:@6123.4]
  wire [3:0] _T_8165; // @[Bitwise.scala 48:55:@6124.4]
  wire [1:0] _T_8166; // @[Bitwise.scala 48:55:@6125.4]
  wire [1:0] _GEN_924; // @[Bitwise.scala 48:55:@6126.4]
  wire [2:0] _T_8167; // @[Bitwise.scala 48:55:@6126.4]
  wire [1:0] _T_8168; // @[Bitwise.scala 48:55:@6127.4]
  wire [1:0] _T_8169; // @[Bitwise.scala 48:55:@6128.4]
  wire [2:0] _T_8170; // @[Bitwise.scala 48:55:@6129.4]
  wire [3:0] _T_8171; // @[Bitwise.scala 48:55:@6130.4]
  wire [4:0] _T_8172; // @[Bitwise.scala 48:55:@6131.4]
  wire [5:0] _T_8173; // @[Bitwise.scala 48:55:@6132.4]
  wire [1:0] _T_8174; // @[Bitwise.scala 48:55:@6133.4]
  wire [1:0] _GEN_925; // @[Bitwise.scala 48:55:@6134.4]
  wire [2:0] _T_8175; // @[Bitwise.scala 48:55:@6134.4]
  wire [1:0] _T_8176; // @[Bitwise.scala 48:55:@6135.4]
  wire [1:0] _GEN_926; // @[Bitwise.scala 48:55:@6136.4]
  wire [2:0] _T_8177; // @[Bitwise.scala 48:55:@6136.4]
  wire [3:0] _T_8178; // @[Bitwise.scala 48:55:@6137.4]
  wire [1:0] _T_8179; // @[Bitwise.scala 48:55:@6138.4]
  wire [1:0] _GEN_927; // @[Bitwise.scala 48:55:@6139.4]
  wire [2:0] _T_8180; // @[Bitwise.scala 48:55:@6139.4]
  wire [1:0] _T_8181; // @[Bitwise.scala 48:55:@6140.4]
  wire [1:0] _T_8182; // @[Bitwise.scala 48:55:@6141.4]
  wire [2:0] _T_8183; // @[Bitwise.scala 48:55:@6142.4]
  wire [3:0] _T_8184; // @[Bitwise.scala 48:55:@6143.4]
  wire [4:0] _T_8185; // @[Bitwise.scala 48:55:@6144.4]
  wire [1:0] _T_8186; // @[Bitwise.scala 48:55:@6145.4]
  wire [1:0] _GEN_928; // @[Bitwise.scala 48:55:@6146.4]
  wire [2:0] _T_8187; // @[Bitwise.scala 48:55:@6146.4]
  wire [1:0] _T_8188; // @[Bitwise.scala 48:55:@6147.4]
  wire [1:0] _GEN_929; // @[Bitwise.scala 48:55:@6148.4]
  wire [2:0] _T_8189; // @[Bitwise.scala 48:55:@6148.4]
  wire [3:0] _T_8190; // @[Bitwise.scala 48:55:@6149.4]
  wire [1:0] _T_8191; // @[Bitwise.scala 48:55:@6150.4]
  wire [1:0] _GEN_930; // @[Bitwise.scala 48:55:@6151.4]
  wire [2:0] _T_8192; // @[Bitwise.scala 48:55:@6151.4]
  wire [1:0] _T_8193; // @[Bitwise.scala 48:55:@6152.4]
  wire [1:0] _T_8194; // @[Bitwise.scala 48:55:@6153.4]
  wire [2:0] _T_8195; // @[Bitwise.scala 48:55:@6154.4]
  wire [3:0] _T_8196; // @[Bitwise.scala 48:55:@6155.4]
  wire [4:0] _T_8197; // @[Bitwise.scala 48:55:@6156.4]
  wire [5:0] _T_8198; // @[Bitwise.scala 48:55:@6157.4]
  wire [6:0] _T_8199; // @[Bitwise.scala 48:55:@6158.4]
  wire [52:0] _T_8263; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6223.4]
  wire  _T_8264; // @[Bitwise.scala 50:65:@6224.4]
  wire  _T_8265; // @[Bitwise.scala 50:65:@6225.4]
  wire  _T_8266; // @[Bitwise.scala 50:65:@6226.4]
  wire  _T_8267; // @[Bitwise.scala 50:65:@6227.4]
  wire  _T_8268; // @[Bitwise.scala 50:65:@6228.4]
  wire  _T_8269; // @[Bitwise.scala 50:65:@6229.4]
  wire  _T_8270; // @[Bitwise.scala 50:65:@6230.4]
  wire  _T_8271; // @[Bitwise.scala 50:65:@6231.4]
  wire  _T_8272; // @[Bitwise.scala 50:65:@6232.4]
  wire  _T_8273; // @[Bitwise.scala 50:65:@6233.4]
  wire  _T_8274; // @[Bitwise.scala 50:65:@6234.4]
  wire  _T_8275; // @[Bitwise.scala 50:65:@6235.4]
  wire  _T_8276; // @[Bitwise.scala 50:65:@6236.4]
  wire  _T_8277; // @[Bitwise.scala 50:65:@6237.4]
  wire  _T_8278; // @[Bitwise.scala 50:65:@6238.4]
  wire  _T_8279; // @[Bitwise.scala 50:65:@6239.4]
  wire  _T_8280; // @[Bitwise.scala 50:65:@6240.4]
  wire  _T_8281; // @[Bitwise.scala 50:65:@6241.4]
  wire  _T_8282; // @[Bitwise.scala 50:65:@6242.4]
  wire  _T_8283; // @[Bitwise.scala 50:65:@6243.4]
  wire  _T_8284; // @[Bitwise.scala 50:65:@6244.4]
  wire  _T_8285; // @[Bitwise.scala 50:65:@6245.4]
  wire  _T_8286; // @[Bitwise.scala 50:65:@6246.4]
  wire  _T_8287; // @[Bitwise.scala 50:65:@6247.4]
  wire  _T_8288; // @[Bitwise.scala 50:65:@6248.4]
  wire  _T_8289; // @[Bitwise.scala 50:65:@6249.4]
  wire  _T_8290; // @[Bitwise.scala 50:65:@6250.4]
  wire  _T_8291; // @[Bitwise.scala 50:65:@6251.4]
  wire  _T_8292; // @[Bitwise.scala 50:65:@6252.4]
  wire  _T_8293; // @[Bitwise.scala 50:65:@6253.4]
  wire  _T_8294; // @[Bitwise.scala 50:65:@6254.4]
  wire  _T_8295; // @[Bitwise.scala 50:65:@6255.4]
  wire  _T_8296; // @[Bitwise.scala 50:65:@6256.4]
  wire  _T_8297; // @[Bitwise.scala 50:65:@6257.4]
  wire  _T_8298; // @[Bitwise.scala 50:65:@6258.4]
  wire  _T_8299; // @[Bitwise.scala 50:65:@6259.4]
  wire  _T_8300; // @[Bitwise.scala 50:65:@6260.4]
  wire  _T_8301; // @[Bitwise.scala 50:65:@6261.4]
  wire  _T_8302; // @[Bitwise.scala 50:65:@6262.4]
  wire  _T_8303; // @[Bitwise.scala 50:65:@6263.4]
  wire  _T_8304; // @[Bitwise.scala 50:65:@6264.4]
  wire  _T_8305; // @[Bitwise.scala 50:65:@6265.4]
  wire  _T_8306; // @[Bitwise.scala 50:65:@6266.4]
  wire  _T_8307; // @[Bitwise.scala 50:65:@6267.4]
  wire  _T_8308; // @[Bitwise.scala 50:65:@6268.4]
  wire  _T_8309; // @[Bitwise.scala 50:65:@6269.4]
  wire  _T_8310; // @[Bitwise.scala 50:65:@6270.4]
  wire  _T_8311; // @[Bitwise.scala 50:65:@6271.4]
  wire  _T_8312; // @[Bitwise.scala 50:65:@6272.4]
  wire  _T_8313; // @[Bitwise.scala 50:65:@6273.4]
  wire  _T_8314; // @[Bitwise.scala 50:65:@6274.4]
  wire  _T_8315; // @[Bitwise.scala 50:65:@6275.4]
  wire  _T_8316; // @[Bitwise.scala 50:65:@6276.4]
  wire [1:0] _T_8317; // @[Bitwise.scala 48:55:@6277.4]
  wire [1:0] _GEN_931; // @[Bitwise.scala 48:55:@6278.4]
  wire [2:0] _T_8318; // @[Bitwise.scala 48:55:@6278.4]
  wire [1:0] _T_8319; // @[Bitwise.scala 48:55:@6279.4]
  wire [1:0] _GEN_932; // @[Bitwise.scala 48:55:@6280.4]
  wire [2:0] _T_8320; // @[Bitwise.scala 48:55:@6280.4]
  wire [3:0] _T_8321; // @[Bitwise.scala 48:55:@6281.4]
  wire [1:0] _T_8322; // @[Bitwise.scala 48:55:@6282.4]
  wire [1:0] _GEN_933; // @[Bitwise.scala 48:55:@6283.4]
  wire [2:0] _T_8323; // @[Bitwise.scala 48:55:@6283.4]
  wire [1:0] _T_8324; // @[Bitwise.scala 48:55:@6284.4]
  wire [1:0] _T_8325; // @[Bitwise.scala 48:55:@6285.4]
  wire [2:0] _T_8326; // @[Bitwise.scala 48:55:@6286.4]
  wire [3:0] _T_8327; // @[Bitwise.scala 48:55:@6287.4]
  wire [4:0] _T_8328; // @[Bitwise.scala 48:55:@6288.4]
  wire [1:0] _T_8329; // @[Bitwise.scala 48:55:@6289.4]
  wire [1:0] _GEN_934; // @[Bitwise.scala 48:55:@6290.4]
  wire [2:0] _T_8330; // @[Bitwise.scala 48:55:@6290.4]
  wire [1:0] _T_8331; // @[Bitwise.scala 48:55:@6291.4]
  wire [1:0] _GEN_935; // @[Bitwise.scala 48:55:@6292.4]
  wire [2:0] _T_8332; // @[Bitwise.scala 48:55:@6292.4]
  wire [3:0] _T_8333; // @[Bitwise.scala 48:55:@6293.4]
  wire [1:0] _T_8334; // @[Bitwise.scala 48:55:@6294.4]
  wire [1:0] _GEN_936; // @[Bitwise.scala 48:55:@6295.4]
  wire [2:0] _T_8335; // @[Bitwise.scala 48:55:@6295.4]
  wire [1:0] _T_8336; // @[Bitwise.scala 48:55:@6296.4]
  wire [1:0] _T_8337; // @[Bitwise.scala 48:55:@6297.4]
  wire [2:0] _T_8338; // @[Bitwise.scala 48:55:@6298.4]
  wire [3:0] _T_8339; // @[Bitwise.scala 48:55:@6299.4]
  wire [4:0] _T_8340; // @[Bitwise.scala 48:55:@6300.4]
  wire [5:0] _T_8341; // @[Bitwise.scala 48:55:@6301.4]
  wire [1:0] _T_8342; // @[Bitwise.scala 48:55:@6302.4]
  wire [1:0] _GEN_937; // @[Bitwise.scala 48:55:@6303.4]
  wire [2:0] _T_8343; // @[Bitwise.scala 48:55:@6303.4]
  wire [1:0] _T_8344; // @[Bitwise.scala 48:55:@6304.4]
  wire [1:0] _GEN_938; // @[Bitwise.scala 48:55:@6305.4]
  wire [2:0] _T_8345; // @[Bitwise.scala 48:55:@6305.4]
  wire [3:0] _T_8346; // @[Bitwise.scala 48:55:@6306.4]
  wire [1:0] _T_8347; // @[Bitwise.scala 48:55:@6307.4]
  wire [1:0] _GEN_939; // @[Bitwise.scala 48:55:@6308.4]
  wire [2:0] _T_8348; // @[Bitwise.scala 48:55:@6308.4]
  wire [1:0] _T_8349; // @[Bitwise.scala 48:55:@6309.4]
  wire [1:0] _T_8350; // @[Bitwise.scala 48:55:@6310.4]
  wire [2:0] _T_8351; // @[Bitwise.scala 48:55:@6311.4]
  wire [3:0] _T_8352; // @[Bitwise.scala 48:55:@6312.4]
  wire [4:0] _T_8353; // @[Bitwise.scala 48:55:@6313.4]
  wire [1:0] _T_8354; // @[Bitwise.scala 48:55:@6314.4]
  wire [1:0] _GEN_940; // @[Bitwise.scala 48:55:@6315.4]
  wire [2:0] _T_8355; // @[Bitwise.scala 48:55:@6315.4]
  wire [1:0] _T_8356; // @[Bitwise.scala 48:55:@6316.4]
  wire [1:0] _T_8357; // @[Bitwise.scala 48:55:@6317.4]
  wire [2:0] _T_8358; // @[Bitwise.scala 48:55:@6318.4]
  wire [3:0] _T_8359; // @[Bitwise.scala 48:55:@6319.4]
  wire [1:0] _T_8360; // @[Bitwise.scala 48:55:@6320.4]
  wire [1:0] _GEN_941; // @[Bitwise.scala 48:55:@6321.4]
  wire [2:0] _T_8361; // @[Bitwise.scala 48:55:@6321.4]
  wire [1:0] _T_8362; // @[Bitwise.scala 48:55:@6322.4]
  wire [1:0] _T_8363; // @[Bitwise.scala 48:55:@6323.4]
  wire [2:0] _T_8364; // @[Bitwise.scala 48:55:@6324.4]
  wire [3:0] _T_8365; // @[Bitwise.scala 48:55:@6325.4]
  wire [4:0] _T_8366; // @[Bitwise.scala 48:55:@6326.4]
  wire [5:0] _T_8367; // @[Bitwise.scala 48:55:@6327.4]
  wire [6:0] _T_8368; // @[Bitwise.scala 48:55:@6328.4]
  wire [53:0] _T_8432; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6393.4]
  wire  _T_8433; // @[Bitwise.scala 50:65:@6394.4]
  wire  _T_8434; // @[Bitwise.scala 50:65:@6395.4]
  wire  _T_8435; // @[Bitwise.scala 50:65:@6396.4]
  wire  _T_8436; // @[Bitwise.scala 50:65:@6397.4]
  wire  _T_8437; // @[Bitwise.scala 50:65:@6398.4]
  wire  _T_8438; // @[Bitwise.scala 50:65:@6399.4]
  wire  _T_8439; // @[Bitwise.scala 50:65:@6400.4]
  wire  _T_8440; // @[Bitwise.scala 50:65:@6401.4]
  wire  _T_8441; // @[Bitwise.scala 50:65:@6402.4]
  wire  _T_8442; // @[Bitwise.scala 50:65:@6403.4]
  wire  _T_8443; // @[Bitwise.scala 50:65:@6404.4]
  wire  _T_8444; // @[Bitwise.scala 50:65:@6405.4]
  wire  _T_8445; // @[Bitwise.scala 50:65:@6406.4]
  wire  _T_8446; // @[Bitwise.scala 50:65:@6407.4]
  wire  _T_8447; // @[Bitwise.scala 50:65:@6408.4]
  wire  _T_8448; // @[Bitwise.scala 50:65:@6409.4]
  wire  _T_8449; // @[Bitwise.scala 50:65:@6410.4]
  wire  _T_8450; // @[Bitwise.scala 50:65:@6411.4]
  wire  _T_8451; // @[Bitwise.scala 50:65:@6412.4]
  wire  _T_8452; // @[Bitwise.scala 50:65:@6413.4]
  wire  _T_8453; // @[Bitwise.scala 50:65:@6414.4]
  wire  _T_8454; // @[Bitwise.scala 50:65:@6415.4]
  wire  _T_8455; // @[Bitwise.scala 50:65:@6416.4]
  wire  _T_8456; // @[Bitwise.scala 50:65:@6417.4]
  wire  _T_8457; // @[Bitwise.scala 50:65:@6418.4]
  wire  _T_8458; // @[Bitwise.scala 50:65:@6419.4]
  wire  _T_8459; // @[Bitwise.scala 50:65:@6420.4]
  wire  _T_8460; // @[Bitwise.scala 50:65:@6421.4]
  wire  _T_8461; // @[Bitwise.scala 50:65:@6422.4]
  wire  _T_8462; // @[Bitwise.scala 50:65:@6423.4]
  wire  _T_8463; // @[Bitwise.scala 50:65:@6424.4]
  wire  _T_8464; // @[Bitwise.scala 50:65:@6425.4]
  wire  _T_8465; // @[Bitwise.scala 50:65:@6426.4]
  wire  _T_8466; // @[Bitwise.scala 50:65:@6427.4]
  wire  _T_8467; // @[Bitwise.scala 50:65:@6428.4]
  wire  _T_8468; // @[Bitwise.scala 50:65:@6429.4]
  wire  _T_8469; // @[Bitwise.scala 50:65:@6430.4]
  wire  _T_8470; // @[Bitwise.scala 50:65:@6431.4]
  wire  _T_8471; // @[Bitwise.scala 50:65:@6432.4]
  wire  _T_8472; // @[Bitwise.scala 50:65:@6433.4]
  wire  _T_8473; // @[Bitwise.scala 50:65:@6434.4]
  wire  _T_8474; // @[Bitwise.scala 50:65:@6435.4]
  wire  _T_8475; // @[Bitwise.scala 50:65:@6436.4]
  wire  _T_8476; // @[Bitwise.scala 50:65:@6437.4]
  wire  _T_8477; // @[Bitwise.scala 50:65:@6438.4]
  wire  _T_8478; // @[Bitwise.scala 50:65:@6439.4]
  wire  _T_8479; // @[Bitwise.scala 50:65:@6440.4]
  wire  _T_8480; // @[Bitwise.scala 50:65:@6441.4]
  wire  _T_8481; // @[Bitwise.scala 50:65:@6442.4]
  wire  _T_8482; // @[Bitwise.scala 50:65:@6443.4]
  wire  _T_8483; // @[Bitwise.scala 50:65:@6444.4]
  wire  _T_8484; // @[Bitwise.scala 50:65:@6445.4]
  wire  _T_8485; // @[Bitwise.scala 50:65:@6446.4]
  wire  _T_8486; // @[Bitwise.scala 50:65:@6447.4]
  wire [1:0] _T_8487; // @[Bitwise.scala 48:55:@6448.4]
  wire [1:0] _GEN_942; // @[Bitwise.scala 48:55:@6449.4]
  wire [2:0] _T_8488; // @[Bitwise.scala 48:55:@6449.4]
  wire [1:0] _T_8489; // @[Bitwise.scala 48:55:@6450.4]
  wire [1:0] _GEN_943; // @[Bitwise.scala 48:55:@6451.4]
  wire [2:0] _T_8490; // @[Bitwise.scala 48:55:@6451.4]
  wire [3:0] _T_8491; // @[Bitwise.scala 48:55:@6452.4]
  wire [1:0] _T_8492; // @[Bitwise.scala 48:55:@6453.4]
  wire [1:0] _GEN_944; // @[Bitwise.scala 48:55:@6454.4]
  wire [2:0] _T_8493; // @[Bitwise.scala 48:55:@6454.4]
  wire [1:0] _T_8494; // @[Bitwise.scala 48:55:@6455.4]
  wire [1:0] _T_8495; // @[Bitwise.scala 48:55:@6456.4]
  wire [2:0] _T_8496; // @[Bitwise.scala 48:55:@6457.4]
  wire [3:0] _T_8497; // @[Bitwise.scala 48:55:@6458.4]
  wire [4:0] _T_8498; // @[Bitwise.scala 48:55:@6459.4]
  wire [1:0] _T_8499; // @[Bitwise.scala 48:55:@6460.4]
  wire [1:0] _GEN_945; // @[Bitwise.scala 48:55:@6461.4]
  wire [2:0] _T_8500; // @[Bitwise.scala 48:55:@6461.4]
  wire [1:0] _T_8501; // @[Bitwise.scala 48:55:@6462.4]
  wire [1:0] _T_8502; // @[Bitwise.scala 48:55:@6463.4]
  wire [2:0] _T_8503; // @[Bitwise.scala 48:55:@6464.4]
  wire [3:0] _T_8504; // @[Bitwise.scala 48:55:@6465.4]
  wire [1:0] _T_8505; // @[Bitwise.scala 48:55:@6466.4]
  wire [1:0] _GEN_946; // @[Bitwise.scala 48:55:@6467.4]
  wire [2:0] _T_8506; // @[Bitwise.scala 48:55:@6467.4]
  wire [1:0] _T_8507; // @[Bitwise.scala 48:55:@6468.4]
  wire [1:0] _T_8508; // @[Bitwise.scala 48:55:@6469.4]
  wire [2:0] _T_8509; // @[Bitwise.scala 48:55:@6470.4]
  wire [3:0] _T_8510; // @[Bitwise.scala 48:55:@6471.4]
  wire [4:0] _T_8511; // @[Bitwise.scala 48:55:@6472.4]
  wire [5:0] _T_8512; // @[Bitwise.scala 48:55:@6473.4]
  wire [1:0] _T_8513; // @[Bitwise.scala 48:55:@6474.4]
  wire [1:0] _GEN_947; // @[Bitwise.scala 48:55:@6475.4]
  wire [2:0] _T_8514; // @[Bitwise.scala 48:55:@6475.4]
  wire [1:0] _T_8515; // @[Bitwise.scala 48:55:@6476.4]
  wire [1:0] _GEN_948; // @[Bitwise.scala 48:55:@6477.4]
  wire [2:0] _T_8516; // @[Bitwise.scala 48:55:@6477.4]
  wire [3:0] _T_8517; // @[Bitwise.scala 48:55:@6478.4]
  wire [1:0] _T_8518; // @[Bitwise.scala 48:55:@6479.4]
  wire [1:0] _GEN_949; // @[Bitwise.scala 48:55:@6480.4]
  wire [2:0] _T_8519; // @[Bitwise.scala 48:55:@6480.4]
  wire [1:0] _T_8520; // @[Bitwise.scala 48:55:@6481.4]
  wire [1:0] _T_8521; // @[Bitwise.scala 48:55:@6482.4]
  wire [2:0] _T_8522; // @[Bitwise.scala 48:55:@6483.4]
  wire [3:0] _T_8523; // @[Bitwise.scala 48:55:@6484.4]
  wire [4:0] _T_8524; // @[Bitwise.scala 48:55:@6485.4]
  wire [1:0] _T_8525; // @[Bitwise.scala 48:55:@6486.4]
  wire [1:0] _GEN_950; // @[Bitwise.scala 48:55:@6487.4]
  wire [2:0] _T_8526; // @[Bitwise.scala 48:55:@6487.4]
  wire [1:0] _T_8527; // @[Bitwise.scala 48:55:@6488.4]
  wire [1:0] _T_8528; // @[Bitwise.scala 48:55:@6489.4]
  wire [2:0] _T_8529; // @[Bitwise.scala 48:55:@6490.4]
  wire [3:0] _T_8530; // @[Bitwise.scala 48:55:@6491.4]
  wire [1:0] _T_8531; // @[Bitwise.scala 48:55:@6492.4]
  wire [1:0] _GEN_951; // @[Bitwise.scala 48:55:@6493.4]
  wire [2:0] _T_8532; // @[Bitwise.scala 48:55:@6493.4]
  wire [1:0] _T_8533; // @[Bitwise.scala 48:55:@6494.4]
  wire [1:0] _T_8534; // @[Bitwise.scala 48:55:@6495.4]
  wire [2:0] _T_8535; // @[Bitwise.scala 48:55:@6496.4]
  wire [3:0] _T_8536; // @[Bitwise.scala 48:55:@6497.4]
  wire [4:0] _T_8537; // @[Bitwise.scala 48:55:@6498.4]
  wire [5:0] _T_8538; // @[Bitwise.scala 48:55:@6499.4]
  wire [6:0] _T_8539; // @[Bitwise.scala 48:55:@6500.4]
  wire [54:0] _T_8603; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6565.4]
  wire  _T_8604; // @[Bitwise.scala 50:65:@6566.4]
  wire  _T_8605; // @[Bitwise.scala 50:65:@6567.4]
  wire  _T_8606; // @[Bitwise.scala 50:65:@6568.4]
  wire  _T_8607; // @[Bitwise.scala 50:65:@6569.4]
  wire  _T_8608; // @[Bitwise.scala 50:65:@6570.4]
  wire  _T_8609; // @[Bitwise.scala 50:65:@6571.4]
  wire  _T_8610; // @[Bitwise.scala 50:65:@6572.4]
  wire  _T_8611; // @[Bitwise.scala 50:65:@6573.4]
  wire  _T_8612; // @[Bitwise.scala 50:65:@6574.4]
  wire  _T_8613; // @[Bitwise.scala 50:65:@6575.4]
  wire  _T_8614; // @[Bitwise.scala 50:65:@6576.4]
  wire  _T_8615; // @[Bitwise.scala 50:65:@6577.4]
  wire  _T_8616; // @[Bitwise.scala 50:65:@6578.4]
  wire  _T_8617; // @[Bitwise.scala 50:65:@6579.4]
  wire  _T_8618; // @[Bitwise.scala 50:65:@6580.4]
  wire  _T_8619; // @[Bitwise.scala 50:65:@6581.4]
  wire  _T_8620; // @[Bitwise.scala 50:65:@6582.4]
  wire  _T_8621; // @[Bitwise.scala 50:65:@6583.4]
  wire  _T_8622; // @[Bitwise.scala 50:65:@6584.4]
  wire  _T_8623; // @[Bitwise.scala 50:65:@6585.4]
  wire  _T_8624; // @[Bitwise.scala 50:65:@6586.4]
  wire  _T_8625; // @[Bitwise.scala 50:65:@6587.4]
  wire  _T_8626; // @[Bitwise.scala 50:65:@6588.4]
  wire  _T_8627; // @[Bitwise.scala 50:65:@6589.4]
  wire  _T_8628; // @[Bitwise.scala 50:65:@6590.4]
  wire  _T_8629; // @[Bitwise.scala 50:65:@6591.4]
  wire  _T_8630; // @[Bitwise.scala 50:65:@6592.4]
  wire  _T_8631; // @[Bitwise.scala 50:65:@6593.4]
  wire  _T_8632; // @[Bitwise.scala 50:65:@6594.4]
  wire  _T_8633; // @[Bitwise.scala 50:65:@6595.4]
  wire  _T_8634; // @[Bitwise.scala 50:65:@6596.4]
  wire  _T_8635; // @[Bitwise.scala 50:65:@6597.4]
  wire  _T_8636; // @[Bitwise.scala 50:65:@6598.4]
  wire  _T_8637; // @[Bitwise.scala 50:65:@6599.4]
  wire  _T_8638; // @[Bitwise.scala 50:65:@6600.4]
  wire  _T_8639; // @[Bitwise.scala 50:65:@6601.4]
  wire  _T_8640; // @[Bitwise.scala 50:65:@6602.4]
  wire  _T_8641; // @[Bitwise.scala 50:65:@6603.4]
  wire  _T_8642; // @[Bitwise.scala 50:65:@6604.4]
  wire  _T_8643; // @[Bitwise.scala 50:65:@6605.4]
  wire  _T_8644; // @[Bitwise.scala 50:65:@6606.4]
  wire  _T_8645; // @[Bitwise.scala 50:65:@6607.4]
  wire  _T_8646; // @[Bitwise.scala 50:65:@6608.4]
  wire  _T_8647; // @[Bitwise.scala 50:65:@6609.4]
  wire  _T_8648; // @[Bitwise.scala 50:65:@6610.4]
  wire  _T_8649; // @[Bitwise.scala 50:65:@6611.4]
  wire  _T_8650; // @[Bitwise.scala 50:65:@6612.4]
  wire  _T_8651; // @[Bitwise.scala 50:65:@6613.4]
  wire  _T_8652; // @[Bitwise.scala 50:65:@6614.4]
  wire  _T_8653; // @[Bitwise.scala 50:65:@6615.4]
  wire  _T_8654; // @[Bitwise.scala 50:65:@6616.4]
  wire  _T_8655; // @[Bitwise.scala 50:65:@6617.4]
  wire  _T_8656; // @[Bitwise.scala 50:65:@6618.4]
  wire  _T_8657; // @[Bitwise.scala 50:65:@6619.4]
  wire  _T_8658; // @[Bitwise.scala 50:65:@6620.4]
  wire [1:0] _T_8659; // @[Bitwise.scala 48:55:@6621.4]
  wire [1:0] _GEN_952; // @[Bitwise.scala 48:55:@6622.4]
  wire [2:0] _T_8660; // @[Bitwise.scala 48:55:@6622.4]
  wire [1:0] _T_8661; // @[Bitwise.scala 48:55:@6623.4]
  wire [1:0] _GEN_953; // @[Bitwise.scala 48:55:@6624.4]
  wire [2:0] _T_8662; // @[Bitwise.scala 48:55:@6624.4]
  wire [3:0] _T_8663; // @[Bitwise.scala 48:55:@6625.4]
  wire [1:0] _T_8664; // @[Bitwise.scala 48:55:@6626.4]
  wire [1:0] _GEN_954; // @[Bitwise.scala 48:55:@6627.4]
  wire [2:0] _T_8665; // @[Bitwise.scala 48:55:@6627.4]
  wire [1:0] _T_8666; // @[Bitwise.scala 48:55:@6628.4]
  wire [1:0] _T_8667; // @[Bitwise.scala 48:55:@6629.4]
  wire [2:0] _T_8668; // @[Bitwise.scala 48:55:@6630.4]
  wire [3:0] _T_8669; // @[Bitwise.scala 48:55:@6631.4]
  wire [4:0] _T_8670; // @[Bitwise.scala 48:55:@6632.4]
  wire [1:0] _T_8671; // @[Bitwise.scala 48:55:@6633.4]
  wire [1:0] _GEN_955; // @[Bitwise.scala 48:55:@6634.4]
  wire [2:0] _T_8672; // @[Bitwise.scala 48:55:@6634.4]
  wire [1:0] _T_8673; // @[Bitwise.scala 48:55:@6635.4]
  wire [1:0] _T_8674; // @[Bitwise.scala 48:55:@6636.4]
  wire [2:0] _T_8675; // @[Bitwise.scala 48:55:@6637.4]
  wire [3:0] _T_8676; // @[Bitwise.scala 48:55:@6638.4]
  wire [1:0] _T_8677; // @[Bitwise.scala 48:55:@6639.4]
  wire [1:0] _GEN_956; // @[Bitwise.scala 48:55:@6640.4]
  wire [2:0] _T_8678; // @[Bitwise.scala 48:55:@6640.4]
  wire [1:0] _T_8679; // @[Bitwise.scala 48:55:@6641.4]
  wire [1:0] _T_8680; // @[Bitwise.scala 48:55:@6642.4]
  wire [2:0] _T_8681; // @[Bitwise.scala 48:55:@6643.4]
  wire [3:0] _T_8682; // @[Bitwise.scala 48:55:@6644.4]
  wire [4:0] _T_8683; // @[Bitwise.scala 48:55:@6645.4]
  wire [5:0] _T_8684; // @[Bitwise.scala 48:55:@6646.4]
  wire [1:0] _T_8685; // @[Bitwise.scala 48:55:@6647.4]
  wire [1:0] _GEN_957; // @[Bitwise.scala 48:55:@6648.4]
  wire [2:0] _T_8686; // @[Bitwise.scala 48:55:@6648.4]
  wire [1:0] _T_8687; // @[Bitwise.scala 48:55:@6649.4]
  wire [1:0] _T_8688; // @[Bitwise.scala 48:55:@6650.4]
  wire [2:0] _T_8689; // @[Bitwise.scala 48:55:@6651.4]
  wire [3:0] _T_8690; // @[Bitwise.scala 48:55:@6652.4]
  wire [1:0] _T_8691; // @[Bitwise.scala 48:55:@6653.4]
  wire [1:0] _GEN_958; // @[Bitwise.scala 48:55:@6654.4]
  wire [2:0] _T_8692; // @[Bitwise.scala 48:55:@6654.4]
  wire [1:0] _T_8693; // @[Bitwise.scala 48:55:@6655.4]
  wire [1:0] _T_8694; // @[Bitwise.scala 48:55:@6656.4]
  wire [2:0] _T_8695; // @[Bitwise.scala 48:55:@6657.4]
  wire [3:0] _T_8696; // @[Bitwise.scala 48:55:@6658.4]
  wire [4:0] _T_8697; // @[Bitwise.scala 48:55:@6659.4]
  wire [1:0] _T_8698; // @[Bitwise.scala 48:55:@6660.4]
  wire [1:0] _GEN_959; // @[Bitwise.scala 48:55:@6661.4]
  wire [2:0] _T_8699; // @[Bitwise.scala 48:55:@6661.4]
  wire [1:0] _T_8700; // @[Bitwise.scala 48:55:@6662.4]
  wire [1:0] _T_8701; // @[Bitwise.scala 48:55:@6663.4]
  wire [2:0] _T_8702; // @[Bitwise.scala 48:55:@6664.4]
  wire [3:0] _T_8703; // @[Bitwise.scala 48:55:@6665.4]
  wire [1:0] _T_8704; // @[Bitwise.scala 48:55:@6666.4]
  wire [1:0] _GEN_960; // @[Bitwise.scala 48:55:@6667.4]
  wire [2:0] _T_8705; // @[Bitwise.scala 48:55:@6667.4]
  wire [1:0] _T_8706; // @[Bitwise.scala 48:55:@6668.4]
  wire [1:0] _T_8707; // @[Bitwise.scala 48:55:@6669.4]
  wire [2:0] _T_8708; // @[Bitwise.scala 48:55:@6670.4]
  wire [3:0] _T_8709; // @[Bitwise.scala 48:55:@6671.4]
  wire [4:0] _T_8710; // @[Bitwise.scala 48:55:@6672.4]
  wire [5:0] _T_8711; // @[Bitwise.scala 48:55:@6673.4]
  wire [6:0] _T_8712; // @[Bitwise.scala 48:55:@6674.4]
  wire [55:0] _T_8776; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6739.4]
  wire  _T_8777; // @[Bitwise.scala 50:65:@6740.4]
  wire  _T_8778; // @[Bitwise.scala 50:65:@6741.4]
  wire  _T_8779; // @[Bitwise.scala 50:65:@6742.4]
  wire  _T_8780; // @[Bitwise.scala 50:65:@6743.4]
  wire  _T_8781; // @[Bitwise.scala 50:65:@6744.4]
  wire  _T_8782; // @[Bitwise.scala 50:65:@6745.4]
  wire  _T_8783; // @[Bitwise.scala 50:65:@6746.4]
  wire  _T_8784; // @[Bitwise.scala 50:65:@6747.4]
  wire  _T_8785; // @[Bitwise.scala 50:65:@6748.4]
  wire  _T_8786; // @[Bitwise.scala 50:65:@6749.4]
  wire  _T_8787; // @[Bitwise.scala 50:65:@6750.4]
  wire  _T_8788; // @[Bitwise.scala 50:65:@6751.4]
  wire  _T_8789; // @[Bitwise.scala 50:65:@6752.4]
  wire  _T_8790; // @[Bitwise.scala 50:65:@6753.4]
  wire  _T_8791; // @[Bitwise.scala 50:65:@6754.4]
  wire  _T_8792; // @[Bitwise.scala 50:65:@6755.4]
  wire  _T_8793; // @[Bitwise.scala 50:65:@6756.4]
  wire  _T_8794; // @[Bitwise.scala 50:65:@6757.4]
  wire  _T_8795; // @[Bitwise.scala 50:65:@6758.4]
  wire  _T_8796; // @[Bitwise.scala 50:65:@6759.4]
  wire  _T_8797; // @[Bitwise.scala 50:65:@6760.4]
  wire  _T_8798; // @[Bitwise.scala 50:65:@6761.4]
  wire  _T_8799; // @[Bitwise.scala 50:65:@6762.4]
  wire  _T_8800; // @[Bitwise.scala 50:65:@6763.4]
  wire  _T_8801; // @[Bitwise.scala 50:65:@6764.4]
  wire  _T_8802; // @[Bitwise.scala 50:65:@6765.4]
  wire  _T_8803; // @[Bitwise.scala 50:65:@6766.4]
  wire  _T_8804; // @[Bitwise.scala 50:65:@6767.4]
  wire  _T_8805; // @[Bitwise.scala 50:65:@6768.4]
  wire  _T_8806; // @[Bitwise.scala 50:65:@6769.4]
  wire  _T_8807; // @[Bitwise.scala 50:65:@6770.4]
  wire  _T_8808; // @[Bitwise.scala 50:65:@6771.4]
  wire  _T_8809; // @[Bitwise.scala 50:65:@6772.4]
  wire  _T_8810; // @[Bitwise.scala 50:65:@6773.4]
  wire  _T_8811; // @[Bitwise.scala 50:65:@6774.4]
  wire  _T_8812; // @[Bitwise.scala 50:65:@6775.4]
  wire  _T_8813; // @[Bitwise.scala 50:65:@6776.4]
  wire  _T_8814; // @[Bitwise.scala 50:65:@6777.4]
  wire  _T_8815; // @[Bitwise.scala 50:65:@6778.4]
  wire  _T_8816; // @[Bitwise.scala 50:65:@6779.4]
  wire  _T_8817; // @[Bitwise.scala 50:65:@6780.4]
  wire  _T_8818; // @[Bitwise.scala 50:65:@6781.4]
  wire  _T_8819; // @[Bitwise.scala 50:65:@6782.4]
  wire  _T_8820; // @[Bitwise.scala 50:65:@6783.4]
  wire  _T_8821; // @[Bitwise.scala 50:65:@6784.4]
  wire  _T_8822; // @[Bitwise.scala 50:65:@6785.4]
  wire  _T_8823; // @[Bitwise.scala 50:65:@6786.4]
  wire  _T_8824; // @[Bitwise.scala 50:65:@6787.4]
  wire  _T_8825; // @[Bitwise.scala 50:65:@6788.4]
  wire  _T_8826; // @[Bitwise.scala 50:65:@6789.4]
  wire  _T_8827; // @[Bitwise.scala 50:65:@6790.4]
  wire  _T_8828; // @[Bitwise.scala 50:65:@6791.4]
  wire  _T_8829; // @[Bitwise.scala 50:65:@6792.4]
  wire  _T_8830; // @[Bitwise.scala 50:65:@6793.4]
  wire  _T_8831; // @[Bitwise.scala 50:65:@6794.4]
  wire  _T_8832; // @[Bitwise.scala 50:65:@6795.4]
  wire [1:0] _T_8833; // @[Bitwise.scala 48:55:@6796.4]
  wire [1:0] _GEN_961; // @[Bitwise.scala 48:55:@6797.4]
  wire [2:0] _T_8834; // @[Bitwise.scala 48:55:@6797.4]
  wire [1:0] _T_8835; // @[Bitwise.scala 48:55:@6798.4]
  wire [1:0] _T_8836; // @[Bitwise.scala 48:55:@6799.4]
  wire [2:0] _T_8837; // @[Bitwise.scala 48:55:@6800.4]
  wire [3:0] _T_8838; // @[Bitwise.scala 48:55:@6801.4]
  wire [1:0] _T_8839; // @[Bitwise.scala 48:55:@6802.4]
  wire [1:0] _GEN_962; // @[Bitwise.scala 48:55:@6803.4]
  wire [2:0] _T_8840; // @[Bitwise.scala 48:55:@6803.4]
  wire [1:0] _T_8841; // @[Bitwise.scala 48:55:@6804.4]
  wire [1:0] _T_8842; // @[Bitwise.scala 48:55:@6805.4]
  wire [2:0] _T_8843; // @[Bitwise.scala 48:55:@6806.4]
  wire [3:0] _T_8844; // @[Bitwise.scala 48:55:@6807.4]
  wire [4:0] _T_8845; // @[Bitwise.scala 48:55:@6808.4]
  wire [1:0] _T_8846; // @[Bitwise.scala 48:55:@6809.4]
  wire [1:0] _GEN_963; // @[Bitwise.scala 48:55:@6810.4]
  wire [2:0] _T_8847; // @[Bitwise.scala 48:55:@6810.4]
  wire [1:0] _T_8848; // @[Bitwise.scala 48:55:@6811.4]
  wire [1:0] _T_8849; // @[Bitwise.scala 48:55:@6812.4]
  wire [2:0] _T_8850; // @[Bitwise.scala 48:55:@6813.4]
  wire [3:0] _T_8851; // @[Bitwise.scala 48:55:@6814.4]
  wire [1:0] _T_8852; // @[Bitwise.scala 48:55:@6815.4]
  wire [1:0] _GEN_964; // @[Bitwise.scala 48:55:@6816.4]
  wire [2:0] _T_8853; // @[Bitwise.scala 48:55:@6816.4]
  wire [1:0] _T_8854; // @[Bitwise.scala 48:55:@6817.4]
  wire [1:0] _T_8855; // @[Bitwise.scala 48:55:@6818.4]
  wire [2:0] _T_8856; // @[Bitwise.scala 48:55:@6819.4]
  wire [3:0] _T_8857; // @[Bitwise.scala 48:55:@6820.4]
  wire [4:0] _T_8858; // @[Bitwise.scala 48:55:@6821.4]
  wire [5:0] _T_8859; // @[Bitwise.scala 48:55:@6822.4]
  wire [1:0] _T_8860; // @[Bitwise.scala 48:55:@6823.4]
  wire [1:0] _GEN_965; // @[Bitwise.scala 48:55:@6824.4]
  wire [2:0] _T_8861; // @[Bitwise.scala 48:55:@6824.4]
  wire [1:0] _T_8862; // @[Bitwise.scala 48:55:@6825.4]
  wire [1:0] _T_8863; // @[Bitwise.scala 48:55:@6826.4]
  wire [2:0] _T_8864; // @[Bitwise.scala 48:55:@6827.4]
  wire [3:0] _T_8865; // @[Bitwise.scala 48:55:@6828.4]
  wire [1:0] _T_8866; // @[Bitwise.scala 48:55:@6829.4]
  wire [1:0] _GEN_966; // @[Bitwise.scala 48:55:@6830.4]
  wire [2:0] _T_8867; // @[Bitwise.scala 48:55:@6830.4]
  wire [1:0] _T_8868; // @[Bitwise.scala 48:55:@6831.4]
  wire [1:0] _T_8869; // @[Bitwise.scala 48:55:@6832.4]
  wire [2:0] _T_8870; // @[Bitwise.scala 48:55:@6833.4]
  wire [3:0] _T_8871; // @[Bitwise.scala 48:55:@6834.4]
  wire [4:0] _T_8872; // @[Bitwise.scala 48:55:@6835.4]
  wire [1:0] _T_8873; // @[Bitwise.scala 48:55:@6836.4]
  wire [1:0] _GEN_967; // @[Bitwise.scala 48:55:@6837.4]
  wire [2:0] _T_8874; // @[Bitwise.scala 48:55:@6837.4]
  wire [1:0] _T_8875; // @[Bitwise.scala 48:55:@6838.4]
  wire [1:0] _T_8876; // @[Bitwise.scala 48:55:@6839.4]
  wire [2:0] _T_8877; // @[Bitwise.scala 48:55:@6840.4]
  wire [3:0] _T_8878; // @[Bitwise.scala 48:55:@6841.4]
  wire [1:0] _T_8879; // @[Bitwise.scala 48:55:@6842.4]
  wire [1:0] _GEN_968; // @[Bitwise.scala 48:55:@6843.4]
  wire [2:0] _T_8880; // @[Bitwise.scala 48:55:@6843.4]
  wire [1:0] _T_8881; // @[Bitwise.scala 48:55:@6844.4]
  wire [1:0] _T_8882; // @[Bitwise.scala 48:55:@6845.4]
  wire [2:0] _T_8883; // @[Bitwise.scala 48:55:@6846.4]
  wire [3:0] _T_8884; // @[Bitwise.scala 48:55:@6847.4]
  wire [4:0] _T_8885; // @[Bitwise.scala 48:55:@6848.4]
  wire [5:0] _T_8886; // @[Bitwise.scala 48:55:@6849.4]
  wire [6:0] _T_8887; // @[Bitwise.scala 48:55:@6850.4]
  wire [56:0] _T_8951; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6915.4]
  wire  _T_8952; // @[Bitwise.scala 50:65:@6916.4]
  wire  _T_8953; // @[Bitwise.scala 50:65:@6917.4]
  wire  _T_8954; // @[Bitwise.scala 50:65:@6918.4]
  wire  _T_8955; // @[Bitwise.scala 50:65:@6919.4]
  wire  _T_8956; // @[Bitwise.scala 50:65:@6920.4]
  wire  _T_8957; // @[Bitwise.scala 50:65:@6921.4]
  wire  _T_8958; // @[Bitwise.scala 50:65:@6922.4]
  wire  _T_8959; // @[Bitwise.scala 50:65:@6923.4]
  wire  _T_8960; // @[Bitwise.scala 50:65:@6924.4]
  wire  _T_8961; // @[Bitwise.scala 50:65:@6925.4]
  wire  _T_8962; // @[Bitwise.scala 50:65:@6926.4]
  wire  _T_8963; // @[Bitwise.scala 50:65:@6927.4]
  wire  _T_8964; // @[Bitwise.scala 50:65:@6928.4]
  wire  _T_8965; // @[Bitwise.scala 50:65:@6929.4]
  wire  _T_8966; // @[Bitwise.scala 50:65:@6930.4]
  wire  _T_8967; // @[Bitwise.scala 50:65:@6931.4]
  wire  _T_8968; // @[Bitwise.scala 50:65:@6932.4]
  wire  _T_8969; // @[Bitwise.scala 50:65:@6933.4]
  wire  _T_8970; // @[Bitwise.scala 50:65:@6934.4]
  wire  _T_8971; // @[Bitwise.scala 50:65:@6935.4]
  wire  _T_8972; // @[Bitwise.scala 50:65:@6936.4]
  wire  _T_8973; // @[Bitwise.scala 50:65:@6937.4]
  wire  _T_8974; // @[Bitwise.scala 50:65:@6938.4]
  wire  _T_8975; // @[Bitwise.scala 50:65:@6939.4]
  wire  _T_8976; // @[Bitwise.scala 50:65:@6940.4]
  wire  _T_8977; // @[Bitwise.scala 50:65:@6941.4]
  wire  _T_8978; // @[Bitwise.scala 50:65:@6942.4]
  wire  _T_8979; // @[Bitwise.scala 50:65:@6943.4]
  wire  _T_8980; // @[Bitwise.scala 50:65:@6944.4]
  wire  _T_8981; // @[Bitwise.scala 50:65:@6945.4]
  wire  _T_8982; // @[Bitwise.scala 50:65:@6946.4]
  wire  _T_8983; // @[Bitwise.scala 50:65:@6947.4]
  wire  _T_8984; // @[Bitwise.scala 50:65:@6948.4]
  wire  _T_8985; // @[Bitwise.scala 50:65:@6949.4]
  wire  _T_8986; // @[Bitwise.scala 50:65:@6950.4]
  wire  _T_8987; // @[Bitwise.scala 50:65:@6951.4]
  wire  _T_8988; // @[Bitwise.scala 50:65:@6952.4]
  wire  _T_8989; // @[Bitwise.scala 50:65:@6953.4]
  wire  _T_8990; // @[Bitwise.scala 50:65:@6954.4]
  wire  _T_8991; // @[Bitwise.scala 50:65:@6955.4]
  wire  _T_8992; // @[Bitwise.scala 50:65:@6956.4]
  wire  _T_8993; // @[Bitwise.scala 50:65:@6957.4]
  wire  _T_8994; // @[Bitwise.scala 50:65:@6958.4]
  wire  _T_8995; // @[Bitwise.scala 50:65:@6959.4]
  wire  _T_8996; // @[Bitwise.scala 50:65:@6960.4]
  wire  _T_8997; // @[Bitwise.scala 50:65:@6961.4]
  wire  _T_8998; // @[Bitwise.scala 50:65:@6962.4]
  wire  _T_8999; // @[Bitwise.scala 50:65:@6963.4]
  wire  _T_9000; // @[Bitwise.scala 50:65:@6964.4]
  wire  _T_9001; // @[Bitwise.scala 50:65:@6965.4]
  wire  _T_9002; // @[Bitwise.scala 50:65:@6966.4]
  wire  _T_9003; // @[Bitwise.scala 50:65:@6967.4]
  wire  _T_9004; // @[Bitwise.scala 50:65:@6968.4]
  wire  _T_9005; // @[Bitwise.scala 50:65:@6969.4]
  wire  _T_9006; // @[Bitwise.scala 50:65:@6970.4]
  wire  _T_9007; // @[Bitwise.scala 50:65:@6971.4]
  wire  _T_9008; // @[Bitwise.scala 50:65:@6972.4]
  wire [1:0] _T_9009; // @[Bitwise.scala 48:55:@6973.4]
  wire [1:0] _GEN_969; // @[Bitwise.scala 48:55:@6974.4]
  wire [2:0] _T_9010; // @[Bitwise.scala 48:55:@6974.4]
  wire [1:0] _T_9011; // @[Bitwise.scala 48:55:@6975.4]
  wire [1:0] _T_9012; // @[Bitwise.scala 48:55:@6976.4]
  wire [2:0] _T_9013; // @[Bitwise.scala 48:55:@6977.4]
  wire [3:0] _T_9014; // @[Bitwise.scala 48:55:@6978.4]
  wire [1:0] _T_9015; // @[Bitwise.scala 48:55:@6979.4]
  wire [1:0] _GEN_970; // @[Bitwise.scala 48:55:@6980.4]
  wire [2:0] _T_9016; // @[Bitwise.scala 48:55:@6980.4]
  wire [1:0] _T_9017; // @[Bitwise.scala 48:55:@6981.4]
  wire [1:0] _T_9018; // @[Bitwise.scala 48:55:@6982.4]
  wire [2:0] _T_9019; // @[Bitwise.scala 48:55:@6983.4]
  wire [3:0] _T_9020; // @[Bitwise.scala 48:55:@6984.4]
  wire [4:0] _T_9021; // @[Bitwise.scala 48:55:@6985.4]
  wire [1:0] _T_9022; // @[Bitwise.scala 48:55:@6986.4]
  wire [1:0] _GEN_971; // @[Bitwise.scala 48:55:@6987.4]
  wire [2:0] _T_9023; // @[Bitwise.scala 48:55:@6987.4]
  wire [1:0] _T_9024; // @[Bitwise.scala 48:55:@6988.4]
  wire [1:0] _T_9025; // @[Bitwise.scala 48:55:@6989.4]
  wire [2:0] _T_9026; // @[Bitwise.scala 48:55:@6990.4]
  wire [3:0] _T_9027; // @[Bitwise.scala 48:55:@6991.4]
  wire [1:0] _T_9028; // @[Bitwise.scala 48:55:@6992.4]
  wire [1:0] _GEN_972; // @[Bitwise.scala 48:55:@6993.4]
  wire [2:0] _T_9029; // @[Bitwise.scala 48:55:@6993.4]
  wire [1:0] _T_9030; // @[Bitwise.scala 48:55:@6994.4]
  wire [1:0] _T_9031; // @[Bitwise.scala 48:55:@6995.4]
  wire [2:0] _T_9032; // @[Bitwise.scala 48:55:@6996.4]
  wire [3:0] _T_9033; // @[Bitwise.scala 48:55:@6997.4]
  wire [4:0] _T_9034; // @[Bitwise.scala 48:55:@6998.4]
  wire [5:0] _T_9035; // @[Bitwise.scala 48:55:@6999.4]
  wire [1:0] _T_9036; // @[Bitwise.scala 48:55:@7000.4]
  wire [1:0] _GEN_973; // @[Bitwise.scala 48:55:@7001.4]
  wire [2:0] _T_9037; // @[Bitwise.scala 48:55:@7001.4]
  wire [1:0] _T_9038; // @[Bitwise.scala 48:55:@7002.4]
  wire [1:0] _T_9039; // @[Bitwise.scala 48:55:@7003.4]
  wire [2:0] _T_9040; // @[Bitwise.scala 48:55:@7004.4]
  wire [3:0] _T_9041; // @[Bitwise.scala 48:55:@7005.4]
  wire [1:0] _T_9042; // @[Bitwise.scala 48:55:@7006.4]
  wire [1:0] _GEN_974; // @[Bitwise.scala 48:55:@7007.4]
  wire [2:0] _T_9043; // @[Bitwise.scala 48:55:@7007.4]
  wire [1:0] _T_9044; // @[Bitwise.scala 48:55:@7008.4]
  wire [1:0] _T_9045; // @[Bitwise.scala 48:55:@7009.4]
  wire [2:0] _T_9046; // @[Bitwise.scala 48:55:@7010.4]
  wire [3:0] _T_9047; // @[Bitwise.scala 48:55:@7011.4]
  wire [4:0] _T_9048; // @[Bitwise.scala 48:55:@7012.4]
  wire [1:0] _T_9049; // @[Bitwise.scala 48:55:@7013.4]
  wire [1:0] _GEN_975; // @[Bitwise.scala 48:55:@7014.4]
  wire [2:0] _T_9050; // @[Bitwise.scala 48:55:@7014.4]
  wire [1:0] _T_9051; // @[Bitwise.scala 48:55:@7015.4]
  wire [1:0] _T_9052; // @[Bitwise.scala 48:55:@7016.4]
  wire [2:0] _T_9053; // @[Bitwise.scala 48:55:@7017.4]
  wire [3:0] _T_9054; // @[Bitwise.scala 48:55:@7018.4]
  wire [1:0] _T_9055; // @[Bitwise.scala 48:55:@7019.4]
  wire [1:0] _T_9056; // @[Bitwise.scala 48:55:@7020.4]
  wire [2:0] _T_9057; // @[Bitwise.scala 48:55:@7021.4]
  wire [1:0] _T_9058; // @[Bitwise.scala 48:55:@7022.4]
  wire [1:0] _T_9059; // @[Bitwise.scala 48:55:@7023.4]
  wire [2:0] _T_9060; // @[Bitwise.scala 48:55:@7024.4]
  wire [3:0] _T_9061; // @[Bitwise.scala 48:55:@7025.4]
  wire [4:0] _T_9062; // @[Bitwise.scala 48:55:@7026.4]
  wire [5:0] _T_9063; // @[Bitwise.scala 48:55:@7027.4]
  wire [6:0] _T_9064; // @[Bitwise.scala 48:55:@7028.4]
  wire [57:0] _T_9128; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7093.4]
  wire  _T_9129; // @[Bitwise.scala 50:65:@7094.4]
  wire  _T_9130; // @[Bitwise.scala 50:65:@7095.4]
  wire  _T_9131; // @[Bitwise.scala 50:65:@7096.4]
  wire  _T_9132; // @[Bitwise.scala 50:65:@7097.4]
  wire  _T_9133; // @[Bitwise.scala 50:65:@7098.4]
  wire  _T_9134; // @[Bitwise.scala 50:65:@7099.4]
  wire  _T_9135; // @[Bitwise.scala 50:65:@7100.4]
  wire  _T_9136; // @[Bitwise.scala 50:65:@7101.4]
  wire  _T_9137; // @[Bitwise.scala 50:65:@7102.4]
  wire  _T_9138; // @[Bitwise.scala 50:65:@7103.4]
  wire  _T_9139; // @[Bitwise.scala 50:65:@7104.4]
  wire  _T_9140; // @[Bitwise.scala 50:65:@7105.4]
  wire  _T_9141; // @[Bitwise.scala 50:65:@7106.4]
  wire  _T_9142; // @[Bitwise.scala 50:65:@7107.4]
  wire  _T_9143; // @[Bitwise.scala 50:65:@7108.4]
  wire  _T_9144; // @[Bitwise.scala 50:65:@7109.4]
  wire  _T_9145; // @[Bitwise.scala 50:65:@7110.4]
  wire  _T_9146; // @[Bitwise.scala 50:65:@7111.4]
  wire  _T_9147; // @[Bitwise.scala 50:65:@7112.4]
  wire  _T_9148; // @[Bitwise.scala 50:65:@7113.4]
  wire  _T_9149; // @[Bitwise.scala 50:65:@7114.4]
  wire  _T_9150; // @[Bitwise.scala 50:65:@7115.4]
  wire  _T_9151; // @[Bitwise.scala 50:65:@7116.4]
  wire  _T_9152; // @[Bitwise.scala 50:65:@7117.4]
  wire  _T_9153; // @[Bitwise.scala 50:65:@7118.4]
  wire  _T_9154; // @[Bitwise.scala 50:65:@7119.4]
  wire  _T_9155; // @[Bitwise.scala 50:65:@7120.4]
  wire  _T_9156; // @[Bitwise.scala 50:65:@7121.4]
  wire  _T_9157; // @[Bitwise.scala 50:65:@7122.4]
  wire  _T_9158; // @[Bitwise.scala 50:65:@7123.4]
  wire  _T_9159; // @[Bitwise.scala 50:65:@7124.4]
  wire  _T_9160; // @[Bitwise.scala 50:65:@7125.4]
  wire  _T_9161; // @[Bitwise.scala 50:65:@7126.4]
  wire  _T_9162; // @[Bitwise.scala 50:65:@7127.4]
  wire  _T_9163; // @[Bitwise.scala 50:65:@7128.4]
  wire  _T_9164; // @[Bitwise.scala 50:65:@7129.4]
  wire  _T_9165; // @[Bitwise.scala 50:65:@7130.4]
  wire  _T_9166; // @[Bitwise.scala 50:65:@7131.4]
  wire  _T_9167; // @[Bitwise.scala 50:65:@7132.4]
  wire  _T_9168; // @[Bitwise.scala 50:65:@7133.4]
  wire  _T_9169; // @[Bitwise.scala 50:65:@7134.4]
  wire  _T_9170; // @[Bitwise.scala 50:65:@7135.4]
  wire  _T_9171; // @[Bitwise.scala 50:65:@7136.4]
  wire  _T_9172; // @[Bitwise.scala 50:65:@7137.4]
  wire  _T_9173; // @[Bitwise.scala 50:65:@7138.4]
  wire  _T_9174; // @[Bitwise.scala 50:65:@7139.4]
  wire  _T_9175; // @[Bitwise.scala 50:65:@7140.4]
  wire  _T_9176; // @[Bitwise.scala 50:65:@7141.4]
  wire  _T_9177; // @[Bitwise.scala 50:65:@7142.4]
  wire  _T_9178; // @[Bitwise.scala 50:65:@7143.4]
  wire  _T_9179; // @[Bitwise.scala 50:65:@7144.4]
  wire  _T_9180; // @[Bitwise.scala 50:65:@7145.4]
  wire  _T_9181; // @[Bitwise.scala 50:65:@7146.4]
  wire  _T_9182; // @[Bitwise.scala 50:65:@7147.4]
  wire  _T_9183; // @[Bitwise.scala 50:65:@7148.4]
  wire  _T_9184; // @[Bitwise.scala 50:65:@7149.4]
  wire  _T_9185; // @[Bitwise.scala 50:65:@7150.4]
  wire  _T_9186; // @[Bitwise.scala 50:65:@7151.4]
  wire [1:0] _T_9187; // @[Bitwise.scala 48:55:@7152.4]
  wire [1:0] _GEN_976; // @[Bitwise.scala 48:55:@7153.4]
  wire [2:0] _T_9188; // @[Bitwise.scala 48:55:@7153.4]
  wire [1:0] _T_9189; // @[Bitwise.scala 48:55:@7154.4]
  wire [1:0] _T_9190; // @[Bitwise.scala 48:55:@7155.4]
  wire [2:0] _T_9191; // @[Bitwise.scala 48:55:@7156.4]
  wire [3:0] _T_9192; // @[Bitwise.scala 48:55:@7157.4]
  wire [1:0] _T_9193; // @[Bitwise.scala 48:55:@7158.4]
  wire [1:0] _GEN_977; // @[Bitwise.scala 48:55:@7159.4]
  wire [2:0] _T_9194; // @[Bitwise.scala 48:55:@7159.4]
  wire [1:0] _T_9195; // @[Bitwise.scala 48:55:@7160.4]
  wire [1:0] _T_9196; // @[Bitwise.scala 48:55:@7161.4]
  wire [2:0] _T_9197; // @[Bitwise.scala 48:55:@7162.4]
  wire [3:0] _T_9198; // @[Bitwise.scala 48:55:@7163.4]
  wire [4:0] _T_9199; // @[Bitwise.scala 48:55:@7164.4]
  wire [1:0] _T_9200; // @[Bitwise.scala 48:55:@7165.4]
  wire [1:0] _GEN_978; // @[Bitwise.scala 48:55:@7166.4]
  wire [2:0] _T_9201; // @[Bitwise.scala 48:55:@7166.4]
  wire [1:0] _T_9202; // @[Bitwise.scala 48:55:@7167.4]
  wire [1:0] _T_9203; // @[Bitwise.scala 48:55:@7168.4]
  wire [2:0] _T_9204; // @[Bitwise.scala 48:55:@7169.4]
  wire [3:0] _T_9205; // @[Bitwise.scala 48:55:@7170.4]
  wire [1:0] _T_9206; // @[Bitwise.scala 48:55:@7171.4]
  wire [1:0] _T_9207; // @[Bitwise.scala 48:55:@7172.4]
  wire [2:0] _T_9208; // @[Bitwise.scala 48:55:@7173.4]
  wire [1:0] _T_9209; // @[Bitwise.scala 48:55:@7174.4]
  wire [1:0] _T_9210; // @[Bitwise.scala 48:55:@7175.4]
  wire [2:0] _T_9211; // @[Bitwise.scala 48:55:@7176.4]
  wire [3:0] _T_9212; // @[Bitwise.scala 48:55:@7177.4]
  wire [4:0] _T_9213; // @[Bitwise.scala 48:55:@7178.4]
  wire [5:0] _T_9214; // @[Bitwise.scala 48:55:@7179.4]
  wire [1:0] _T_9215; // @[Bitwise.scala 48:55:@7180.4]
  wire [1:0] _GEN_979; // @[Bitwise.scala 48:55:@7181.4]
  wire [2:0] _T_9216; // @[Bitwise.scala 48:55:@7181.4]
  wire [1:0] _T_9217; // @[Bitwise.scala 48:55:@7182.4]
  wire [1:0] _T_9218; // @[Bitwise.scala 48:55:@7183.4]
  wire [2:0] _T_9219; // @[Bitwise.scala 48:55:@7184.4]
  wire [3:0] _T_9220; // @[Bitwise.scala 48:55:@7185.4]
  wire [1:0] _T_9221; // @[Bitwise.scala 48:55:@7186.4]
  wire [1:0] _GEN_980; // @[Bitwise.scala 48:55:@7187.4]
  wire [2:0] _T_9222; // @[Bitwise.scala 48:55:@7187.4]
  wire [1:0] _T_9223; // @[Bitwise.scala 48:55:@7188.4]
  wire [1:0] _T_9224; // @[Bitwise.scala 48:55:@7189.4]
  wire [2:0] _T_9225; // @[Bitwise.scala 48:55:@7190.4]
  wire [3:0] _T_9226; // @[Bitwise.scala 48:55:@7191.4]
  wire [4:0] _T_9227; // @[Bitwise.scala 48:55:@7192.4]
  wire [1:0] _T_9228; // @[Bitwise.scala 48:55:@7193.4]
  wire [1:0] _GEN_981; // @[Bitwise.scala 48:55:@7194.4]
  wire [2:0] _T_9229; // @[Bitwise.scala 48:55:@7194.4]
  wire [1:0] _T_9230; // @[Bitwise.scala 48:55:@7195.4]
  wire [1:0] _T_9231; // @[Bitwise.scala 48:55:@7196.4]
  wire [2:0] _T_9232; // @[Bitwise.scala 48:55:@7197.4]
  wire [3:0] _T_9233; // @[Bitwise.scala 48:55:@7198.4]
  wire [1:0] _T_9234; // @[Bitwise.scala 48:55:@7199.4]
  wire [1:0] _T_9235; // @[Bitwise.scala 48:55:@7200.4]
  wire [2:0] _T_9236; // @[Bitwise.scala 48:55:@7201.4]
  wire [1:0] _T_9237; // @[Bitwise.scala 48:55:@7202.4]
  wire [1:0] _T_9238; // @[Bitwise.scala 48:55:@7203.4]
  wire [2:0] _T_9239; // @[Bitwise.scala 48:55:@7204.4]
  wire [3:0] _T_9240; // @[Bitwise.scala 48:55:@7205.4]
  wire [4:0] _T_9241; // @[Bitwise.scala 48:55:@7206.4]
  wire [5:0] _T_9242; // @[Bitwise.scala 48:55:@7207.4]
  wire [6:0] _T_9243; // @[Bitwise.scala 48:55:@7208.4]
  wire [58:0] _T_9307; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7273.4]
  wire  _T_9308; // @[Bitwise.scala 50:65:@7274.4]
  wire  _T_9309; // @[Bitwise.scala 50:65:@7275.4]
  wire  _T_9310; // @[Bitwise.scala 50:65:@7276.4]
  wire  _T_9311; // @[Bitwise.scala 50:65:@7277.4]
  wire  _T_9312; // @[Bitwise.scala 50:65:@7278.4]
  wire  _T_9313; // @[Bitwise.scala 50:65:@7279.4]
  wire  _T_9314; // @[Bitwise.scala 50:65:@7280.4]
  wire  _T_9315; // @[Bitwise.scala 50:65:@7281.4]
  wire  _T_9316; // @[Bitwise.scala 50:65:@7282.4]
  wire  _T_9317; // @[Bitwise.scala 50:65:@7283.4]
  wire  _T_9318; // @[Bitwise.scala 50:65:@7284.4]
  wire  _T_9319; // @[Bitwise.scala 50:65:@7285.4]
  wire  _T_9320; // @[Bitwise.scala 50:65:@7286.4]
  wire  _T_9321; // @[Bitwise.scala 50:65:@7287.4]
  wire  _T_9322; // @[Bitwise.scala 50:65:@7288.4]
  wire  _T_9323; // @[Bitwise.scala 50:65:@7289.4]
  wire  _T_9324; // @[Bitwise.scala 50:65:@7290.4]
  wire  _T_9325; // @[Bitwise.scala 50:65:@7291.4]
  wire  _T_9326; // @[Bitwise.scala 50:65:@7292.4]
  wire  _T_9327; // @[Bitwise.scala 50:65:@7293.4]
  wire  _T_9328; // @[Bitwise.scala 50:65:@7294.4]
  wire  _T_9329; // @[Bitwise.scala 50:65:@7295.4]
  wire  _T_9330; // @[Bitwise.scala 50:65:@7296.4]
  wire  _T_9331; // @[Bitwise.scala 50:65:@7297.4]
  wire  _T_9332; // @[Bitwise.scala 50:65:@7298.4]
  wire  _T_9333; // @[Bitwise.scala 50:65:@7299.4]
  wire  _T_9334; // @[Bitwise.scala 50:65:@7300.4]
  wire  _T_9335; // @[Bitwise.scala 50:65:@7301.4]
  wire  _T_9336; // @[Bitwise.scala 50:65:@7302.4]
  wire  _T_9337; // @[Bitwise.scala 50:65:@7303.4]
  wire  _T_9338; // @[Bitwise.scala 50:65:@7304.4]
  wire  _T_9339; // @[Bitwise.scala 50:65:@7305.4]
  wire  _T_9340; // @[Bitwise.scala 50:65:@7306.4]
  wire  _T_9341; // @[Bitwise.scala 50:65:@7307.4]
  wire  _T_9342; // @[Bitwise.scala 50:65:@7308.4]
  wire  _T_9343; // @[Bitwise.scala 50:65:@7309.4]
  wire  _T_9344; // @[Bitwise.scala 50:65:@7310.4]
  wire  _T_9345; // @[Bitwise.scala 50:65:@7311.4]
  wire  _T_9346; // @[Bitwise.scala 50:65:@7312.4]
  wire  _T_9347; // @[Bitwise.scala 50:65:@7313.4]
  wire  _T_9348; // @[Bitwise.scala 50:65:@7314.4]
  wire  _T_9349; // @[Bitwise.scala 50:65:@7315.4]
  wire  _T_9350; // @[Bitwise.scala 50:65:@7316.4]
  wire  _T_9351; // @[Bitwise.scala 50:65:@7317.4]
  wire  _T_9352; // @[Bitwise.scala 50:65:@7318.4]
  wire  _T_9353; // @[Bitwise.scala 50:65:@7319.4]
  wire  _T_9354; // @[Bitwise.scala 50:65:@7320.4]
  wire  _T_9355; // @[Bitwise.scala 50:65:@7321.4]
  wire  _T_9356; // @[Bitwise.scala 50:65:@7322.4]
  wire  _T_9357; // @[Bitwise.scala 50:65:@7323.4]
  wire  _T_9358; // @[Bitwise.scala 50:65:@7324.4]
  wire  _T_9359; // @[Bitwise.scala 50:65:@7325.4]
  wire  _T_9360; // @[Bitwise.scala 50:65:@7326.4]
  wire  _T_9361; // @[Bitwise.scala 50:65:@7327.4]
  wire  _T_9362; // @[Bitwise.scala 50:65:@7328.4]
  wire  _T_9363; // @[Bitwise.scala 50:65:@7329.4]
  wire  _T_9364; // @[Bitwise.scala 50:65:@7330.4]
  wire  _T_9365; // @[Bitwise.scala 50:65:@7331.4]
  wire  _T_9366; // @[Bitwise.scala 50:65:@7332.4]
  wire [1:0] _T_9367; // @[Bitwise.scala 48:55:@7333.4]
  wire [1:0] _GEN_982; // @[Bitwise.scala 48:55:@7334.4]
  wire [2:0] _T_9368; // @[Bitwise.scala 48:55:@7334.4]
  wire [1:0] _T_9369; // @[Bitwise.scala 48:55:@7335.4]
  wire [1:0] _T_9370; // @[Bitwise.scala 48:55:@7336.4]
  wire [2:0] _T_9371; // @[Bitwise.scala 48:55:@7337.4]
  wire [3:0] _T_9372; // @[Bitwise.scala 48:55:@7338.4]
  wire [1:0] _T_9373; // @[Bitwise.scala 48:55:@7339.4]
  wire [1:0] _GEN_983; // @[Bitwise.scala 48:55:@7340.4]
  wire [2:0] _T_9374; // @[Bitwise.scala 48:55:@7340.4]
  wire [1:0] _T_9375; // @[Bitwise.scala 48:55:@7341.4]
  wire [1:0] _T_9376; // @[Bitwise.scala 48:55:@7342.4]
  wire [2:0] _T_9377; // @[Bitwise.scala 48:55:@7343.4]
  wire [3:0] _T_9378; // @[Bitwise.scala 48:55:@7344.4]
  wire [4:0] _T_9379; // @[Bitwise.scala 48:55:@7345.4]
  wire [1:0] _T_9380; // @[Bitwise.scala 48:55:@7346.4]
  wire [1:0] _GEN_984; // @[Bitwise.scala 48:55:@7347.4]
  wire [2:0] _T_9381; // @[Bitwise.scala 48:55:@7347.4]
  wire [1:0] _T_9382; // @[Bitwise.scala 48:55:@7348.4]
  wire [1:0] _T_9383; // @[Bitwise.scala 48:55:@7349.4]
  wire [2:0] _T_9384; // @[Bitwise.scala 48:55:@7350.4]
  wire [3:0] _T_9385; // @[Bitwise.scala 48:55:@7351.4]
  wire [1:0] _T_9386; // @[Bitwise.scala 48:55:@7352.4]
  wire [1:0] _T_9387; // @[Bitwise.scala 48:55:@7353.4]
  wire [2:0] _T_9388; // @[Bitwise.scala 48:55:@7354.4]
  wire [1:0] _T_9389; // @[Bitwise.scala 48:55:@7355.4]
  wire [1:0] _T_9390; // @[Bitwise.scala 48:55:@7356.4]
  wire [2:0] _T_9391; // @[Bitwise.scala 48:55:@7357.4]
  wire [3:0] _T_9392; // @[Bitwise.scala 48:55:@7358.4]
  wire [4:0] _T_9393; // @[Bitwise.scala 48:55:@7359.4]
  wire [5:0] _T_9394; // @[Bitwise.scala 48:55:@7360.4]
  wire [1:0] _T_9395; // @[Bitwise.scala 48:55:@7361.4]
  wire [1:0] _GEN_985; // @[Bitwise.scala 48:55:@7362.4]
  wire [2:0] _T_9396; // @[Bitwise.scala 48:55:@7362.4]
  wire [1:0] _T_9397; // @[Bitwise.scala 48:55:@7363.4]
  wire [1:0] _T_9398; // @[Bitwise.scala 48:55:@7364.4]
  wire [2:0] _T_9399; // @[Bitwise.scala 48:55:@7365.4]
  wire [3:0] _T_9400; // @[Bitwise.scala 48:55:@7366.4]
  wire [1:0] _T_9401; // @[Bitwise.scala 48:55:@7367.4]
  wire [1:0] _T_9402; // @[Bitwise.scala 48:55:@7368.4]
  wire [2:0] _T_9403; // @[Bitwise.scala 48:55:@7369.4]
  wire [1:0] _T_9404; // @[Bitwise.scala 48:55:@7370.4]
  wire [1:0] _T_9405; // @[Bitwise.scala 48:55:@7371.4]
  wire [2:0] _T_9406; // @[Bitwise.scala 48:55:@7372.4]
  wire [3:0] _T_9407; // @[Bitwise.scala 48:55:@7373.4]
  wire [4:0] _T_9408; // @[Bitwise.scala 48:55:@7374.4]
  wire [1:0] _T_9409; // @[Bitwise.scala 48:55:@7375.4]
  wire [1:0] _GEN_986; // @[Bitwise.scala 48:55:@7376.4]
  wire [2:0] _T_9410; // @[Bitwise.scala 48:55:@7376.4]
  wire [1:0] _T_9411; // @[Bitwise.scala 48:55:@7377.4]
  wire [1:0] _T_9412; // @[Bitwise.scala 48:55:@7378.4]
  wire [2:0] _T_9413; // @[Bitwise.scala 48:55:@7379.4]
  wire [3:0] _T_9414; // @[Bitwise.scala 48:55:@7380.4]
  wire [1:0] _T_9415; // @[Bitwise.scala 48:55:@7381.4]
  wire [1:0] _T_9416; // @[Bitwise.scala 48:55:@7382.4]
  wire [2:0] _T_9417; // @[Bitwise.scala 48:55:@7383.4]
  wire [1:0] _T_9418; // @[Bitwise.scala 48:55:@7384.4]
  wire [1:0] _T_9419; // @[Bitwise.scala 48:55:@7385.4]
  wire [2:0] _T_9420; // @[Bitwise.scala 48:55:@7386.4]
  wire [3:0] _T_9421; // @[Bitwise.scala 48:55:@7387.4]
  wire [4:0] _T_9422; // @[Bitwise.scala 48:55:@7388.4]
  wire [5:0] _T_9423; // @[Bitwise.scala 48:55:@7389.4]
  wire [6:0] _T_9424; // @[Bitwise.scala 48:55:@7390.4]
  wire [59:0] _T_9488; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7455.4]
  wire  _T_9489; // @[Bitwise.scala 50:65:@7456.4]
  wire  _T_9490; // @[Bitwise.scala 50:65:@7457.4]
  wire  _T_9491; // @[Bitwise.scala 50:65:@7458.4]
  wire  _T_9492; // @[Bitwise.scala 50:65:@7459.4]
  wire  _T_9493; // @[Bitwise.scala 50:65:@7460.4]
  wire  _T_9494; // @[Bitwise.scala 50:65:@7461.4]
  wire  _T_9495; // @[Bitwise.scala 50:65:@7462.4]
  wire  _T_9496; // @[Bitwise.scala 50:65:@7463.4]
  wire  _T_9497; // @[Bitwise.scala 50:65:@7464.4]
  wire  _T_9498; // @[Bitwise.scala 50:65:@7465.4]
  wire  _T_9499; // @[Bitwise.scala 50:65:@7466.4]
  wire  _T_9500; // @[Bitwise.scala 50:65:@7467.4]
  wire  _T_9501; // @[Bitwise.scala 50:65:@7468.4]
  wire  _T_9502; // @[Bitwise.scala 50:65:@7469.4]
  wire  _T_9503; // @[Bitwise.scala 50:65:@7470.4]
  wire  _T_9504; // @[Bitwise.scala 50:65:@7471.4]
  wire  _T_9505; // @[Bitwise.scala 50:65:@7472.4]
  wire  _T_9506; // @[Bitwise.scala 50:65:@7473.4]
  wire  _T_9507; // @[Bitwise.scala 50:65:@7474.4]
  wire  _T_9508; // @[Bitwise.scala 50:65:@7475.4]
  wire  _T_9509; // @[Bitwise.scala 50:65:@7476.4]
  wire  _T_9510; // @[Bitwise.scala 50:65:@7477.4]
  wire  _T_9511; // @[Bitwise.scala 50:65:@7478.4]
  wire  _T_9512; // @[Bitwise.scala 50:65:@7479.4]
  wire  _T_9513; // @[Bitwise.scala 50:65:@7480.4]
  wire  _T_9514; // @[Bitwise.scala 50:65:@7481.4]
  wire  _T_9515; // @[Bitwise.scala 50:65:@7482.4]
  wire  _T_9516; // @[Bitwise.scala 50:65:@7483.4]
  wire  _T_9517; // @[Bitwise.scala 50:65:@7484.4]
  wire  _T_9518; // @[Bitwise.scala 50:65:@7485.4]
  wire  _T_9519; // @[Bitwise.scala 50:65:@7486.4]
  wire  _T_9520; // @[Bitwise.scala 50:65:@7487.4]
  wire  _T_9521; // @[Bitwise.scala 50:65:@7488.4]
  wire  _T_9522; // @[Bitwise.scala 50:65:@7489.4]
  wire  _T_9523; // @[Bitwise.scala 50:65:@7490.4]
  wire  _T_9524; // @[Bitwise.scala 50:65:@7491.4]
  wire  _T_9525; // @[Bitwise.scala 50:65:@7492.4]
  wire  _T_9526; // @[Bitwise.scala 50:65:@7493.4]
  wire  _T_9527; // @[Bitwise.scala 50:65:@7494.4]
  wire  _T_9528; // @[Bitwise.scala 50:65:@7495.4]
  wire  _T_9529; // @[Bitwise.scala 50:65:@7496.4]
  wire  _T_9530; // @[Bitwise.scala 50:65:@7497.4]
  wire  _T_9531; // @[Bitwise.scala 50:65:@7498.4]
  wire  _T_9532; // @[Bitwise.scala 50:65:@7499.4]
  wire  _T_9533; // @[Bitwise.scala 50:65:@7500.4]
  wire  _T_9534; // @[Bitwise.scala 50:65:@7501.4]
  wire  _T_9535; // @[Bitwise.scala 50:65:@7502.4]
  wire  _T_9536; // @[Bitwise.scala 50:65:@7503.4]
  wire  _T_9537; // @[Bitwise.scala 50:65:@7504.4]
  wire  _T_9538; // @[Bitwise.scala 50:65:@7505.4]
  wire  _T_9539; // @[Bitwise.scala 50:65:@7506.4]
  wire  _T_9540; // @[Bitwise.scala 50:65:@7507.4]
  wire  _T_9541; // @[Bitwise.scala 50:65:@7508.4]
  wire  _T_9542; // @[Bitwise.scala 50:65:@7509.4]
  wire  _T_9543; // @[Bitwise.scala 50:65:@7510.4]
  wire  _T_9544; // @[Bitwise.scala 50:65:@7511.4]
  wire  _T_9545; // @[Bitwise.scala 50:65:@7512.4]
  wire  _T_9546; // @[Bitwise.scala 50:65:@7513.4]
  wire  _T_9547; // @[Bitwise.scala 50:65:@7514.4]
  wire  _T_9548; // @[Bitwise.scala 50:65:@7515.4]
  wire [1:0] _T_9549; // @[Bitwise.scala 48:55:@7516.4]
  wire [1:0] _GEN_987; // @[Bitwise.scala 48:55:@7517.4]
  wire [2:0] _T_9550; // @[Bitwise.scala 48:55:@7517.4]
  wire [1:0] _T_9551; // @[Bitwise.scala 48:55:@7518.4]
  wire [1:0] _T_9552; // @[Bitwise.scala 48:55:@7519.4]
  wire [2:0] _T_9553; // @[Bitwise.scala 48:55:@7520.4]
  wire [3:0] _T_9554; // @[Bitwise.scala 48:55:@7521.4]
  wire [1:0] _T_9555; // @[Bitwise.scala 48:55:@7522.4]
  wire [1:0] _T_9556; // @[Bitwise.scala 48:55:@7523.4]
  wire [2:0] _T_9557; // @[Bitwise.scala 48:55:@7524.4]
  wire [1:0] _T_9558; // @[Bitwise.scala 48:55:@7525.4]
  wire [1:0] _T_9559; // @[Bitwise.scala 48:55:@7526.4]
  wire [2:0] _T_9560; // @[Bitwise.scala 48:55:@7527.4]
  wire [3:0] _T_9561; // @[Bitwise.scala 48:55:@7528.4]
  wire [4:0] _T_9562; // @[Bitwise.scala 48:55:@7529.4]
  wire [1:0] _T_9563; // @[Bitwise.scala 48:55:@7530.4]
  wire [1:0] _GEN_988; // @[Bitwise.scala 48:55:@7531.4]
  wire [2:0] _T_9564; // @[Bitwise.scala 48:55:@7531.4]
  wire [1:0] _T_9565; // @[Bitwise.scala 48:55:@7532.4]
  wire [1:0] _T_9566; // @[Bitwise.scala 48:55:@7533.4]
  wire [2:0] _T_9567; // @[Bitwise.scala 48:55:@7534.4]
  wire [3:0] _T_9568; // @[Bitwise.scala 48:55:@7535.4]
  wire [1:0] _T_9569; // @[Bitwise.scala 48:55:@7536.4]
  wire [1:0] _T_9570; // @[Bitwise.scala 48:55:@7537.4]
  wire [2:0] _T_9571; // @[Bitwise.scala 48:55:@7538.4]
  wire [1:0] _T_9572; // @[Bitwise.scala 48:55:@7539.4]
  wire [1:0] _T_9573; // @[Bitwise.scala 48:55:@7540.4]
  wire [2:0] _T_9574; // @[Bitwise.scala 48:55:@7541.4]
  wire [3:0] _T_9575; // @[Bitwise.scala 48:55:@7542.4]
  wire [4:0] _T_9576; // @[Bitwise.scala 48:55:@7543.4]
  wire [5:0] _T_9577; // @[Bitwise.scala 48:55:@7544.4]
  wire [1:0] _T_9578; // @[Bitwise.scala 48:55:@7545.4]
  wire [1:0] _GEN_989; // @[Bitwise.scala 48:55:@7546.4]
  wire [2:0] _T_9579; // @[Bitwise.scala 48:55:@7546.4]
  wire [1:0] _T_9580; // @[Bitwise.scala 48:55:@7547.4]
  wire [1:0] _T_9581; // @[Bitwise.scala 48:55:@7548.4]
  wire [2:0] _T_9582; // @[Bitwise.scala 48:55:@7549.4]
  wire [3:0] _T_9583; // @[Bitwise.scala 48:55:@7550.4]
  wire [1:0] _T_9584; // @[Bitwise.scala 48:55:@7551.4]
  wire [1:0] _T_9585; // @[Bitwise.scala 48:55:@7552.4]
  wire [2:0] _T_9586; // @[Bitwise.scala 48:55:@7553.4]
  wire [1:0] _T_9587; // @[Bitwise.scala 48:55:@7554.4]
  wire [1:0] _T_9588; // @[Bitwise.scala 48:55:@7555.4]
  wire [2:0] _T_9589; // @[Bitwise.scala 48:55:@7556.4]
  wire [3:0] _T_9590; // @[Bitwise.scala 48:55:@7557.4]
  wire [4:0] _T_9591; // @[Bitwise.scala 48:55:@7558.4]
  wire [1:0] _T_9592; // @[Bitwise.scala 48:55:@7559.4]
  wire [1:0] _GEN_990; // @[Bitwise.scala 48:55:@7560.4]
  wire [2:0] _T_9593; // @[Bitwise.scala 48:55:@7560.4]
  wire [1:0] _T_9594; // @[Bitwise.scala 48:55:@7561.4]
  wire [1:0] _T_9595; // @[Bitwise.scala 48:55:@7562.4]
  wire [2:0] _T_9596; // @[Bitwise.scala 48:55:@7563.4]
  wire [3:0] _T_9597; // @[Bitwise.scala 48:55:@7564.4]
  wire [1:0] _T_9598; // @[Bitwise.scala 48:55:@7565.4]
  wire [1:0] _T_9599; // @[Bitwise.scala 48:55:@7566.4]
  wire [2:0] _T_9600; // @[Bitwise.scala 48:55:@7567.4]
  wire [1:0] _T_9601; // @[Bitwise.scala 48:55:@7568.4]
  wire [1:0] _T_9602; // @[Bitwise.scala 48:55:@7569.4]
  wire [2:0] _T_9603; // @[Bitwise.scala 48:55:@7570.4]
  wire [3:0] _T_9604; // @[Bitwise.scala 48:55:@7571.4]
  wire [4:0] _T_9605; // @[Bitwise.scala 48:55:@7572.4]
  wire [5:0] _T_9606; // @[Bitwise.scala 48:55:@7573.4]
  wire [6:0] _T_9607; // @[Bitwise.scala 48:55:@7574.4]
  wire [60:0] _T_9671; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7639.4]
  wire  _T_9672; // @[Bitwise.scala 50:65:@7640.4]
  wire  _T_9673; // @[Bitwise.scala 50:65:@7641.4]
  wire  _T_9674; // @[Bitwise.scala 50:65:@7642.4]
  wire  _T_9675; // @[Bitwise.scala 50:65:@7643.4]
  wire  _T_9676; // @[Bitwise.scala 50:65:@7644.4]
  wire  _T_9677; // @[Bitwise.scala 50:65:@7645.4]
  wire  _T_9678; // @[Bitwise.scala 50:65:@7646.4]
  wire  _T_9679; // @[Bitwise.scala 50:65:@7647.4]
  wire  _T_9680; // @[Bitwise.scala 50:65:@7648.4]
  wire  _T_9681; // @[Bitwise.scala 50:65:@7649.4]
  wire  _T_9682; // @[Bitwise.scala 50:65:@7650.4]
  wire  _T_9683; // @[Bitwise.scala 50:65:@7651.4]
  wire  _T_9684; // @[Bitwise.scala 50:65:@7652.4]
  wire  _T_9685; // @[Bitwise.scala 50:65:@7653.4]
  wire  _T_9686; // @[Bitwise.scala 50:65:@7654.4]
  wire  _T_9687; // @[Bitwise.scala 50:65:@7655.4]
  wire  _T_9688; // @[Bitwise.scala 50:65:@7656.4]
  wire  _T_9689; // @[Bitwise.scala 50:65:@7657.4]
  wire  _T_9690; // @[Bitwise.scala 50:65:@7658.4]
  wire  _T_9691; // @[Bitwise.scala 50:65:@7659.4]
  wire  _T_9692; // @[Bitwise.scala 50:65:@7660.4]
  wire  _T_9693; // @[Bitwise.scala 50:65:@7661.4]
  wire  _T_9694; // @[Bitwise.scala 50:65:@7662.4]
  wire  _T_9695; // @[Bitwise.scala 50:65:@7663.4]
  wire  _T_9696; // @[Bitwise.scala 50:65:@7664.4]
  wire  _T_9697; // @[Bitwise.scala 50:65:@7665.4]
  wire  _T_9698; // @[Bitwise.scala 50:65:@7666.4]
  wire  _T_9699; // @[Bitwise.scala 50:65:@7667.4]
  wire  _T_9700; // @[Bitwise.scala 50:65:@7668.4]
  wire  _T_9701; // @[Bitwise.scala 50:65:@7669.4]
  wire  _T_9702; // @[Bitwise.scala 50:65:@7670.4]
  wire  _T_9703; // @[Bitwise.scala 50:65:@7671.4]
  wire  _T_9704; // @[Bitwise.scala 50:65:@7672.4]
  wire  _T_9705; // @[Bitwise.scala 50:65:@7673.4]
  wire  _T_9706; // @[Bitwise.scala 50:65:@7674.4]
  wire  _T_9707; // @[Bitwise.scala 50:65:@7675.4]
  wire  _T_9708; // @[Bitwise.scala 50:65:@7676.4]
  wire  _T_9709; // @[Bitwise.scala 50:65:@7677.4]
  wire  _T_9710; // @[Bitwise.scala 50:65:@7678.4]
  wire  _T_9711; // @[Bitwise.scala 50:65:@7679.4]
  wire  _T_9712; // @[Bitwise.scala 50:65:@7680.4]
  wire  _T_9713; // @[Bitwise.scala 50:65:@7681.4]
  wire  _T_9714; // @[Bitwise.scala 50:65:@7682.4]
  wire  _T_9715; // @[Bitwise.scala 50:65:@7683.4]
  wire  _T_9716; // @[Bitwise.scala 50:65:@7684.4]
  wire  _T_9717; // @[Bitwise.scala 50:65:@7685.4]
  wire  _T_9718; // @[Bitwise.scala 50:65:@7686.4]
  wire  _T_9719; // @[Bitwise.scala 50:65:@7687.4]
  wire  _T_9720; // @[Bitwise.scala 50:65:@7688.4]
  wire  _T_9721; // @[Bitwise.scala 50:65:@7689.4]
  wire  _T_9722; // @[Bitwise.scala 50:65:@7690.4]
  wire  _T_9723; // @[Bitwise.scala 50:65:@7691.4]
  wire  _T_9724; // @[Bitwise.scala 50:65:@7692.4]
  wire  _T_9725; // @[Bitwise.scala 50:65:@7693.4]
  wire  _T_9726; // @[Bitwise.scala 50:65:@7694.4]
  wire  _T_9727; // @[Bitwise.scala 50:65:@7695.4]
  wire  _T_9728; // @[Bitwise.scala 50:65:@7696.4]
  wire  _T_9729; // @[Bitwise.scala 50:65:@7697.4]
  wire  _T_9730; // @[Bitwise.scala 50:65:@7698.4]
  wire  _T_9731; // @[Bitwise.scala 50:65:@7699.4]
  wire  _T_9732; // @[Bitwise.scala 50:65:@7700.4]
  wire [1:0] _T_9733; // @[Bitwise.scala 48:55:@7701.4]
  wire [1:0] _GEN_991; // @[Bitwise.scala 48:55:@7702.4]
  wire [2:0] _T_9734; // @[Bitwise.scala 48:55:@7702.4]
  wire [1:0] _T_9735; // @[Bitwise.scala 48:55:@7703.4]
  wire [1:0] _T_9736; // @[Bitwise.scala 48:55:@7704.4]
  wire [2:0] _T_9737; // @[Bitwise.scala 48:55:@7705.4]
  wire [3:0] _T_9738; // @[Bitwise.scala 48:55:@7706.4]
  wire [1:0] _T_9739; // @[Bitwise.scala 48:55:@7707.4]
  wire [1:0] _T_9740; // @[Bitwise.scala 48:55:@7708.4]
  wire [2:0] _T_9741; // @[Bitwise.scala 48:55:@7709.4]
  wire [1:0] _T_9742; // @[Bitwise.scala 48:55:@7710.4]
  wire [1:0] _T_9743; // @[Bitwise.scala 48:55:@7711.4]
  wire [2:0] _T_9744; // @[Bitwise.scala 48:55:@7712.4]
  wire [3:0] _T_9745; // @[Bitwise.scala 48:55:@7713.4]
  wire [4:0] _T_9746; // @[Bitwise.scala 48:55:@7714.4]
  wire [1:0] _T_9747; // @[Bitwise.scala 48:55:@7715.4]
  wire [1:0] _GEN_992; // @[Bitwise.scala 48:55:@7716.4]
  wire [2:0] _T_9748; // @[Bitwise.scala 48:55:@7716.4]
  wire [1:0] _T_9749; // @[Bitwise.scala 48:55:@7717.4]
  wire [1:0] _T_9750; // @[Bitwise.scala 48:55:@7718.4]
  wire [2:0] _T_9751; // @[Bitwise.scala 48:55:@7719.4]
  wire [3:0] _T_9752; // @[Bitwise.scala 48:55:@7720.4]
  wire [1:0] _T_9753; // @[Bitwise.scala 48:55:@7721.4]
  wire [1:0] _T_9754; // @[Bitwise.scala 48:55:@7722.4]
  wire [2:0] _T_9755; // @[Bitwise.scala 48:55:@7723.4]
  wire [1:0] _T_9756; // @[Bitwise.scala 48:55:@7724.4]
  wire [1:0] _T_9757; // @[Bitwise.scala 48:55:@7725.4]
  wire [2:0] _T_9758; // @[Bitwise.scala 48:55:@7726.4]
  wire [3:0] _T_9759; // @[Bitwise.scala 48:55:@7727.4]
  wire [4:0] _T_9760; // @[Bitwise.scala 48:55:@7728.4]
  wire [5:0] _T_9761; // @[Bitwise.scala 48:55:@7729.4]
  wire [1:0] _T_9762; // @[Bitwise.scala 48:55:@7730.4]
  wire [1:0] _GEN_993; // @[Bitwise.scala 48:55:@7731.4]
  wire [2:0] _T_9763; // @[Bitwise.scala 48:55:@7731.4]
  wire [1:0] _T_9764; // @[Bitwise.scala 48:55:@7732.4]
  wire [1:0] _T_9765; // @[Bitwise.scala 48:55:@7733.4]
  wire [2:0] _T_9766; // @[Bitwise.scala 48:55:@7734.4]
  wire [3:0] _T_9767; // @[Bitwise.scala 48:55:@7735.4]
  wire [1:0] _T_9768; // @[Bitwise.scala 48:55:@7736.4]
  wire [1:0] _T_9769; // @[Bitwise.scala 48:55:@7737.4]
  wire [2:0] _T_9770; // @[Bitwise.scala 48:55:@7738.4]
  wire [1:0] _T_9771; // @[Bitwise.scala 48:55:@7739.4]
  wire [1:0] _T_9772; // @[Bitwise.scala 48:55:@7740.4]
  wire [2:0] _T_9773; // @[Bitwise.scala 48:55:@7741.4]
  wire [3:0] _T_9774; // @[Bitwise.scala 48:55:@7742.4]
  wire [4:0] _T_9775; // @[Bitwise.scala 48:55:@7743.4]
  wire [1:0] _T_9776; // @[Bitwise.scala 48:55:@7744.4]
  wire [1:0] _T_9777; // @[Bitwise.scala 48:55:@7745.4]
  wire [2:0] _T_9778; // @[Bitwise.scala 48:55:@7746.4]
  wire [1:0] _T_9779; // @[Bitwise.scala 48:55:@7747.4]
  wire [1:0] _T_9780; // @[Bitwise.scala 48:55:@7748.4]
  wire [2:0] _T_9781; // @[Bitwise.scala 48:55:@7749.4]
  wire [3:0] _T_9782; // @[Bitwise.scala 48:55:@7750.4]
  wire [1:0] _T_9783; // @[Bitwise.scala 48:55:@7751.4]
  wire [1:0] _T_9784; // @[Bitwise.scala 48:55:@7752.4]
  wire [2:0] _T_9785; // @[Bitwise.scala 48:55:@7753.4]
  wire [1:0] _T_9786; // @[Bitwise.scala 48:55:@7754.4]
  wire [1:0] _T_9787; // @[Bitwise.scala 48:55:@7755.4]
  wire [2:0] _T_9788; // @[Bitwise.scala 48:55:@7756.4]
  wire [3:0] _T_9789; // @[Bitwise.scala 48:55:@7757.4]
  wire [4:0] _T_9790; // @[Bitwise.scala 48:55:@7758.4]
  wire [5:0] _T_9791; // @[Bitwise.scala 48:55:@7759.4]
  wire [6:0] _T_9792; // @[Bitwise.scala 48:55:@7760.4]
  wire [61:0] _T_9856; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7825.4]
  wire  _T_9857; // @[Bitwise.scala 50:65:@7826.4]
  wire  _T_9858; // @[Bitwise.scala 50:65:@7827.4]
  wire  _T_9859; // @[Bitwise.scala 50:65:@7828.4]
  wire  _T_9860; // @[Bitwise.scala 50:65:@7829.4]
  wire  _T_9861; // @[Bitwise.scala 50:65:@7830.4]
  wire  _T_9862; // @[Bitwise.scala 50:65:@7831.4]
  wire  _T_9863; // @[Bitwise.scala 50:65:@7832.4]
  wire  _T_9864; // @[Bitwise.scala 50:65:@7833.4]
  wire  _T_9865; // @[Bitwise.scala 50:65:@7834.4]
  wire  _T_9866; // @[Bitwise.scala 50:65:@7835.4]
  wire  _T_9867; // @[Bitwise.scala 50:65:@7836.4]
  wire  _T_9868; // @[Bitwise.scala 50:65:@7837.4]
  wire  _T_9869; // @[Bitwise.scala 50:65:@7838.4]
  wire  _T_9870; // @[Bitwise.scala 50:65:@7839.4]
  wire  _T_9871; // @[Bitwise.scala 50:65:@7840.4]
  wire  _T_9872; // @[Bitwise.scala 50:65:@7841.4]
  wire  _T_9873; // @[Bitwise.scala 50:65:@7842.4]
  wire  _T_9874; // @[Bitwise.scala 50:65:@7843.4]
  wire  _T_9875; // @[Bitwise.scala 50:65:@7844.4]
  wire  _T_9876; // @[Bitwise.scala 50:65:@7845.4]
  wire  _T_9877; // @[Bitwise.scala 50:65:@7846.4]
  wire  _T_9878; // @[Bitwise.scala 50:65:@7847.4]
  wire  _T_9879; // @[Bitwise.scala 50:65:@7848.4]
  wire  _T_9880; // @[Bitwise.scala 50:65:@7849.4]
  wire  _T_9881; // @[Bitwise.scala 50:65:@7850.4]
  wire  _T_9882; // @[Bitwise.scala 50:65:@7851.4]
  wire  _T_9883; // @[Bitwise.scala 50:65:@7852.4]
  wire  _T_9884; // @[Bitwise.scala 50:65:@7853.4]
  wire  _T_9885; // @[Bitwise.scala 50:65:@7854.4]
  wire  _T_9886; // @[Bitwise.scala 50:65:@7855.4]
  wire  _T_9887; // @[Bitwise.scala 50:65:@7856.4]
  wire  _T_9888; // @[Bitwise.scala 50:65:@7857.4]
  wire  _T_9889; // @[Bitwise.scala 50:65:@7858.4]
  wire  _T_9890; // @[Bitwise.scala 50:65:@7859.4]
  wire  _T_9891; // @[Bitwise.scala 50:65:@7860.4]
  wire  _T_9892; // @[Bitwise.scala 50:65:@7861.4]
  wire  _T_9893; // @[Bitwise.scala 50:65:@7862.4]
  wire  _T_9894; // @[Bitwise.scala 50:65:@7863.4]
  wire  _T_9895; // @[Bitwise.scala 50:65:@7864.4]
  wire  _T_9896; // @[Bitwise.scala 50:65:@7865.4]
  wire  _T_9897; // @[Bitwise.scala 50:65:@7866.4]
  wire  _T_9898; // @[Bitwise.scala 50:65:@7867.4]
  wire  _T_9899; // @[Bitwise.scala 50:65:@7868.4]
  wire  _T_9900; // @[Bitwise.scala 50:65:@7869.4]
  wire  _T_9901; // @[Bitwise.scala 50:65:@7870.4]
  wire  _T_9902; // @[Bitwise.scala 50:65:@7871.4]
  wire  _T_9903; // @[Bitwise.scala 50:65:@7872.4]
  wire  _T_9904; // @[Bitwise.scala 50:65:@7873.4]
  wire  _T_9905; // @[Bitwise.scala 50:65:@7874.4]
  wire  _T_9906; // @[Bitwise.scala 50:65:@7875.4]
  wire  _T_9907; // @[Bitwise.scala 50:65:@7876.4]
  wire  _T_9908; // @[Bitwise.scala 50:65:@7877.4]
  wire  _T_9909; // @[Bitwise.scala 50:65:@7878.4]
  wire  _T_9910; // @[Bitwise.scala 50:65:@7879.4]
  wire  _T_9911; // @[Bitwise.scala 50:65:@7880.4]
  wire  _T_9912; // @[Bitwise.scala 50:65:@7881.4]
  wire  _T_9913; // @[Bitwise.scala 50:65:@7882.4]
  wire  _T_9914; // @[Bitwise.scala 50:65:@7883.4]
  wire  _T_9915; // @[Bitwise.scala 50:65:@7884.4]
  wire  _T_9916; // @[Bitwise.scala 50:65:@7885.4]
  wire  _T_9917; // @[Bitwise.scala 50:65:@7886.4]
  wire  _T_9918; // @[Bitwise.scala 50:65:@7887.4]
  wire [1:0] _T_9919; // @[Bitwise.scala 48:55:@7888.4]
  wire [1:0] _GEN_994; // @[Bitwise.scala 48:55:@7889.4]
  wire [2:0] _T_9920; // @[Bitwise.scala 48:55:@7889.4]
  wire [1:0] _T_9921; // @[Bitwise.scala 48:55:@7890.4]
  wire [1:0] _T_9922; // @[Bitwise.scala 48:55:@7891.4]
  wire [2:0] _T_9923; // @[Bitwise.scala 48:55:@7892.4]
  wire [3:0] _T_9924; // @[Bitwise.scala 48:55:@7893.4]
  wire [1:0] _T_9925; // @[Bitwise.scala 48:55:@7894.4]
  wire [1:0] _T_9926; // @[Bitwise.scala 48:55:@7895.4]
  wire [2:0] _T_9927; // @[Bitwise.scala 48:55:@7896.4]
  wire [1:0] _T_9928; // @[Bitwise.scala 48:55:@7897.4]
  wire [1:0] _T_9929; // @[Bitwise.scala 48:55:@7898.4]
  wire [2:0] _T_9930; // @[Bitwise.scala 48:55:@7899.4]
  wire [3:0] _T_9931; // @[Bitwise.scala 48:55:@7900.4]
  wire [4:0] _T_9932; // @[Bitwise.scala 48:55:@7901.4]
  wire [1:0] _T_9933; // @[Bitwise.scala 48:55:@7902.4]
  wire [1:0] _T_9934; // @[Bitwise.scala 48:55:@7903.4]
  wire [2:0] _T_9935; // @[Bitwise.scala 48:55:@7904.4]
  wire [1:0] _T_9936; // @[Bitwise.scala 48:55:@7905.4]
  wire [1:0] _T_9937; // @[Bitwise.scala 48:55:@7906.4]
  wire [2:0] _T_9938; // @[Bitwise.scala 48:55:@7907.4]
  wire [3:0] _T_9939; // @[Bitwise.scala 48:55:@7908.4]
  wire [1:0] _T_9940; // @[Bitwise.scala 48:55:@7909.4]
  wire [1:0] _T_9941; // @[Bitwise.scala 48:55:@7910.4]
  wire [2:0] _T_9942; // @[Bitwise.scala 48:55:@7911.4]
  wire [1:0] _T_9943; // @[Bitwise.scala 48:55:@7912.4]
  wire [1:0] _T_9944; // @[Bitwise.scala 48:55:@7913.4]
  wire [2:0] _T_9945; // @[Bitwise.scala 48:55:@7914.4]
  wire [3:0] _T_9946; // @[Bitwise.scala 48:55:@7915.4]
  wire [4:0] _T_9947; // @[Bitwise.scala 48:55:@7916.4]
  wire [5:0] _T_9948; // @[Bitwise.scala 48:55:@7917.4]
  wire [1:0] _T_9949; // @[Bitwise.scala 48:55:@7918.4]
  wire [1:0] _GEN_995; // @[Bitwise.scala 48:55:@7919.4]
  wire [2:0] _T_9950; // @[Bitwise.scala 48:55:@7919.4]
  wire [1:0] _T_9951; // @[Bitwise.scala 48:55:@7920.4]
  wire [1:0] _T_9952; // @[Bitwise.scala 48:55:@7921.4]
  wire [2:0] _T_9953; // @[Bitwise.scala 48:55:@7922.4]
  wire [3:0] _T_9954; // @[Bitwise.scala 48:55:@7923.4]
  wire [1:0] _T_9955; // @[Bitwise.scala 48:55:@7924.4]
  wire [1:0] _T_9956; // @[Bitwise.scala 48:55:@7925.4]
  wire [2:0] _T_9957; // @[Bitwise.scala 48:55:@7926.4]
  wire [1:0] _T_9958; // @[Bitwise.scala 48:55:@7927.4]
  wire [1:0] _T_9959; // @[Bitwise.scala 48:55:@7928.4]
  wire [2:0] _T_9960; // @[Bitwise.scala 48:55:@7929.4]
  wire [3:0] _T_9961; // @[Bitwise.scala 48:55:@7930.4]
  wire [4:0] _T_9962; // @[Bitwise.scala 48:55:@7931.4]
  wire [1:0] _T_9963; // @[Bitwise.scala 48:55:@7932.4]
  wire [1:0] _T_9964; // @[Bitwise.scala 48:55:@7933.4]
  wire [2:0] _T_9965; // @[Bitwise.scala 48:55:@7934.4]
  wire [1:0] _T_9966; // @[Bitwise.scala 48:55:@7935.4]
  wire [1:0] _T_9967; // @[Bitwise.scala 48:55:@7936.4]
  wire [2:0] _T_9968; // @[Bitwise.scala 48:55:@7937.4]
  wire [3:0] _T_9969; // @[Bitwise.scala 48:55:@7938.4]
  wire [1:0] _T_9970; // @[Bitwise.scala 48:55:@7939.4]
  wire [1:0] _T_9971; // @[Bitwise.scala 48:55:@7940.4]
  wire [2:0] _T_9972; // @[Bitwise.scala 48:55:@7941.4]
  wire [1:0] _T_9973; // @[Bitwise.scala 48:55:@7942.4]
  wire [1:0] _T_9974; // @[Bitwise.scala 48:55:@7943.4]
  wire [2:0] _T_9975; // @[Bitwise.scala 48:55:@7944.4]
  wire [3:0] _T_9976; // @[Bitwise.scala 48:55:@7945.4]
  wire [4:0] _T_9977; // @[Bitwise.scala 48:55:@7946.4]
  wire [5:0] _T_9978; // @[Bitwise.scala 48:55:@7947.4]
  wire [6:0] _T_9979; // @[Bitwise.scala 48:55:@7948.4]
  wire [62:0] _T_10043; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8013.4]
  wire  _T_10044; // @[Bitwise.scala 50:65:@8014.4]
  wire  _T_10045; // @[Bitwise.scala 50:65:@8015.4]
  wire  _T_10046; // @[Bitwise.scala 50:65:@8016.4]
  wire  _T_10047; // @[Bitwise.scala 50:65:@8017.4]
  wire  _T_10048; // @[Bitwise.scala 50:65:@8018.4]
  wire  _T_10049; // @[Bitwise.scala 50:65:@8019.4]
  wire  _T_10050; // @[Bitwise.scala 50:65:@8020.4]
  wire  _T_10051; // @[Bitwise.scala 50:65:@8021.4]
  wire  _T_10052; // @[Bitwise.scala 50:65:@8022.4]
  wire  _T_10053; // @[Bitwise.scala 50:65:@8023.4]
  wire  _T_10054; // @[Bitwise.scala 50:65:@8024.4]
  wire  _T_10055; // @[Bitwise.scala 50:65:@8025.4]
  wire  _T_10056; // @[Bitwise.scala 50:65:@8026.4]
  wire  _T_10057; // @[Bitwise.scala 50:65:@8027.4]
  wire  _T_10058; // @[Bitwise.scala 50:65:@8028.4]
  wire  _T_10059; // @[Bitwise.scala 50:65:@8029.4]
  wire  _T_10060; // @[Bitwise.scala 50:65:@8030.4]
  wire  _T_10061; // @[Bitwise.scala 50:65:@8031.4]
  wire  _T_10062; // @[Bitwise.scala 50:65:@8032.4]
  wire  _T_10063; // @[Bitwise.scala 50:65:@8033.4]
  wire  _T_10064; // @[Bitwise.scala 50:65:@8034.4]
  wire  _T_10065; // @[Bitwise.scala 50:65:@8035.4]
  wire  _T_10066; // @[Bitwise.scala 50:65:@8036.4]
  wire  _T_10067; // @[Bitwise.scala 50:65:@8037.4]
  wire  _T_10068; // @[Bitwise.scala 50:65:@8038.4]
  wire  _T_10069; // @[Bitwise.scala 50:65:@8039.4]
  wire  _T_10070; // @[Bitwise.scala 50:65:@8040.4]
  wire  _T_10071; // @[Bitwise.scala 50:65:@8041.4]
  wire  _T_10072; // @[Bitwise.scala 50:65:@8042.4]
  wire  _T_10073; // @[Bitwise.scala 50:65:@8043.4]
  wire  _T_10074; // @[Bitwise.scala 50:65:@8044.4]
  wire  _T_10075; // @[Bitwise.scala 50:65:@8045.4]
  wire  _T_10076; // @[Bitwise.scala 50:65:@8046.4]
  wire  _T_10077; // @[Bitwise.scala 50:65:@8047.4]
  wire  _T_10078; // @[Bitwise.scala 50:65:@8048.4]
  wire  _T_10079; // @[Bitwise.scala 50:65:@8049.4]
  wire  _T_10080; // @[Bitwise.scala 50:65:@8050.4]
  wire  _T_10081; // @[Bitwise.scala 50:65:@8051.4]
  wire  _T_10082; // @[Bitwise.scala 50:65:@8052.4]
  wire  _T_10083; // @[Bitwise.scala 50:65:@8053.4]
  wire  _T_10084; // @[Bitwise.scala 50:65:@8054.4]
  wire  _T_10085; // @[Bitwise.scala 50:65:@8055.4]
  wire  _T_10086; // @[Bitwise.scala 50:65:@8056.4]
  wire  _T_10087; // @[Bitwise.scala 50:65:@8057.4]
  wire  _T_10088; // @[Bitwise.scala 50:65:@8058.4]
  wire  _T_10089; // @[Bitwise.scala 50:65:@8059.4]
  wire  _T_10090; // @[Bitwise.scala 50:65:@8060.4]
  wire  _T_10091; // @[Bitwise.scala 50:65:@8061.4]
  wire  _T_10092; // @[Bitwise.scala 50:65:@8062.4]
  wire  _T_10093; // @[Bitwise.scala 50:65:@8063.4]
  wire  _T_10094; // @[Bitwise.scala 50:65:@8064.4]
  wire  _T_10095; // @[Bitwise.scala 50:65:@8065.4]
  wire  _T_10096; // @[Bitwise.scala 50:65:@8066.4]
  wire  _T_10097; // @[Bitwise.scala 50:65:@8067.4]
  wire  _T_10098; // @[Bitwise.scala 50:65:@8068.4]
  wire  _T_10099; // @[Bitwise.scala 50:65:@8069.4]
  wire  _T_10100; // @[Bitwise.scala 50:65:@8070.4]
  wire  _T_10101; // @[Bitwise.scala 50:65:@8071.4]
  wire  _T_10102; // @[Bitwise.scala 50:65:@8072.4]
  wire  _T_10103; // @[Bitwise.scala 50:65:@8073.4]
  wire  _T_10104; // @[Bitwise.scala 50:65:@8074.4]
  wire  _T_10105; // @[Bitwise.scala 50:65:@8075.4]
  wire  _T_10106; // @[Bitwise.scala 50:65:@8076.4]
  wire [1:0] _T_10107; // @[Bitwise.scala 48:55:@8077.4]
  wire [1:0] _GEN_996; // @[Bitwise.scala 48:55:@8078.4]
  wire [2:0] _T_10108; // @[Bitwise.scala 48:55:@8078.4]
  wire [1:0] _T_10109; // @[Bitwise.scala 48:55:@8079.4]
  wire [1:0] _T_10110; // @[Bitwise.scala 48:55:@8080.4]
  wire [2:0] _T_10111; // @[Bitwise.scala 48:55:@8081.4]
  wire [3:0] _T_10112; // @[Bitwise.scala 48:55:@8082.4]
  wire [1:0] _T_10113; // @[Bitwise.scala 48:55:@8083.4]
  wire [1:0] _T_10114; // @[Bitwise.scala 48:55:@8084.4]
  wire [2:0] _T_10115; // @[Bitwise.scala 48:55:@8085.4]
  wire [1:0] _T_10116; // @[Bitwise.scala 48:55:@8086.4]
  wire [1:0] _T_10117; // @[Bitwise.scala 48:55:@8087.4]
  wire [2:0] _T_10118; // @[Bitwise.scala 48:55:@8088.4]
  wire [3:0] _T_10119; // @[Bitwise.scala 48:55:@8089.4]
  wire [4:0] _T_10120; // @[Bitwise.scala 48:55:@8090.4]
  wire [1:0] _T_10121; // @[Bitwise.scala 48:55:@8091.4]
  wire [1:0] _T_10122; // @[Bitwise.scala 48:55:@8092.4]
  wire [2:0] _T_10123; // @[Bitwise.scala 48:55:@8093.4]
  wire [1:0] _T_10124; // @[Bitwise.scala 48:55:@8094.4]
  wire [1:0] _T_10125; // @[Bitwise.scala 48:55:@8095.4]
  wire [2:0] _T_10126; // @[Bitwise.scala 48:55:@8096.4]
  wire [3:0] _T_10127; // @[Bitwise.scala 48:55:@8097.4]
  wire [1:0] _T_10128; // @[Bitwise.scala 48:55:@8098.4]
  wire [1:0] _T_10129; // @[Bitwise.scala 48:55:@8099.4]
  wire [2:0] _T_10130; // @[Bitwise.scala 48:55:@8100.4]
  wire [1:0] _T_10131; // @[Bitwise.scala 48:55:@8101.4]
  wire [1:0] _T_10132; // @[Bitwise.scala 48:55:@8102.4]
  wire [2:0] _T_10133; // @[Bitwise.scala 48:55:@8103.4]
  wire [3:0] _T_10134; // @[Bitwise.scala 48:55:@8104.4]
  wire [4:0] _T_10135; // @[Bitwise.scala 48:55:@8105.4]
  wire [5:0] _T_10136; // @[Bitwise.scala 48:55:@8106.4]
  wire [1:0] _T_10137; // @[Bitwise.scala 48:55:@8107.4]
  wire [1:0] _T_10138; // @[Bitwise.scala 48:55:@8108.4]
  wire [2:0] _T_10139; // @[Bitwise.scala 48:55:@8109.4]
  wire [1:0] _T_10140; // @[Bitwise.scala 48:55:@8110.4]
  wire [1:0] _T_10141; // @[Bitwise.scala 48:55:@8111.4]
  wire [2:0] _T_10142; // @[Bitwise.scala 48:55:@8112.4]
  wire [3:0] _T_10143; // @[Bitwise.scala 48:55:@8113.4]
  wire [1:0] _T_10144; // @[Bitwise.scala 48:55:@8114.4]
  wire [1:0] _T_10145; // @[Bitwise.scala 48:55:@8115.4]
  wire [2:0] _T_10146; // @[Bitwise.scala 48:55:@8116.4]
  wire [1:0] _T_10147; // @[Bitwise.scala 48:55:@8117.4]
  wire [1:0] _T_10148; // @[Bitwise.scala 48:55:@8118.4]
  wire [2:0] _T_10149; // @[Bitwise.scala 48:55:@8119.4]
  wire [3:0] _T_10150; // @[Bitwise.scala 48:55:@8120.4]
  wire [4:0] _T_10151; // @[Bitwise.scala 48:55:@8121.4]
  wire [1:0] _T_10152; // @[Bitwise.scala 48:55:@8122.4]
  wire [1:0] _T_10153; // @[Bitwise.scala 48:55:@8123.4]
  wire [2:0] _T_10154; // @[Bitwise.scala 48:55:@8124.4]
  wire [1:0] _T_10155; // @[Bitwise.scala 48:55:@8125.4]
  wire [1:0] _T_10156; // @[Bitwise.scala 48:55:@8126.4]
  wire [2:0] _T_10157; // @[Bitwise.scala 48:55:@8127.4]
  wire [3:0] _T_10158; // @[Bitwise.scala 48:55:@8128.4]
  wire [1:0] _T_10159; // @[Bitwise.scala 48:55:@8129.4]
  wire [1:0] _T_10160; // @[Bitwise.scala 48:55:@8130.4]
  wire [2:0] _T_10161; // @[Bitwise.scala 48:55:@8131.4]
  wire [1:0] _T_10162; // @[Bitwise.scala 48:55:@8132.4]
  wire [1:0] _T_10163; // @[Bitwise.scala 48:55:@8133.4]
  wire [2:0] _T_10164; // @[Bitwise.scala 48:55:@8134.4]
  wire [3:0] _T_10165; // @[Bitwise.scala 48:55:@8135.4]
  wire [4:0] _T_10166; // @[Bitwise.scala 48:55:@8136.4]
  wire [5:0] _T_10167; // @[Bitwise.scala 48:55:@8137.4]
  wire [6:0] _T_10168; // @[Bitwise.scala 48:55:@8138.4]
  wire  _T_10234; // @[Bitwise.scala 50:65:@8205.4]
  wire  _T_10235; // @[Bitwise.scala 50:65:@8206.4]
  wire  _T_10236; // @[Bitwise.scala 50:65:@8207.4]
  wire  _T_10237; // @[Bitwise.scala 50:65:@8208.4]
  wire  _T_10238; // @[Bitwise.scala 50:65:@8209.4]
  wire  _T_10239; // @[Bitwise.scala 50:65:@8210.4]
  wire  _T_10240; // @[Bitwise.scala 50:65:@8211.4]
  wire  _T_10241; // @[Bitwise.scala 50:65:@8212.4]
  wire  _T_10242; // @[Bitwise.scala 50:65:@8213.4]
  wire  _T_10243; // @[Bitwise.scala 50:65:@8214.4]
  wire  _T_10244; // @[Bitwise.scala 50:65:@8215.4]
  wire  _T_10245; // @[Bitwise.scala 50:65:@8216.4]
  wire  _T_10246; // @[Bitwise.scala 50:65:@8217.4]
  wire  _T_10247; // @[Bitwise.scala 50:65:@8218.4]
  wire  _T_10248; // @[Bitwise.scala 50:65:@8219.4]
  wire  _T_10249; // @[Bitwise.scala 50:65:@8220.4]
  wire  _T_10250; // @[Bitwise.scala 50:65:@8221.4]
  wire  _T_10251; // @[Bitwise.scala 50:65:@8222.4]
  wire  _T_10252; // @[Bitwise.scala 50:65:@8223.4]
  wire  _T_10253; // @[Bitwise.scala 50:65:@8224.4]
  wire  _T_10254; // @[Bitwise.scala 50:65:@8225.4]
  wire  _T_10255; // @[Bitwise.scala 50:65:@8226.4]
  wire  _T_10256; // @[Bitwise.scala 50:65:@8227.4]
  wire  _T_10257; // @[Bitwise.scala 50:65:@8228.4]
  wire  _T_10258; // @[Bitwise.scala 50:65:@8229.4]
  wire  _T_10259; // @[Bitwise.scala 50:65:@8230.4]
  wire  _T_10260; // @[Bitwise.scala 50:65:@8231.4]
  wire  _T_10261; // @[Bitwise.scala 50:65:@8232.4]
  wire  _T_10262; // @[Bitwise.scala 50:65:@8233.4]
  wire  _T_10263; // @[Bitwise.scala 50:65:@8234.4]
  wire  _T_10264; // @[Bitwise.scala 50:65:@8235.4]
  wire  _T_10265; // @[Bitwise.scala 50:65:@8236.4]
  wire  _T_10266; // @[Bitwise.scala 50:65:@8237.4]
  wire  _T_10267; // @[Bitwise.scala 50:65:@8238.4]
  wire  _T_10268; // @[Bitwise.scala 50:65:@8239.4]
  wire  _T_10269; // @[Bitwise.scala 50:65:@8240.4]
  wire  _T_10270; // @[Bitwise.scala 50:65:@8241.4]
  wire  _T_10271; // @[Bitwise.scala 50:65:@8242.4]
  wire  _T_10272; // @[Bitwise.scala 50:65:@8243.4]
  wire  _T_10273; // @[Bitwise.scala 50:65:@8244.4]
  wire  _T_10274; // @[Bitwise.scala 50:65:@8245.4]
  wire  _T_10275; // @[Bitwise.scala 50:65:@8246.4]
  wire  _T_10276; // @[Bitwise.scala 50:65:@8247.4]
  wire  _T_10277; // @[Bitwise.scala 50:65:@8248.4]
  wire  _T_10278; // @[Bitwise.scala 50:65:@8249.4]
  wire  _T_10279; // @[Bitwise.scala 50:65:@8250.4]
  wire  _T_10280; // @[Bitwise.scala 50:65:@8251.4]
  wire  _T_10281; // @[Bitwise.scala 50:65:@8252.4]
  wire  _T_10282; // @[Bitwise.scala 50:65:@8253.4]
  wire  _T_10283; // @[Bitwise.scala 50:65:@8254.4]
  wire  _T_10284; // @[Bitwise.scala 50:65:@8255.4]
  wire  _T_10285; // @[Bitwise.scala 50:65:@8256.4]
  wire  _T_10286; // @[Bitwise.scala 50:65:@8257.4]
  wire  _T_10287; // @[Bitwise.scala 50:65:@8258.4]
  wire  _T_10288; // @[Bitwise.scala 50:65:@8259.4]
  wire  _T_10289; // @[Bitwise.scala 50:65:@8260.4]
  wire  _T_10290; // @[Bitwise.scala 50:65:@8261.4]
  wire  _T_10291; // @[Bitwise.scala 50:65:@8262.4]
  wire  _T_10292; // @[Bitwise.scala 50:65:@8263.4]
  wire  _T_10293; // @[Bitwise.scala 50:65:@8264.4]
  wire  _T_10294; // @[Bitwise.scala 50:65:@8265.4]
  wire  _T_10295; // @[Bitwise.scala 50:65:@8266.4]
  wire  _T_10296; // @[Bitwise.scala 50:65:@8267.4]
  wire [1:0] _T_10297; // @[Bitwise.scala 48:55:@8268.4]
  wire [1:0] _T_10298; // @[Bitwise.scala 48:55:@8269.4]
  wire [2:0] _T_10299; // @[Bitwise.scala 48:55:@8270.4]
  wire [1:0] _T_10300; // @[Bitwise.scala 48:55:@8271.4]
  wire [1:0] _T_10301; // @[Bitwise.scala 48:55:@8272.4]
  wire [2:0] _T_10302; // @[Bitwise.scala 48:55:@8273.4]
  wire [3:0] _T_10303; // @[Bitwise.scala 48:55:@8274.4]
  wire [1:0] _T_10304; // @[Bitwise.scala 48:55:@8275.4]
  wire [1:0] _T_10305; // @[Bitwise.scala 48:55:@8276.4]
  wire [2:0] _T_10306; // @[Bitwise.scala 48:55:@8277.4]
  wire [1:0] _T_10307; // @[Bitwise.scala 48:55:@8278.4]
  wire [1:0] _T_10308; // @[Bitwise.scala 48:55:@8279.4]
  wire [2:0] _T_10309; // @[Bitwise.scala 48:55:@8280.4]
  wire [3:0] _T_10310; // @[Bitwise.scala 48:55:@8281.4]
  wire [4:0] _T_10311; // @[Bitwise.scala 48:55:@8282.4]
  wire [1:0] _T_10312; // @[Bitwise.scala 48:55:@8283.4]
  wire [1:0] _T_10313; // @[Bitwise.scala 48:55:@8284.4]
  wire [2:0] _T_10314; // @[Bitwise.scala 48:55:@8285.4]
  wire [1:0] _T_10315; // @[Bitwise.scala 48:55:@8286.4]
  wire [1:0] _T_10316; // @[Bitwise.scala 48:55:@8287.4]
  wire [2:0] _T_10317; // @[Bitwise.scala 48:55:@8288.4]
  wire [3:0] _T_10318; // @[Bitwise.scala 48:55:@8289.4]
  wire [1:0] _T_10319; // @[Bitwise.scala 48:55:@8290.4]
  wire [1:0] _T_10320; // @[Bitwise.scala 48:55:@8291.4]
  wire [2:0] _T_10321; // @[Bitwise.scala 48:55:@8292.4]
  wire [1:0] _T_10322; // @[Bitwise.scala 48:55:@8293.4]
  wire [1:0] _T_10323; // @[Bitwise.scala 48:55:@8294.4]
  wire [2:0] _T_10324; // @[Bitwise.scala 48:55:@8295.4]
  wire [3:0] _T_10325; // @[Bitwise.scala 48:55:@8296.4]
  wire [4:0] _T_10326; // @[Bitwise.scala 48:55:@8297.4]
  wire [5:0] _T_10327; // @[Bitwise.scala 48:55:@8298.4]
  wire [1:0] _T_10328; // @[Bitwise.scala 48:55:@8299.4]
  wire [1:0] _T_10329; // @[Bitwise.scala 48:55:@8300.4]
  wire [2:0] _T_10330; // @[Bitwise.scala 48:55:@8301.4]
  wire [1:0] _T_10331; // @[Bitwise.scala 48:55:@8302.4]
  wire [1:0] _T_10332; // @[Bitwise.scala 48:55:@8303.4]
  wire [2:0] _T_10333; // @[Bitwise.scala 48:55:@8304.4]
  wire [3:0] _T_10334; // @[Bitwise.scala 48:55:@8305.4]
  wire [1:0] _T_10335; // @[Bitwise.scala 48:55:@8306.4]
  wire [1:0] _T_10336; // @[Bitwise.scala 48:55:@8307.4]
  wire [2:0] _T_10337; // @[Bitwise.scala 48:55:@8308.4]
  wire [1:0] _T_10338; // @[Bitwise.scala 48:55:@8309.4]
  wire [1:0] _T_10339; // @[Bitwise.scala 48:55:@8310.4]
  wire [2:0] _T_10340; // @[Bitwise.scala 48:55:@8311.4]
  wire [3:0] _T_10341; // @[Bitwise.scala 48:55:@8312.4]
  wire [4:0] _T_10342; // @[Bitwise.scala 48:55:@8313.4]
  wire [1:0] _T_10343; // @[Bitwise.scala 48:55:@8314.4]
  wire [1:0] _T_10344; // @[Bitwise.scala 48:55:@8315.4]
  wire [2:0] _T_10345; // @[Bitwise.scala 48:55:@8316.4]
  wire [1:0] _T_10346; // @[Bitwise.scala 48:55:@8317.4]
  wire [1:0] _T_10347; // @[Bitwise.scala 48:55:@8318.4]
  wire [2:0] _T_10348; // @[Bitwise.scala 48:55:@8319.4]
  wire [3:0] _T_10349; // @[Bitwise.scala 48:55:@8320.4]
  wire [1:0] _T_10350; // @[Bitwise.scala 48:55:@8321.4]
  wire [1:0] _T_10351; // @[Bitwise.scala 48:55:@8322.4]
  wire [2:0] _T_10352; // @[Bitwise.scala 48:55:@8323.4]
  wire [1:0] _T_10353; // @[Bitwise.scala 48:55:@8324.4]
  wire [1:0] _T_10354; // @[Bitwise.scala 48:55:@8325.4]
  wire [2:0] _T_10355; // @[Bitwise.scala 48:55:@8326.4]
  wire [3:0] _T_10356; // @[Bitwise.scala 48:55:@8327.4]
  wire [4:0] _T_10357; // @[Bitwise.scala 48:55:@8328.4]
  wire [5:0] _T_10358; // @[Bitwise.scala 48:55:@8329.4]
  wire [6:0] _T_10359; // @[Bitwise.scala 48:55:@8330.4]
  reg  _T_10362; // @[NV_NVDLA_CSC_WL_dec.scala 64:27:@8332.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_10366_0; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_10366_1; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_10366_2; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_10366_3; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_10366_4; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_10366_5; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_10366_6; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_10366_7; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_10366_8; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_10366_9; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_10366_10; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_10366_11; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_10366_12; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_10366_13; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_10366_14; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_10366_15; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_10366_16; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_10366_17; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_10366_18; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_10366_19; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_10366_20; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_10366_21; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_10366_22; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_10366_23; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_10366_24; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_10366_25; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_10366_26; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_10366_27; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_10366_28; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_10366_29; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_10366_30; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_10366_31; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_10366_32; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_10366_33; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_10366_34; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_10366_35; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_10366_36; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_10366_37; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_10366_38; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_10366_39; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_10366_40; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_10366_41; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_10366_42; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_10366_43; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_10366_44; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_10366_45; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_10366_46; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_10366_47; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_10366_48; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_10366_49; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_10366_50; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_10366_51; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_10366_52; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_10366_53; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_10366_54; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_10366_55; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_10366_56; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_10366_57; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_10366_58; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_10366_59; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_10366_60; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_10366_61; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_10366_62; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_10366_63; // @[NV_NVDLA_CSC_WL_dec.scala 65:22:@8333.4]
  reg [31:0] _RAND_64;
  reg  _T_10436_0; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_65;
  reg  _T_10436_1; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_66;
  reg  _T_10436_2; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_67;
  reg  _T_10436_3; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_68;
  reg  _T_10436_4; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_69;
  reg  _T_10436_5; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_70;
  reg  _T_10436_6; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_71;
  reg  _T_10436_7; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_72;
  reg  _T_10436_8; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_73;
  reg  _T_10436_9; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_74;
  reg  _T_10436_10; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_75;
  reg  _T_10436_11; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_76;
  reg  _T_10436_12; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_77;
  reg  _T_10436_13; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_78;
  reg  _T_10436_14; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_79;
  reg  _T_10436_15; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_80;
  reg  _T_10436_16; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_81;
  reg  _T_10436_17; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_82;
  reg  _T_10436_18; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_83;
  reg  _T_10436_19; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_84;
  reg  _T_10436_20; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_85;
  reg  _T_10436_21; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_86;
  reg  _T_10436_22; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_87;
  reg  _T_10436_23; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_88;
  reg  _T_10436_24; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_89;
  reg  _T_10436_25; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_90;
  reg  _T_10436_26; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_91;
  reg  _T_10436_27; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_92;
  reg  _T_10436_28; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_93;
  reg  _T_10436_29; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_94;
  reg  _T_10436_30; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_95;
  reg  _T_10436_31; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_96;
  reg  _T_10436_32; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_97;
  reg  _T_10436_33; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_98;
  reg  _T_10436_34; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_99;
  reg  _T_10436_35; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_100;
  reg  _T_10436_36; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_101;
  reg  _T_10436_37; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_102;
  reg  _T_10436_38; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_103;
  reg  _T_10436_39; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_104;
  reg  _T_10436_40; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_105;
  reg  _T_10436_41; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_106;
  reg  _T_10436_42; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_107;
  reg  _T_10436_43; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_108;
  reg  _T_10436_44; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_109;
  reg  _T_10436_45; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_110;
  reg  _T_10436_46; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_111;
  reg  _T_10436_47; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_112;
  reg  _T_10436_48; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_113;
  reg  _T_10436_49; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_114;
  reg  _T_10436_50; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_115;
  reg  _T_10436_51; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_116;
  reg  _T_10436_52; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_117;
  reg  _T_10436_53; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_118;
  reg  _T_10436_54; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_119;
  reg  _T_10436_55; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_120;
  reg  _T_10436_56; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_121;
  reg  _T_10436_57; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_122;
  reg  _T_10436_58; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_123;
  reg  _T_10436_59; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_124;
  reg  _T_10436_60; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_125;
  reg  _T_10436_61; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_126;
  reg  _T_10436_62; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_127;
  reg  _T_10436_63; // @[NV_NVDLA_CSC_WL_dec.scala 66:22:@8334.4]
  reg [31:0] _RAND_128;
  reg  _T_10641_0; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_129;
  reg  _T_10641_1; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_130;
  reg  _T_10641_2; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_131;
  reg  _T_10641_3; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_132;
  reg  _T_10641_4; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_133;
  reg  _T_10641_5; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_134;
  reg  _T_10641_6; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_135;
  reg  _T_10641_7; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_136;
  reg  _T_10641_8; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_137;
  reg  _T_10641_9; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_138;
  reg  _T_10641_10; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_139;
  reg  _T_10641_11; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_140;
  reg  _T_10641_12; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_141;
  reg  _T_10641_13; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_142;
  reg  _T_10641_14; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_143;
  reg  _T_10641_15; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_144;
  reg  _T_10641_16; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_145;
  reg  _T_10641_17; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_146;
  reg  _T_10641_18; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_147;
  reg  _T_10641_19; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_148;
  reg  _T_10641_20; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_149;
  reg  _T_10641_21; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_150;
  reg  _T_10641_22; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_151;
  reg  _T_10641_23; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_152;
  reg  _T_10641_24; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_153;
  reg  _T_10641_25; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_154;
  reg  _T_10641_26; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_155;
  reg  _T_10641_27; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_156;
  reg  _T_10641_28; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_157;
  reg  _T_10641_29; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_158;
  reg  _T_10641_30; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_159;
  reg  _T_10641_31; // @[NV_NVDLA_CSC_WL_dec.scala 67:25:@8368.4]
  reg [31:0] _RAND_160;
  reg [6:0] _T_11317_63; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_161;
  reg [5:0] _T_11317_62; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_162;
  reg [5:0] _T_11317_61; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_163;
  reg [5:0] _T_11317_60; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_164;
  reg [5:0] _T_11317_59; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_165;
  reg [5:0] _T_11317_58; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_166;
  reg [5:0] _T_11317_57; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_167;
  reg [5:0] _T_11317_56; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_168;
  reg [5:0] _T_11317_55; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_169;
  reg [5:0] _T_11317_54; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_170;
  reg [5:0] _T_11317_53; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_171;
  reg [5:0] _T_11317_52; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_172;
  reg [5:0] _T_11317_51; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_173;
  reg [5:0] _T_11317_50; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_174;
  reg [5:0] _T_11317_49; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_175;
  reg [5:0] _T_11317_48; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_176;
  reg [5:0] _T_11317_47; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_177;
  reg [5:0] _T_11317_46; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_178;
  reg [5:0] _T_11317_45; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_179;
  reg [5:0] _T_11317_44; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_180;
  reg [5:0] _T_11317_43; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_181;
  reg [5:0] _T_11317_42; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_182;
  reg [5:0] _T_11317_41; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_183;
  reg [5:0] _T_11317_40; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_184;
  reg [5:0] _T_11317_39; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_185;
  reg [5:0] _T_11317_38; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_186;
  reg [5:0] _T_11317_37; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_187;
  reg [5:0] _T_11317_36; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_188;
  reg [5:0] _T_11317_35; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_189;
  reg [5:0] _T_11317_34; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_190;
  reg [5:0] _T_11317_33; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_191;
  reg [5:0] _T_11317_32; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_192;
  reg [5:0] _T_11317_31; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_193;
  reg [4:0] _T_11317_30; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_194;
  reg [4:0] _T_11317_29; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_195;
  reg [4:0] _T_11317_28; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_196;
  reg [4:0] _T_11317_27; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_197;
  reg [4:0] _T_11317_26; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_198;
  reg [4:0] _T_11317_25; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_199;
  reg [4:0] _T_11317_24; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_200;
  reg [4:0] _T_11317_23; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_201;
  reg [4:0] _T_11317_22; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_202;
  reg [4:0] _T_11317_21; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_203;
  reg [4:0] _T_11317_20; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_204;
  reg [4:0] _T_11317_19; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_205;
  reg [4:0] _T_11317_18; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_206;
  reg [4:0] _T_11317_17; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_207;
  reg [4:0] _T_11317_16; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_208;
  reg [4:0] _T_11317_15; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_209;
  reg [3:0] _T_11317_14; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_210;
  reg [3:0] _T_11317_13; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_211;
  reg [3:0] _T_11317_12; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_212;
  reg [3:0] _T_11317_11; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_213;
  reg [3:0] _T_11317_10; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_214;
  reg [3:0] _T_11317_9; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_215;
  reg [3:0] _T_11317_8; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_216;
  reg [3:0] _T_11317_7; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_217;
  reg [2:0] _T_11317_6; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_218;
  reg [2:0] _T_11317_5; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_219;
  reg [2:0] _T_11317_4; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_220;
  reg [2:0] _T_11317_3; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_221;
  reg [1:0] _T_11317_2; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_222;
  reg [1:0] _T_11317_1; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_223;
  reg  _T_11317_0; // @[NV_NVDLA_CSC_WL_dec.scala 68:29:@8497.4]
  reg [31:0] _RAND_224;
  wire  _GEN_128; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_129; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_130; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_131; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_132; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_133; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_134; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_135; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_136; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_137; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_138; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_139; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_140; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_141; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_142; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_143; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_144; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_145; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_146; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_147; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_148; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_149; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_150; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_151; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_152; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_153; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_154; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_155; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  wire  _T_11318; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8661.4]
  wire  _T_11319; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8662.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8663.4]
  wire [1:0] _GEN_161; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8668.4]
  wire [1:0] _T_2167_2; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@279.4]
  wire [1:0] _GEN_162; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8673.4]
  wire [2:0] _GEN_163; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8678.4]
  wire [2:0] _T_2167_4; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@425.4]
  wire [2:0] _GEN_164; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8683.4]
  wire [2:0] _T_2167_5; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@501.4]
  wire [2:0] _GEN_165; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8688.4]
  wire [2:0] _T_2167_6; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@579.4]
  wire [2:0] _GEN_166; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8693.4]
  wire [3:0] _GEN_167; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8698.4]
  wire  _T_11334; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8701.4]
  wire  _T_11335; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8702.4]
  wire [3:0] _T_2167_8; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@741.4]
  wire [3:0] _GEN_168; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8703.4]
  wire [3:0] _T_2167_9; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@825.4]
  wire [3:0] _GEN_169; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8708.4]
  wire [3:0] _T_2167_10; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@911.4]
  wire [3:0] _GEN_170; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8713.4]
  wire [3:0] _T_2167_11; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@999.4]
  wire [3:0] _GEN_171; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8718.4]
  wire [3:0] _T_2167_12; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1089.4]
  wire [3:0] _GEN_172; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8723.4]
  wire [3:0] _T_2167_13; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1181.4]
  wire [3:0] _GEN_173; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8728.4]
  wire [3:0] _T_2167_14; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1275.4]
  wire [3:0] _GEN_174; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8733.4]
  wire [4:0] _GEN_175; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8738.4]
  wire  _T_11350; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8741.4]
  wire  _T_11351; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8742.4]
  wire [4:0] _T_2167_16; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1469.4]
  wire [4:0] _GEN_176; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8743.4]
  wire [4:0] _T_2167_17; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1569.4]
  wire [4:0] _GEN_177; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8748.4]
  wire [4:0] _T_2167_18; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1671.4]
  wire [4:0] _GEN_178; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8753.4]
  wire [4:0] _T_2167_19; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1775.4]
  wire [4:0] _GEN_179; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8758.4]
  wire [4:0] _T_2167_20; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1881.4]
  wire [4:0] _GEN_180; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8763.4]
  wire [4:0] _T_2167_21; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1989.4]
  wire [4:0] _GEN_181; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8768.4]
  wire [4:0] _T_2167_22; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2099.4]
  wire [4:0] _GEN_182; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8773.4]
  wire [4:0] _T_2167_23; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2211.4]
  wire [4:0] _GEN_183; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8778.4]
  wire  _T_11366; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8781.4]
  wire  _T_11367; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8782.4]
  wire [4:0] _T_2167_24; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2325.4]
  wire [4:0] _GEN_184; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8783.4]
  wire [4:0] _T_2167_25; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2441.4]
  wire [4:0] _GEN_185; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8788.4]
  wire [4:0] _T_2167_26; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2559.4]
  wire [4:0] _GEN_186; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8793.4]
  wire [4:0] _T_2167_27; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2679.4]
  wire [4:0] _GEN_187; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8798.4]
  wire [4:0] _T_2167_28; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2801.4]
  wire [4:0] _GEN_188; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8803.4]
  wire [4:0] _T_2167_29; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2925.4]
  wire [4:0] _GEN_189; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8808.4]
  wire [4:0] _T_2167_30; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3051.4]
  wire [4:0] _GEN_190; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8813.4]
  wire [5:0] _GEN_191; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8818.4]
  wire  _T_11382; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8821.4]
  wire  _T_11383; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8822.4]
  wire [5:0] _T_2167_32; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3309.4]
  wire [5:0] _GEN_192; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8823.4]
  wire [5:0] _T_2167_33; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3441.4]
  wire [5:0] _GEN_193; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8828.4]
  wire [5:0] _T_2167_34; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3575.4]
  wire [5:0] _GEN_194; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8833.4]
  wire [5:0] _T_2167_35; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3711.4]
  wire [5:0] _GEN_195; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8838.4]
  wire [5:0] _T_2167_36; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3849.4]
  wire [5:0] _GEN_196; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8843.4]
  wire [5:0] _T_2167_37; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3989.4]
  wire [5:0] _GEN_197; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8848.4]
  wire [5:0] _T_2167_38; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4131.4]
  wire [5:0] _GEN_198; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8853.4]
  wire [5:0] _T_2167_39; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4275.4]
  wire [5:0] _GEN_199; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8858.4]
  wire  _T_11398; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8861.4]
  wire  _T_11399; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8862.4]
  wire [5:0] _T_2167_40; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4421.4]
  wire [5:0] _GEN_200; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8863.4]
  wire [5:0] _T_2167_41; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4569.4]
  wire [5:0] _GEN_201; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8868.4]
  wire [5:0] _T_2167_42; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4719.4]
  wire [5:0] _GEN_202; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8873.4]
  wire [5:0] _T_2167_43; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4871.4]
  wire [5:0] _GEN_203; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8878.4]
  wire [5:0] _T_2167_44; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5025.4]
  wire [5:0] _GEN_204; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8883.4]
  wire [5:0] _T_2167_45; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5181.4]
  wire [5:0] _GEN_205; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8888.4]
  wire [5:0] _T_2167_46; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5339.4]
  wire [5:0] _GEN_206; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8893.4]
  wire [5:0] _T_2167_47; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5499.4]
  wire [5:0] _GEN_207; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8898.4]
  wire  _T_11414; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8901.4]
  wire  _T_11415; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8902.4]
  wire [5:0] _T_2167_48; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5661.4]
  wire [5:0] _GEN_208; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8903.4]
  wire [5:0] _T_2167_49; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5825.4]
  wire [5:0] _GEN_209; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8908.4]
  wire [5:0] _T_2167_50; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5991.4]
  wire [5:0] _GEN_210; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8913.4]
  wire [5:0] _T_2167_51; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6159.4]
  wire [5:0] _GEN_211; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8918.4]
  wire [5:0] _T_2167_52; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6329.4]
  wire [5:0] _GEN_212; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8923.4]
  wire [5:0] _T_2167_53; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6501.4]
  wire [5:0] _GEN_213; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8928.4]
  wire [5:0] _T_2167_54; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6675.4]
  wire [5:0] _GEN_214; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8933.4]
  wire [5:0] _T_2167_55; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6851.4]
  wire [5:0] _GEN_215; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8938.4]
  wire  _T_11430; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8941.4]
  wire  _T_11431; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8942.4]
  wire [5:0] _T_2167_56; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7029.4]
  wire [5:0] _GEN_216; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8943.4]
  wire [5:0] _T_2167_57; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7209.4]
  wire [5:0] _GEN_217; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8948.4]
  wire [5:0] _T_2167_58; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7391.4]
  wire [5:0] _GEN_218; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8953.4]
  wire [5:0] _T_2167_59; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7575.4]
  wire [5:0] _GEN_219; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8958.4]
  wire [5:0] _T_2167_60; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7761.4]
  wire [5:0] _GEN_220; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8963.4]
  wire [5:0] _T_2167_61; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7949.4]
  wire [5:0] _GEN_221; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8968.4]
  wire [5:0] _T_2167_62; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8139.4]
  wire [5:0] _GEN_222; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8973.4]
  wire [6:0] _GEN_223; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8978.4]
  wire [7:0] _T_11519; // @[Mux.scala 46:16:@8983.4]
  wire  _T_11523; // @[Mux.scala 46:19:@8985.4]
  wire [7:0] _T_11524; // @[Mux.scala 46:16:@8986.4]
  wire  _T_11525; // @[Mux.scala 46:19:@8987.4]
  wire [7:0] _T_11526; // @[Mux.scala 46:16:@8988.4]
  wire  _T_11531; // @[Mux.scala 46:19:@8990.4]
  wire [7:0] _T_11532; // @[Mux.scala 46:16:@8991.4]
  wire  _T_11533; // @[Mux.scala 46:19:@8992.4]
  wire [7:0] _T_11534; // @[Mux.scala 46:16:@8993.4]
  wire  _T_11535; // @[Mux.scala 46:19:@8994.4]
  wire [7:0] _T_11536; // @[Mux.scala 46:16:@8995.4]
  wire  _T_11542; // @[Mux.scala 46:19:@8997.4]
  wire [7:0] _T_11543; // @[Mux.scala 46:16:@8998.4]
  wire  _T_11544; // @[Mux.scala 46:19:@8999.4]
  wire [7:0] _T_11545; // @[Mux.scala 46:16:@9000.4]
  wire  _T_11546; // @[Mux.scala 46:19:@9001.4]
  wire [7:0] _T_11547; // @[Mux.scala 46:16:@9002.4]
  wire  _T_11548; // @[Mux.scala 46:19:@9003.4]
  wire [7:0] _T_11549; // @[Mux.scala 46:16:@9004.4]
  wire  _T_11556; // @[Mux.scala 46:19:@9006.4]
  wire [7:0] _T_11557; // @[Mux.scala 46:16:@9007.4]
  wire  _T_11558; // @[Mux.scala 46:19:@9008.4]
  wire [7:0] _T_11559; // @[Mux.scala 46:16:@9009.4]
  wire  _T_11560; // @[Mux.scala 46:19:@9010.4]
  wire [7:0] _T_11561; // @[Mux.scala 46:16:@9011.4]
  wire  _T_11562; // @[Mux.scala 46:19:@9012.4]
  wire [7:0] _T_11563; // @[Mux.scala 46:16:@9013.4]
  wire  _T_11564; // @[Mux.scala 46:19:@9014.4]
  wire [7:0] _T_11565; // @[Mux.scala 46:16:@9015.4]
  wire  _T_11573; // @[Mux.scala 46:19:@9017.4]
  wire [7:0] _T_11574; // @[Mux.scala 46:16:@9018.4]
  wire  _T_11575; // @[Mux.scala 46:19:@9019.4]
  wire [7:0] _T_11576; // @[Mux.scala 46:16:@9020.4]
  wire  _T_11577; // @[Mux.scala 46:19:@9021.4]
  wire [7:0] _T_11578; // @[Mux.scala 46:16:@9022.4]
  wire  _T_11579; // @[Mux.scala 46:19:@9023.4]
  wire [7:0] _T_11580; // @[Mux.scala 46:16:@9024.4]
  wire  _T_11581; // @[Mux.scala 46:19:@9025.4]
  wire [7:0] _T_11582; // @[Mux.scala 46:16:@9026.4]
  wire  _T_11583; // @[Mux.scala 46:19:@9027.4]
  wire [7:0] _T_11584; // @[Mux.scala 46:16:@9028.4]
  wire  _T_11593; // @[Mux.scala 46:19:@9030.4]
  wire [7:0] _T_11594; // @[Mux.scala 46:16:@9031.4]
  wire  _T_11595; // @[Mux.scala 46:19:@9032.4]
  wire [7:0] _T_11596; // @[Mux.scala 46:16:@9033.4]
  wire  _T_11597; // @[Mux.scala 46:19:@9034.4]
  wire [7:0] _T_11598; // @[Mux.scala 46:16:@9035.4]
  wire  _T_11599; // @[Mux.scala 46:19:@9036.4]
  wire [7:0] _T_11600; // @[Mux.scala 46:16:@9037.4]
  wire  _T_11601; // @[Mux.scala 46:19:@9038.4]
  wire [7:0] _T_11602; // @[Mux.scala 46:16:@9039.4]
  wire  _T_11603; // @[Mux.scala 46:19:@9040.4]
  wire [7:0] _T_11604; // @[Mux.scala 46:16:@9041.4]
  wire  _T_11605; // @[Mux.scala 46:19:@9042.4]
  wire [7:0] _T_11606; // @[Mux.scala 46:16:@9043.4]
  wire  _T_11616; // @[Mux.scala 46:19:@9045.4]
  wire [7:0] _T_11617; // @[Mux.scala 46:16:@9046.4]
  wire  _T_11618; // @[Mux.scala 46:19:@9047.4]
  wire [7:0] _T_11619; // @[Mux.scala 46:16:@9048.4]
  wire  _T_11620; // @[Mux.scala 46:19:@9049.4]
  wire [7:0] _T_11621; // @[Mux.scala 46:16:@9050.4]
  wire  _T_11622; // @[Mux.scala 46:19:@9051.4]
  wire [7:0] _T_11623; // @[Mux.scala 46:16:@9052.4]
  wire  _T_11624; // @[Mux.scala 46:19:@9053.4]
  wire [7:0] _T_11625; // @[Mux.scala 46:16:@9054.4]
  wire  _T_11626; // @[Mux.scala 46:19:@9055.4]
  wire [7:0] _T_11627; // @[Mux.scala 46:16:@9056.4]
  wire  _T_11628; // @[Mux.scala 46:19:@9057.4]
  wire [7:0] _T_11629; // @[Mux.scala 46:16:@9058.4]
  wire  _T_11630; // @[Mux.scala 46:19:@9059.4]
  wire [7:0] _T_11631; // @[Mux.scala 46:16:@9060.4]
  wire  _T_11642; // @[Mux.scala 46:19:@9062.4]
  wire [7:0] _T_11643; // @[Mux.scala 46:16:@9063.4]
  wire  _T_11644; // @[Mux.scala 46:19:@9064.4]
  wire [7:0] _T_11645; // @[Mux.scala 46:16:@9065.4]
  wire  _T_11646; // @[Mux.scala 46:19:@9066.4]
  wire [7:0] _T_11647; // @[Mux.scala 46:16:@9067.4]
  wire  _T_11648; // @[Mux.scala 46:19:@9068.4]
  wire [7:0] _T_11649; // @[Mux.scala 46:16:@9069.4]
  wire  _T_11650; // @[Mux.scala 46:19:@9070.4]
  wire [7:0] _T_11651; // @[Mux.scala 46:16:@9071.4]
  wire  _T_11652; // @[Mux.scala 46:19:@9072.4]
  wire [7:0] _T_11653; // @[Mux.scala 46:16:@9073.4]
  wire  _T_11654; // @[Mux.scala 46:19:@9074.4]
  wire [7:0] _T_11655; // @[Mux.scala 46:16:@9075.4]
  wire  _T_11656; // @[Mux.scala 46:19:@9076.4]
  wire [7:0] _T_11657; // @[Mux.scala 46:16:@9077.4]
  wire  _T_11658; // @[Mux.scala 46:19:@9078.4]
  wire [7:0] _T_11659; // @[Mux.scala 46:16:@9079.4]
  wire  _T_11671; // @[Mux.scala 46:19:@9081.4]
  wire [7:0] _T_11672; // @[Mux.scala 46:16:@9082.4]
  wire  _T_11673; // @[Mux.scala 46:19:@9083.4]
  wire [7:0] _T_11674; // @[Mux.scala 46:16:@9084.4]
  wire  _T_11675; // @[Mux.scala 46:19:@9085.4]
  wire [7:0] _T_11676; // @[Mux.scala 46:16:@9086.4]
  wire  _T_11677; // @[Mux.scala 46:19:@9087.4]
  wire [7:0] _T_11678; // @[Mux.scala 46:16:@9088.4]
  wire  _T_11679; // @[Mux.scala 46:19:@9089.4]
  wire [7:0] _T_11680; // @[Mux.scala 46:16:@9090.4]
  wire  _T_11681; // @[Mux.scala 46:19:@9091.4]
  wire [7:0] _T_11682; // @[Mux.scala 46:16:@9092.4]
  wire  _T_11683; // @[Mux.scala 46:19:@9093.4]
  wire [7:0] _T_11684; // @[Mux.scala 46:16:@9094.4]
  wire  _T_11685; // @[Mux.scala 46:19:@9095.4]
  wire [7:0] _T_11686; // @[Mux.scala 46:16:@9096.4]
  wire  _T_11687; // @[Mux.scala 46:19:@9097.4]
  wire [7:0] _T_11688; // @[Mux.scala 46:16:@9098.4]
  wire  _T_11689; // @[Mux.scala 46:19:@9099.4]
  wire [7:0] _T_11690; // @[Mux.scala 46:16:@9100.4]
  wire  _T_11703; // @[Mux.scala 46:19:@9102.4]
  wire [7:0] _T_11704; // @[Mux.scala 46:16:@9103.4]
  wire  _T_11705; // @[Mux.scala 46:19:@9104.4]
  wire [7:0] _T_11706; // @[Mux.scala 46:16:@9105.4]
  wire  _T_11707; // @[Mux.scala 46:19:@9106.4]
  wire [7:0] _T_11708; // @[Mux.scala 46:16:@9107.4]
  wire  _T_11709; // @[Mux.scala 46:19:@9108.4]
  wire [7:0] _T_11710; // @[Mux.scala 46:16:@9109.4]
  wire  _T_11711; // @[Mux.scala 46:19:@9110.4]
  wire [7:0] _T_11712; // @[Mux.scala 46:16:@9111.4]
  wire  _T_11713; // @[Mux.scala 46:19:@9112.4]
  wire [7:0] _T_11714; // @[Mux.scala 46:16:@9113.4]
  wire  _T_11715; // @[Mux.scala 46:19:@9114.4]
  wire [7:0] _T_11716; // @[Mux.scala 46:16:@9115.4]
  wire  _T_11717; // @[Mux.scala 46:19:@9116.4]
  wire [7:0] _T_11718; // @[Mux.scala 46:16:@9117.4]
  wire  _T_11719; // @[Mux.scala 46:19:@9118.4]
  wire [7:0] _T_11720; // @[Mux.scala 46:16:@9119.4]
  wire  _T_11721; // @[Mux.scala 46:19:@9120.4]
  wire [7:0] _T_11722; // @[Mux.scala 46:16:@9121.4]
  wire  _T_11723; // @[Mux.scala 46:19:@9122.4]
  wire [7:0] _T_11724; // @[Mux.scala 46:16:@9123.4]
  wire  _T_11738; // @[Mux.scala 46:19:@9125.4]
  wire [7:0] _T_11739; // @[Mux.scala 46:16:@9126.4]
  wire  _T_11740; // @[Mux.scala 46:19:@9127.4]
  wire [7:0] _T_11741; // @[Mux.scala 46:16:@9128.4]
  wire  _T_11742; // @[Mux.scala 46:19:@9129.4]
  wire [7:0] _T_11743; // @[Mux.scala 46:16:@9130.4]
  wire  _T_11744; // @[Mux.scala 46:19:@9131.4]
  wire [7:0] _T_11745; // @[Mux.scala 46:16:@9132.4]
  wire  _T_11746; // @[Mux.scala 46:19:@9133.4]
  wire [7:0] _T_11747; // @[Mux.scala 46:16:@9134.4]
  wire  _T_11748; // @[Mux.scala 46:19:@9135.4]
  wire [7:0] _T_11749; // @[Mux.scala 46:16:@9136.4]
  wire  _T_11750; // @[Mux.scala 46:19:@9137.4]
  wire [7:0] _T_11751; // @[Mux.scala 46:16:@9138.4]
  wire  _T_11752; // @[Mux.scala 46:19:@9139.4]
  wire [7:0] _T_11753; // @[Mux.scala 46:16:@9140.4]
  wire  _T_11754; // @[Mux.scala 46:19:@9141.4]
  wire [7:0] _T_11755; // @[Mux.scala 46:16:@9142.4]
  wire  _T_11756; // @[Mux.scala 46:19:@9143.4]
  wire [7:0] _T_11757; // @[Mux.scala 46:16:@9144.4]
  wire  _T_11758; // @[Mux.scala 46:19:@9145.4]
  wire [7:0] _T_11759; // @[Mux.scala 46:16:@9146.4]
  wire  _T_11760; // @[Mux.scala 46:19:@9147.4]
  wire [7:0] _T_11761; // @[Mux.scala 46:16:@9148.4]
  wire  _T_11776; // @[Mux.scala 46:19:@9150.4]
  wire [7:0] _T_11777; // @[Mux.scala 46:16:@9151.4]
  wire  _T_11778; // @[Mux.scala 46:19:@9152.4]
  wire [7:0] _T_11779; // @[Mux.scala 46:16:@9153.4]
  wire  _T_11780; // @[Mux.scala 46:19:@9154.4]
  wire [7:0] _T_11781; // @[Mux.scala 46:16:@9155.4]
  wire  _T_11782; // @[Mux.scala 46:19:@9156.4]
  wire [7:0] _T_11783; // @[Mux.scala 46:16:@9157.4]
  wire  _T_11784; // @[Mux.scala 46:19:@9158.4]
  wire [7:0] _T_11785; // @[Mux.scala 46:16:@9159.4]
  wire  _T_11786; // @[Mux.scala 46:19:@9160.4]
  wire [7:0] _T_11787; // @[Mux.scala 46:16:@9161.4]
  wire  _T_11788; // @[Mux.scala 46:19:@9162.4]
  wire [7:0] _T_11789; // @[Mux.scala 46:16:@9163.4]
  wire  _T_11790; // @[Mux.scala 46:19:@9164.4]
  wire [7:0] _T_11791; // @[Mux.scala 46:16:@9165.4]
  wire  _T_11792; // @[Mux.scala 46:19:@9166.4]
  wire [7:0] _T_11793; // @[Mux.scala 46:16:@9167.4]
  wire  _T_11794; // @[Mux.scala 46:19:@9168.4]
  wire [7:0] _T_11795; // @[Mux.scala 46:16:@9169.4]
  wire  _T_11796; // @[Mux.scala 46:19:@9170.4]
  wire [7:0] _T_11797; // @[Mux.scala 46:16:@9171.4]
  wire  _T_11798; // @[Mux.scala 46:19:@9172.4]
  wire [7:0] _T_11799; // @[Mux.scala 46:16:@9173.4]
  wire  _T_11800; // @[Mux.scala 46:19:@9174.4]
  wire [7:0] _T_11801; // @[Mux.scala 46:16:@9175.4]
  wire  _T_11817; // @[Mux.scala 46:19:@9177.4]
  wire [7:0] _T_11818; // @[Mux.scala 46:16:@9178.4]
  wire  _T_11819; // @[Mux.scala 46:19:@9179.4]
  wire [7:0] _T_11820; // @[Mux.scala 46:16:@9180.4]
  wire  _T_11821; // @[Mux.scala 46:19:@9181.4]
  wire [7:0] _T_11822; // @[Mux.scala 46:16:@9182.4]
  wire  _T_11823; // @[Mux.scala 46:19:@9183.4]
  wire [7:0] _T_11824; // @[Mux.scala 46:16:@9184.4]
  wire  _T_11825; // @[Mux.scala 46:19:@9185.4]
  wire [7:0] _T_11826; // @[Mux.scala 46:16:@9186.4]
  wire  _T_11827; // @[Mux.scala 46:19:@9187.4]
  wire [7:0] _T_11828; // @[Mux.scala 46:16:@9188.4]
  wire  _T_11829; // @[Mux.scala 46:19:@9189.4]
  wire [7:0] _T_11830; // @[Mux.scala 46:16:@9190.4]
  wire  _T_11831; // @[Mux.scala 46:19:@9191.4]
  wire [7:0] _T_11832; // @[Mux.scala 46:16:@9192.4]
  wire  _T_11833; // @[Mux.scala 46:19:@9193.4]
  wire [7:0] _T_11834; // @[Mux.scala 46:16:@9194.4]
  wire  _T_11835; // @[Mux.scala 46:19:@9195.4]
  wire [7:0] _T_11836; // @[Mux.scala 46:16:@9196.4]
  wire  _T_11837; // @[Mux.scala 46:19:@9197.4]
  wire [7:0] _T_11838; // @[Mux.scala 46:16:@9198.4]
  wire  _T_11839; // @[Mux.scala 46:19:@9199.4]
  wire [7:0] _T_11840; // @[Mux.scala 46:16:@9200.4]
  wire  _T_11841; // @[Mux.scala 46:19:@9201.4]
  wire [7:0] _T_11842; // @[Mux.scala 46:16:@9202.4]
  wire  _T_11843; // @[Mux.scala 46:19:@9203.4]
  wire [7:0] _T_11844; // @[Mux.scala 46:16:@9204.4]
  wire  _T_11861; // @[Mux.scala 46:19:@9206.4]
  wire [7:0] _T_11862; // @[Mux.scala 46:16:@9207.4]
  wire  _T_11863; // @[Mux.scala 46:19:@9208.4]
  wire [7:0] _T_11864; // @[Mux.scala 46:16:@9209.4]
  wire  _T_11865; // @[Mux.scala 46:19:@9210.4]
  wire [7:0] _T_11866; // @[Mux.scala 46:16:@9211.4]
  wire  _T_11867; // @[Mux.scala 46:19:@9212.4]
  wire [7:0] _T_11868; // @[Mux.scala 46:16:@9213.4]
  wire  _T_11869; // @[Mux.scala 46:19:@9214.4]
  wire [7:0] _T_11870; // @[Mux.scala 46:16:@9215.4]
  wire  _T_11871; // @[Mux.scala 46:19:@9216.4]
  wire [7:0] _T_11872; // @[Mux.scala 46:16:@9217.4]
  wire  _T_11873; // @[Mux.scala 46:19:@9218.4]
  wire [7:0] _T_11874; // @[Mux.scala 46:16:@9219.4]
  wire  _T_11875; // @[Mux.scala 46:19:@9220.4]
  wire [7:0] _T_11876; // @[Mux.scala 46:16:@9221.4]
  wire  _T_11877; // @[Mux.scala 46:19:@9222.4]
  wire [7:0] _T_11878; // @[Mux.scala 46:16:@9223.4]
  wire  _T_11879; // @[Mux.scala 46:19:@9224.4]
  wire [7:0] _T_11880; // @[Mux.scala 46:16:@9225.4]
  wire  _T_11881; // @[Mux.scala 46:19:@9226.4]
  wire [7:0] _T_11882; // @[Mux.scala 46:16:@9227.4]
  wire  _T_11883; // @[Mux.scala 46:19:@9228.4]
  wire [7:0] _T_11884; // @[Mux.scala 46:16:@9229.4]
  wire  _T_11885; // @[Mux.scala 46:19:@9230.4]
  wire [7:0] _T_11886; // @[Mux.scala 46:16:@9231.4]
  wire  _T_11887; // @[Mux.scala 46:19:@9232.4]
  wire [7:0] _T_11888; // @[Mux.scala 46:16:@9233.4]
  wire  _T_11889; // @[Mux.scala 46:19:@9234.4]
  wire [7:0] _T_11890; // @[Mux.scala 46:16:@9235.4]
  wire  _T_11908; // @[Mux.scala 46:19:@9237.4]
  wire [7:0] _T_11909; // @[Mux.scala 46:16:@9238.4]
  wire  _T_11910; // @[Mux.scala 46:19:@9239.4]
  wire [7:0] _T_11911; // @[Mux.scala 46:16:@9240.4]
  wire  _T_11912; // @[Mux.scala 46:19:@9241.4]
  wire [7:0] _T_11913; // @[Mux.scala 46:16:@9242.4]
  wire  _T_11914; // @[Mux.scala 46:19:@9243.4]
  wire [7:0] _T_11915; // @[Mux.scala 46:16:@9244.4]
  wire  _T_11916; // @[Mux.scala 46:19:@9245.4]
  wire [7:0] _T_11917; // @[Mux.scala 46:16:@9246.4]
  wire  _T_11918; // @[Mux.scala 46:19:@9247.4]
  wire [7:0] _T_11919; // @[Mux.scala 46:16:@9248.4]
  wire  _T_11920; // @[Mux.scala 46:19:@9249.4]
  wire [7:0] _T_11921; // @[Mux.scala 46:16:@9250.4]
  wire  _T_11922; // @[Mux.scala 46:19:@9251.4]
  wire [7:0] _T_11923; // @[Mux.scala 46:16:@9252.4]
  wire  _T_11924; // @[Mux.scala 46:19:@9253.4]
  wire [7:0] _T_11925; // @[Mux.scala 46:16:@9254.4]
  wire  _T_11926; // @[Mux.scala 46:19:@9255.4]
  wire [7:0] _T_11927; // @[Mux.scala 46:16:@9256.4]
  wire  _T_11928; // @[Mux.scala 46:19:@9257.4]
  wire [7:0] _T_11929; // @[Mux.scala 46:16:@9258.4]
  wire  _T_11930; // @[Mux.scala 46:19:@9259.4]
  wire [7:0] _T_11931; // @[Mux.scala 46:16:@9260.4]
  wire  _T_11932; // @[Mux.scala 46:19:@9261.4]
  wire [7:0] _T_11933; // @[Mux.scala 46:16:@9262.4]
  wire  _T_11934; // @[Mux.scala 46:19:@9263.4]
  wire [7:0] _T_11935; // @[Mux.scala 46:16:@9264.4]
  wire  _T_11936; // @[Mux.scala 46:19:@9265.4]
  wire [7:0] _T_11937; // @[Mux.scala 46:16:@9266.4]
  wire  _T_11938; // @[Mux.scala 46:19:@9267.4]
  wire [7:0] _T_11939; // @[Mux.scala 46:16:@9268.4]
  wire  _T_11958; // @[Mux.scala 46:19:@9270.4]
  wire [7:0] _T_11959; // @[Mux.scala 46:16:@9271.4]
  wire  _T_11960; // @[Mux.scala 46:19:@9272.4]
  wire [7:0] _T_11961; // @[Mux.scala 46:16:@9273.4]
  wire  _T_11962; // @[Mux.scala 46:19:@9274.4]
  wire [7:0] _T_11963; // @[Mux.scala 46:16:@9275.4]
  wire  _T_11964; // @[Mux.scala 46:19:@9276.4]
  wire [7:0] _T_11965; // @[Mux.scala 46:16:@9277.4]
  wire  _T_11966; // @[Mux.scala 46:19:@9278.4]
  wire [7:0] _T_11967; // @[Mux.scala 46:16:@9279.4]
  wire  _T_11968; // @[Mux.scala 46:19:@9280.4]
  wire [7:0] _T_11969; // @[Mux.scala 46:16:@9281.4]
  wire  _T_11970; // @[Mux.scala 46:19:@9282.4]
  wire [7:0] _T_11971; // @[Mux.scala 46:16:@9283.4]
  wire  _T_11972; // @[Mux.scala 46:19:@9284.4]
  wire [7:0] _T_11973; // @[Mux.scala 46:16:@9285.4]
  wire  _T_11974; // @[Mux.scala 46:19:@9286.4]
  wire [7:0] _T_11975; // @[Mux.scala 46:16:@9287.4]
  wire  _T_11976; // @[Mux.scala 46:19:@9288.4]
  wire [7:0] _T_11977; // @[Mux.scala 46:16:@9289.4]
  wire  _T_11978; // @[Mux.scala 46:19:@9290.4]
  wire [7:0] _T_11979; // @[Mux.scala 46:16:@9291.4]
  wire  _T_11980; // @[Mux.scala 46:19:@9292.4]
  wire [7:0] _T_11981; // @[Mux.scala 46:16:@9293.4]
  wire  _T_11982; // @[Mux.scala 46:19:@9294.4]
  wire [7:0] _T_11983; // @[Mux.scala 46:16:@9295.4]
  wire  _T_11984; // @[Mux.scala 46:19:@9296.4]
  wire [7:0] _T_11985; // @[Mux.scala 46:16:@9297.4]
  wire  _T_11986; // @[Mux.scala 46:19:@9298.4]
  wire [7:0] _T_11987; // @[Mux.scala 46:16:@9299.4]
  wire  _T_11988; // @[Mux.scala 46:19:@9300.4]
  wire [7:0] _T_11989; // @[Mux.scala 46:16:@9301.4]
  wire  _T_11990; // @[Mux.scala 46:19:@9302.4]
  wire [7:0] _T_11991; // @[Mux.scala 46:16:@9303.4]
  wire  _T_12011; // @[Mux.scala 46:19:@9305.4]
  wire [7:0] _T_12012; // @[Mux.scala 46:16:@9306.4]
  wire  _T_12013; // @[Mux.scala 46:19:@9307.4]
  wire [7:0] _T_12014; // @[Mux.scala 46:16:@9308.4]
  wire  _T_12015; // @[Mux.scala 46:19:@9309.4]
  wire [7:0] _T_12016; // @[Mux.scala 46:16:@9310.4]
  wire  _T_12017; // @[Mux.scala 46:19:@9311.4]
  wire [7:0] _T_12018; // @[Mux.scala 46:16:@9312.4]
  wire  _T_12019; // @[Mux.scala 46:19:@9313.4]
  wire [7:0] _T_12020; // @[Mux.scala 46:16:@9314.4]
  wire  _T_12021; // @[Mux.scala 46:19:@9315.4]
  wire [7:0] _T_12022; // @[Mux.scala 46:16:@9316.4]
  wire  _T_12023; // @[Mux.scala 46:19:@9317.4]
  wire [7:0] _T_12024; // @[Mux.scala 46:16:@9318.4]
  wire  _T_12025; // @[Mux.scala 46:19:@9319.4]
  wire [7:0] _T_12026; // @[Mux.scala 46:16:@9320.4]
  wire  _T_12027; // @[Mux.scala 46:19:@9321.4]
  wire [7:0] _T_12028; // @[Mux.scala 46:16:@9322.4]
  wire  _T_12029; // @[Mux.scala 46:19:@9323.4]
  wire [7:0] _T_12030; // @[Mux.scala 46:16:@9324.4]
  wire  _T_12031; // @[Mux.scala 46:19:@9325.4]
  wire [7:0] _T_12032; // @[Mux.scala 46:16:@9326.4]
  wire  _T_12033; // @[Mux.scala 46:19:@9327.4]
  wire [7:0] _T_12034; // @[Mux.scala 46:16:@9328.4]
  wire  _T_12035; // @[Mux.scala 46:19:@9329.4]
  wire [7:0] _T_12036; // @[Mux.scala 46:16:@9330.4]
  wire  _T_12037; // @[Mux.scala 46:19:@9331.4]
  wire [7:0] _T_12038; // @[Mux.scala 46:16:@9332.4]
  wire  _T_12039; // @[Mux.scala 46:19:@9333.4]
  wire [7:0] _T_12040; // @[Mux.scala 46:16:@9334.4]
  wire  _T_12041; // @[Mux.scala 46:19:@9335.4]
  wire [7:0] _T_12042; // @[Mux.scala 46:16:@9336.4]
  wire  _T_12043; // @[Mux.scala 46:19:@9337.4]
  wire [7:0] _T_12044; // @[Mux.scala 46:16:@9338.4]
  wire  _T_12045; // @[Mux.scala 46:19:@9339.4]
  wire [7:0] _T_12046; // @[Mux.scala 46:16:@9340.4]
  wire  _T_12067; // @[Mux.scala 46:19:@9342.4]
  wire [7:0] _T_12068; // @[Mux.scala 46:16:@9343.4]
  wire  _T_12069; // @[Mux.scala 46:19:@9344.4]
  wire [7:0] _T_12070; // @[Mux.scala 46:16:@9345.4]
  wire  _T_12071; // @[Mux.scala 46:19:@9346.4]
  wire [7:0] _T_12072; // @[Mux.scala 46:16:@9347.4]
  wire  _T_12073; // @[Mux.scala 46:19:@9348.4]
  wire [7:0] _T_12074; // @[Mux.scala 46:16:@9349.4]
  wire  _T_12075; // @[Mux.scala 46:19:@9350.4]
  wire [7:0] _T_12076; // @[Mux.scala 46:16:@9351.4]
  wire  _T_12077; // @[Mux.scala 46:19:@9352.4]
  wire [7:0] _T_12078; // @[Mux.scala 46:16:@9353.4]
  wire  _T_12079; // @[Mux.scala 46:19:@9354.4]
  wire [7:0] _T_12080; // @[Mux.scala 46:16:@9355.4]
  wire  _T_12081; // @[Mux.scala 46:19:@9356.4]
  wire [7:0] _T_12082; // @[Mux.scala 46:16:@9357.4]
  wire  _T_12083; // @[Mux.scala 46:19:@9358.4]
  wire [7:0] _T_12084; // @[Mux.scala 46:16:@9359.4]
  wire  _T_12085; // @[Mux.scala 46:19:@9360.4]
  wire [7:0] _T_12086; // @[Mux.scala 46:16:@9361.4]
  wire  _T_12087; // @[Mux.scala 46:19:@9362.4]
  wire [7:0] _T_12088; // @[Mux.scala 46:16:@9363.4]
  wire  _T_12089; // @[Mux.scala 46:19:@9364.4]
  wire [7:0] _T_12090; // @[Mux.scala 46:16:@9365.4]
  wire  _T_12091; // @[Mux.scala 46:19:@9366.4]
  wire [7:0] _T_12092; // @[Mux.scala 46:16:@9367.4]
  wire  _T_12093; // @[Mux.scala 46:19:@9368.4]
  wire [7:0] _T_12094; // @[Mux.scala 46:16:@9369.4]
  wire  _T_12095; // @[Mux.scala 46:19:@9370.4]
  wire [7:0] _T_12096; // @[Mux.scala 46:16:@9371.4]
  wire  _T_12097; // @[Mux.scala 46:19:@9372.4]
  wire [7:0] _T_12098; // @[Mux.scala 46:16:@9373.4]
  wire  _T_12099; // @[Mux.scala 46:19:@9374.4]
  wire [7:0] _T_12100; // @[Mux.scala 46:16:@9375.4]
  wire  _T_12101; // @[Mux.scala 46:19:@9376.4]
  wire [7:0] _T_12102; // @[Mux.scala 46:16:@9377.4]
  wire  _T_12103; // @[Mux.scala 46:19:@9378.4]
  wire [7:0] _T_12104; // @[Mux.scala 46:16:@9379.4]
  wire  _T_12126; // @[Mux.scala 46:19:@9381.4]
  wire [7:0] _T_12127; // @[Mux.scala 46:16:@9382.4]
  wire  _T_12128; // @[Mux.scala 46:19:@9383.4]
  wire [7:0] _T_12129; // @[Mux.scala 46:16:@9384.4]
  wire  _T_12130; // @[Mux.scala 46:19:@9385.4]
  wire [7:0] _T_12131; // @[Mux.scala 46:16:@9386.4]
  wire  _T_12132; // @[Mux.scala 46:19:@9387.4]
  wire [7:0] _T_12133; // @[Mux.scala 46:16:@9388.4]
  wire  _T_12134; // @[Mux.scala 46:19:@9389.4]
  wire [7:0] _T_12135; // @[Mux.scala 46:16:@9390.4]
  wire  _T_12136; // @[Mux.scala 46:19:@9391.4]
  wire [7:0] _T_12137; // @[Mux.scala 46:16:@9392.4]
  wire  _T_12138; // @[Mux.scala 46:19:@9393.4]
  wire [7:0] _T_12139; // @[Mux.scala 46:16:@9394.4]
  wire  _T_12140; // @[Mux.scala 46:19:@9395.4]
  wire [7:0] _T_12141; // @[Mux.scala 46:16:@9396.4]
  wire  _T_12142; // @[Mux.scala 46:19:@9397.4]
  wire [7:0] _T_12143; // @[Mux.scala 46:16:@9398.4]
  wire  _T_12144; // @[Mux.scala 46:19:@9399.4]
  wire [7:0] _T_12145; // @[Mux.scala 46:16:@9400.4]
  wire  _T_12146; // @[Mux.scala 46:19:@9401.4]
  wire [7:0] _T_12147; // @[Mux.scala 46:16:@9402.4]
  wire  _T_12148; // @[Mux.scala 46:19:@9403.4]
  wire [7:0] _T_12149; // @[Mux.scala 46:16:@9404.4]
  wire  _T_12150; // @[Mux.scala 46:19:@9405.4]
  wire [7:0] _T_12151; // @[Mux.scala 46:16:@9406.4]
  wire  _T_12152; // @[Mux.scala 46:19:@9407.4]
  wire [7:0] _T_12153; // @[Mux.scala 46:16:@9408.4]
  wire  _T_12154; // @[Mux.scala 46:19:@9409.4]
  wire [7:0] _T_12155; // @[Mux.scala 46:16:@9410.4]
  wire  _T_12156; // @[Mux.scala 46:19:@9411.4]
  wire [7:0] _T_12157; // @[Mux.scala 46:16:@9412.4]
  wire  _T_12158; // @[Mux.scala 46:19:@9413.4]
  wire [7:0] _T_12159; // @[Mux.scala 46:16:@9414.4]
  wire  _T_12160; // @[Mux.scala 46:19:@9415.4]
  wire [7:0] _T_12161; // @[Mux.scala 46:16:@9416.4]
  wire  _T_12162; // @[Mux.scala 46:19:@9417.4]
  wire [7:0] _T_12163; // @[Mux.scala 46:16:@9418.4]
  wire  _T_12164; // @[Mux.scala 46:19:@9419.4]
  wire [7:0] _T_12165; // @[Mux.scala 46:16:@9420.4]
  wire  _T_12188; // @[Mux.scala 46:19:@9422.4]
  wire [7:0] _T_12189; // @[Mux.scala 46:16:@9423.4]
  wire  _T_12190; // @[Mux.scala 46:19:@9424.4]
  wire [7:0] _T_12191; // @[Mux.scala 46:16:@9425.4]
  wire  _T_12192; // @[Mux.scala 46:19:@9426.4]
  wire [7:0] _T_12193; // @[Mux.scala 46:16:@9427.4]
  wire  _T_12194; // @[Mux.scala 46:19:@9428.4]
  wire [7:0] _T_12195; // @[Mux.scala 46:16:@9429.4]
  wire  _T_12196; // @[Mux.scala 46:19:@9430.4]
  wire [7:0] _T_12197; // @[Mux.scala 46:16:@9431.4]
  wire  _T_12198; // @[Mux.scala 46:19:@9432.4]
  wire [7:0] _T_12199; // @[Mux.scala 46:16:@9433.4]
  wire  _T_12200; // @[Mux.scala 46:19:@9434.4]
  wire [7:0] _T_12201; // @[Mux.scala 46:16:@9435.4]
  wire  _T_12202; // @[Mux.scala 46:19:@9436.4]
  wire [7:0] _T_12203; // @[Mux.scala 46:16:@9437.4]
  wire  _T_12204; // @[Mux.scala 46:19:@9438.4]
  wire [7:0] _T_12205; // @[Mux.scala 46:16:@9439.4]
  wire  _T_12206; // @[Mux.scala 46:19:@9440.4]
  wire [7:0] _T_12207; // @[Mux.scala 46:16:@9441.4]
  wire  _T_12208; // @[Mux.scala 46:19:@9442.4]
  wire [7:0] _T_12209; // @[Mux.scala 46:16:@9443.4]
  wire  _T_12210; // @[Mux.scala 46:19:@9444.4]
  wire [7:0] _T_12211; // @[Mux.scala 46:16:@9445.4]
  wire  _T_12212; // @[Mux.scala 46:19:@9446.4]
  wire [7:0] _T_12213; // @[Mux.scala 46:16:@9447.4]
  wire  _T_12214; // @[Mux.scala 46:19:@9448.4]
  wire [7:0] _T_12215; // @[Mux.scala 46:16:@9449.4]
  wire  _T_12216; // @[Mux.scala 46:19:@9450.4]
  wire [7:0] _T_12217; // @[Mux.scala 46:16:@9451.4]
  wire  _T_12218; // @[Mux.scala 46:19:@9452.4]
  wire [7:0] _T_12219; // @[Mux.scala 46:16:@9453.4]
  wire  _T_12220; // @[Mux.scala 46:19:@9454.4]
  wire [7:0] _T_12221; // @[Mux.scala 46:16:@9455.4]
  wire  _T_12222; // @[Mux.scala 46:19:@9456.4]
  wire [7:0] _T_12223; // @[Mux.scala 46:16:@9457.4]
  wire  _T_12224; // @[Mux.scala 46:19:@9458.4]
  wire [7:0] _T_12225; // @[Mux.scala 46:16:@9459.4]
  wire  _T_12226; // @[Mux.scala 46:19:@9460.4]
  wire [7:0] _T_12227; // @[Mux.scala 46:16:@9461.4]
  wire  _T_12228; // @[Mux.scala 46:19:@9462.4]
  wire [7:0] _T_12229; // @[Mux.scala 46:16:@9463.4]
  wire  _T_12253; // @[Mux.scala 46:19:@9465.4]
  wire [7:0] _T_12254; // @[Mux.scala 46:16:@9466.4]
  wire  _T_12255; // @[Mux.scala 46:19:@9467.4]
  wire [7:0] _T_12256; // @[Mux.scala 46:16:@9468.4]
  wire  _T_12257; // @[Mux.scala 46:19:@9469.4]
  wire [7:0] _T_12258; // @[Mux.scala 46:16:@9470.4]
  wire  _T_12259; // @[Mux.scala 46:19:@9471.4]
  wire [7:0] _T_12260; // @[Mux.scala 46:16:@9472.4]
  wire  _T_12261; // @[Mux.scala 46:19:@9473.4]
  wire [7:0] _T_12262; // @[Mux.scala 46:16:@9474.4]
  wire  _T_12263; // @[Mux.scala 46:19:@9475.4]
  wire [7:0] _T_12264; // @[Mux.scala 46:16:@9476.4]
  wire  _T_12265; // @[Mux.scala 46:19:@9477.4]
  wire [7:0] _T_12266; // @[Mux.scala 46:16:@9478.4]
  wire  _T_12267; // @[Mux.scala 46:19:@9479.4]
  wire [7:0] _T_12268; // @[Mux.scala 46:16:@9480.4]
  wire  _T_12269; // @[Mux.scala 46:19:@9481.4]
  wire [7:0] _T_12270; // @[Mux.scala 46:16:@9482.4]
  wire  _T_12271; // @[Mux.scala 46:19:@9483.4]
  wire [7:0] _T_12272; // @[Mux.scala 46:16:@9484.4]
  wire  _T_12273; // @[Mux.scala 46:19:@9485.4]
  wire [7:0] _T_12274; // @[Mux.scala 46:16:@9486.4]
  wire  _T_12275; // @[Mux.scala 46:19:@9487.4]
  wire [7:0] _T_12276; // @[Mux.scala 46:16:@9488.4]
  wire  _T_12277; // @[Mux.scala 46:19:@9489.4]
  wire [7:0] _T_12278; // @[Mux.scala 46:16:@9490.4]
  wire  _T_12279; // @[Mux.scala 46:19:@9491.4]
  wire [7:0] _T_12280; // @[Mux.scala 46:16:@9492.4]
  wire  _T_12281; // @[Mux.scala 46:19:@9493.4]
  wire [7:0] _T_12282; // @[Mux.scala 46:16:@9494.4]
  wire  _T_12283; // @[Mux.scala 46:19:@9495.4]
  wire [7:0] _T_12284; // @[Mux.scala 46:16:@9496.4]
  wire  _T_12285; // @[Mux.scala 46:19:@9497.4]
  wire [7:0] _T_12286; // @[Mux.scala 46:16:@9498.4]
  wire  _T_12287; // @[Mux.scala 46:19:@9499.4]
  wire [7:0] _T_12288; // @[Mux.scala 46:16:@9500.4]
  wire  _T_12289; // @[Mux.scala 46:19:@9501.4]
  wire [7:0] _T_12290; // @[Mux.scala 46:16:@9502.4]
  wire  _T_12291; // @[Mux.scala 46:19:@9503.4]
  wire [7:0] _T_12292; // @[Mux.scala 46:16:@9504.4]
  wire  _T_12293; // @[Mux.scala 46:19:@9505.4]
  wire [7:0] _T_12294; // @[Mux.scala 46:16:@9506.4]
  wire  _T_12295; // @[Mux.scala 46:19:@9507.4]
  wire [7:0] _T_12296; // @[Mux.scala 46:16:@9508.4]
  wire  _T_12321; // @[Mux.scala 46:19:@9510.4]
  wire [7:0] _T_12322; // @[Mux.scala 46:16:@9511.4]
  wire  _T_12323; // @[Mux.scala 46:19:@9512.4]
  wire [7:0] _T_12324; // @[Mux.scala 46:16:@9513.4]
  wire  _T_12325; // @[Mux.scala 46:19:@9514.4]
  wire [7:0] _T_12326; // @[Mux.scala 46:16:@9515.4]
  wire  _T_12327; // @[Mux.scala 46:19:@9516.4]
  wire [7:0] _T_12328; // @[Mux.scala 46:16:@9517.4]
  wire  _T_12329; // @[Mux.scala 46:19:@9518.4]
  wire [7:0] _T_12330; // @[Mux.scala 46:16:@9519.4]
  wire  _T_12331; // @[Mux.scala 46:19:@9520.4]
  wire [7:0] _T_12332; // @[Mux.scala 46:16:@9521.4]
  wire  _T_12333; // @[Mux.scala 46:19:@9522.4]
  wire [7:0] _T_12334; // @[Mux.scala 46:16:@9523.4]
  wire  _T_12335; // @[Mux.scala 46:19:@9524.4]
  wire [7:0] _T_12336; // @[Mux.scala 46:16:@9525.4]
  wire  _T_12337; // @[Mux.scala 46:19:@9526.4]
  wire [7:0] _T_12338; // @[Mux.scala 46:16:@9527.4]
  wire  _T_12339; // @[Mux.scala 46:19:@9528.4]
  wire [7:0] _T_12340; // @[Mux.scala 46:16:@9529.4]
  wire  _T_12341; // @[Mux.scala 46:19:@9530.4]
  wire [7:0] _T_12342; // @[Mux.scala 46:16:@9531.4]
  wire  _T_12343; // @[Mux.scala 46:19:@9532.4]
  wire [7:0] _T_12344; // @[Mux.scala 46:16:@9533.4]
  wire  _T_12345; // @[Mux.scala 46:19:@9534.4]
  wire [7:0] _T_12346; // @[Mux.scala 46:16:@9535.4]
  wire  _T_12347; // @[Mux.scala 46:19:@9536.4]
  wire [7:0] _T_12348; // @[Mux.scala 46:16:@9537.4]
  wire  _T_12349; // @[Mux.scala 46:19:@9538.4]
  wire [7:0] _T_12350; // @[Mux.scala 46:16:@9539.4]
  wire  _T_12351; // @[Mux.scala 46:19:@9540.4]
  wire [7:0] _T_12352; // @[Mux.scala 46:16:@9541.4]
  wire  _T_12353; // @[Mux.scala 46:19:@9542.4]
  wire [7:0] _T_12354; // @[Mux.scala 46:16:@9543.4]
  wire  _T_12355; // @[Mux.scala 46:19:@9544.4]
  wire [7:0] _T_12356; // @[Mux.scala 46:16:@9545.4]
  wire  _T_12357; // @[Mux.scala 46:19:@9546.4]
  wire [7:0] _T_12358; // @[Mux.scala 46:16:@9547.4]
  wire  _T_12359; // @[Mux.scala 46:19:@9548.4]
  wire [7:0] _T_12360; // @[Mux.scala 46:16:@9549.4]
  wire  _T_12361; // @[Mux.scala 46:19:@9550.4]
  wire [7:0] _T_12362; // @[Mux.scala 46:16:@9551.4]
  wire  _T_12363; // @[Mux.scala 46:19:@9552.4]
  wire [7:0] _T_12364; // @[Mux.scala 46:16:@9553.4]
  wire  _T_12365; // @[Mux.scala 46:19:@9554.4]
  wire [7:0] _T_12366; // @[Mux.scala 46:16:@9555.4]
  wire  _T_12392; // @[Mux.scala 46:19:@9557.4]
  wire [7:0] _T_12393; // @[Mux.scala 46:16:@9558.4]
  wire  _T_12394; // @[Mux.scala 46:19:@9559.4]
  wire [7:0] _T_12395; // @[Mux.scala 46:16:@9560.4]
  wire  _T_12396; // @[Mux.scala 46:19:@9561.4]
  wire [7:0] _T_12397; // @[Mux.scala 46:16:@9562.4]
  wire  _T_12398; // @[Mux.scala 46:19:@9563.4]
  wire [7:0] _T_12399; // @[Mux.scala 46:16:@9564.4]
  wire  _T_12400; // @[Mux.scala 46:19:@9565.4]
  wire [7:0] _T_12401; // @[Mux.scala 46:16:@9566.4]
  wire  _T_12402; // @[Mux.scala 46:19:@9567.4]
  wire [7:0] _T_12403; // @[Mux.scala 46:16:@9568.4]
  wire  _T_12404; // @[Mux.scala 46:19:@9569.4]
  wire [7:0] _T_12405; // @[Mux.scala 46:16:@9570.4]
  wire  _T_12406; // @[Mux.scala 46:19:@9571.4]
  wire [7:0] _T_12407; // @[Mux.scala 46:16:@9572.4]
  wire  _T_12408; // @[Mux.scala 46:19:@9573.4]
  wire [7:0] _T_12409; // @[Mux.scala 46:16:@9574.4]
  wire  _T_12410; // @[Mux.scala 46:19:@9575.4]
  wire [7:0] _T_12411; // @[Mux.scala 46:16:@9576.4]
  wire  _T_12412; // @[Mux.scala 46:19:@9577.4]
  wire [7:0] _T_12413; // @[Mux.scala 46:16:@9578.4]
  wire  _T_12414; // @[Mux.scala 46:19:@9579.4]
  wire [7:0] _T_12415; // @[Mux.scala 46:16:@9580.4]
  wire  _T_12416; // @[Mux.scala 46:19:@9581.4]
  wire [7:0] _T_12417; // @[Mux.scala 46:16:@9582.4]
  wire  _T_12418; // @[Mux.scala 46:19:@9583.4]
  wire [7:0] _T_12419; // @[Mux.scala 46:16:@9584.4]
  wire  _T_12420; // @[Mux.scala 46:19:@9585.4]
  wire [7:0] _T_12421; // @[Mux.scala 46:16:@9586.4]
  wire  _T_12422; // @[Mux.scala 46:19:@9587.4]
  wire [7:0] _T_12423; // @[Mux.scala 46:16:@9588.4]
  wire  _T_12424; // @[Mux.scala 46:19:@9589.4]
  wire [7:0] _T_12425; // @[Mux.scala 46:16:@9590.4]
  wire  _T_12426; // @[Mux.scala 46:19:@9591.4]
  wire [7:0] _T_12427; // @[Mux.scala 46:16:@9592.4]
  wire  _T_12428; // @[Mux.scala 46:19:@9593.4]
  wire [7:0] _T_12429; // @[Mux.scala 46:16:@9594.4]
  wire  _T_12430; // @[Mux.scala 46:19:@9595.4]
  wire [7:0] _T_12431; // @[Mux.scala 46:16:@9596.4]
  wire  _T_12432; // @[Mux.scala 46:19:@9597.4]
  wire [7:0] _T_12433; // @[Mux.scala 46:16:@9598.4]
  wire  _T_12434; // @[Mux.scala 46:19:@9599.4]
  wire [7:0] _T_12435; // @[Mux.scala 46:16:@9600.4]
  wire  _T_12436; // @[Mux.scala 46:19:@9601.4]
  wire [7:0] _T_12437; // @[Mux.scala 46:16:@9602.4]
  wire  _T_12438; // @[Mux.scala 46:19:@9603.4]
  wire [7:0] _T_12439; // @[Mux.scala 46:16:@9604.4]
  wire  _T_12466; // @[Mux.scala 46:19:@9606.4]
  wire [7:0] _T_12467; // @[Mux.scala 46:16:@9607.4]
  wire  _T_12468; // @[Mux.scala 46:19:@9608.4]
  wire [7:0] _T_12469; // @[Mux.scala 46:16:@9609.4]
  wire  _T_12470; // @[Mux.scala 46:19:@9610.4]
  wire [7:0] _T_12471; // @[Mux.scala 46:16:@9611.4]
  wire  _T_12472; // @[Mux.scala 46:19:@9612.4]
  wire [7:0] _T_12473; // @[Mux.scala 46:16:@9613.4]
  wire  _T_12474; // @[Mux.scala 46:19:@9614.4]
  wire [7:0] _T_12475; // @[Mux.scala 46:16:@9615.4]
  wire  _T_12476; // @[Mux.scala 46:19:@9616.4]
  wire [7:0] _T_12477; // @[Mux.scala 46:16:@9617.4]
  wire  _T_12478; // @[Mux.scala 46:19:@9618.4]
  wire [7:0] _T_12479; // @[Mux.scala 46:16:@9619.4]
  wire  _T_12480; // @[Mux.scala 46:19:@9620.4]
  wire [7:0] _T_12481; // @[Mux.scala 46:16:@9621.4]
  wire  _T_12482; // @[Mux.scala 46:19:@9622.4]
  wire [7:0] _T_12483; // @[Mux.scala 46:16:@9623.4]
  wire  _T_12484; // @[Mux.scala 46:19:@9624.4]
  wire [7:0] _T_12485; // @[Mux.scala 46:16:@9625.4]
  wire  _T_12486; // @[Mux.scala 46:19:@9626.4]
  wire [7:0] _T_12487; // @[Mux.scala 46:16:@9627.4]
  wire  _T_12488; // @[Mux.scala 46:19:@9628.4]
  wire [7:0] _T_12489; // @[Mux.scala 46:16:@9629.4]
  wire  _T_12490; // @[Mux.scala 46:19:@9630.4]
  wire [7:0] _T_12491; // @[Mux.scala 46:16:@9631.4]
  wire  _T_12492; // @[Mux.scala 46:19:@9632.4]
  wire [7:0] _T_12493; // @[Mux.scala 46:16:@9633.4]
  wire  _T_12494; // @[Mux.scala 46:19:@9634.4]
  wire [7:0] _T_12495; // @[Mux.scala 46:16:@9635.4]
  wire  _T_12496; // @[Mux.scala 46:19:@9636.4]
  wire [7:0] _T_12497; // @[Mux.scala 46:16:@9637.4]
  wire  _T_12498; // @[Mux.scala 46:19:@9638.4]
  wire [7:0] _T_12499; // @[Mux.scala 46:16:@9639.4]
  wire  _T_12500; // @[Mux.scala 46:19:@9640.4]
  wire [7:0] _T_12501; // @[Mux.scala 46:16:@9641.4]
  wire  _T_12502; // @[Mux.scala 46:19:@9642.4]
  wire [7:0] _T_12503; // @[Mux.scala 46:16:@9643.4]
  wire  _T_12504; // @[Mux.scala 46:19:@9644.4]
  wire [7:0] _T_12505; // @[Mux.scala 46:16:@9645.4]
  wire  _T_12506; // @[Mux.scala 46:19:@9646.4]
  wire [7:0] _T_12507; // @[Mux.scala 46:16:@9647.4]
  wire  _T_12508; // @[Mux.scala 46:19:@9648.4]
  wire [7:0] _T_12509; // @[Mux.scala 46:16:@9649.4]
  wire  _T_12510; // @[Mux.scala 46:19:@9650.4]
  wire [7:0] _T_12511; // @[Mux.scala 46:16:@9651.4]
  wire  _T_12512; // @[Mux.scala 46:19:@9652.4]
  wire [7:0] _T_12513; // @[Mux.scala 46:16:@9653.4]
  wire  _T_12514; // @[Mux.scala 46:19:@9654.4]
  wire [7:0] _T_12515; // @[Mux.scala 46:16:@9655.4]
  wire  _T_12543; // @[Mux.scala 46:19:@9657.4]
  wire [7:0] _T_12544; // @[Mux.scala 46:16:@9658.4]
  wire  _T_12545; // @[Mux.scala 46:19:@9659.4]
  wire [7:0] _T_12546; // @[Mux.scala 46:16:@9660.4]
  wire  _T_12547; // @[Mux.scala 46:19:@9661.4]
  wire [7:0] _T_12548; // @[Mux.scala 46:16:@9662.4]
  wire  _T_12549; // @[Mux.scala 46:19:@9663.4]
  wire [7:0] _T_12550; // @[Mux.scala 46:16:@9664.4]
  wire  _T_12551; // @[Mux.scala 46:19:@9665.4]
  wire [7:0] _T_12552; // @[Mux.scala 46:16:@9666.4]
  wire  _T_12553; // @[Mux.scala 46:19:@9667.4]
  wire [7:0] _T_12554; // @[Mux.scala 46:16:@9668.4]
  wire  _T_12555; // @[Mux.scala 46:19:@9669.4]
  wire [7:0] _T_12556; // @[Mux.scala 46:16:@9670.4]
  wire  _T_12557; // @[Mux.scala 46:19:@9671.4]
  wire [7:0] _T_12558; // @[Mux.scala 46:16:@9672.4]
  wire  _T_12559; // @[Mux.scala 46:19:@9673.4]
  wire [7:0] _T_12560; // @[Mux.scala 46:16:@9674.4]
  wire  _T_12561; // @[Mux.scala 46:19:@9675.4]
  wire [7:0] _T_12562; // @[Mux.scala 46:16:@9676.4]
  wire  _T_12563; // @[Mux.scala 46:19:@9677.4]
  wire [7:0] _T_12564; // @[Mux.scala 46:16:@9678.4]
  wire  _T_12565; // @[Mux.scala 46:19:@9679.4]
  wire [7:0] _T_12566; // @[Mux.scala 46:16:@9680.4]
  wire  _T_12567; // @[Mux.scala 46:19:@9681.4]
  wire [7:0] _T_12568; // @[Mux.scala 46:16:@9682.4]
  wire  _T_12569; // @[Mux.scala 46:19:@9683.4]
  wire [7:0] _T_12570; // @[Mux.scala 46:16:@9684.4]
  wire  _T_12571; // @[Mux.scala 46:19:@9685.4]
  wire [7:0] _T_12572; // @[Mux.scala 46:16:@9686.4]
  wire  _T_12573; // @[Mux.scala 46:19:@9687.4]
  wire [7:0] _T_12574; // @[Mux.scala 46:16:@9688.4]
  wire  _T_12575; // @[Mux.scala 46:19:@9689.4]
  wire [7:0] _T_12576; // @[Mux.scala 46:16:@9690.4]
  wire  _T_12577; // @[Mux.scala 46:19:@9691.4]
  wire [7:0] _T_12578; // @[Mux.scala 46:16:@9692.4]
  wire  _T_12579; // @[Mux.scala 46:19:@9693.4]
  wire [7:0] _T_12580; // @[Mux.scala 46:16:@9694.4]
  wire  _T_12581; // @[Mux.scala 46:19:@9695.4]
  wire [7:0] _T_12582; // @[Mux.scala 46:16:@9696.4]
  wire  _T_12583; // @[Mux.scala 46:19:@9697.4]
  wire [7:0] _T_12584; // @[Mux.scala 46:16:@9698.4]
  wire  _T_12585; // @[Mux.scala 46:19:@9699.4]
  wire [7:0] _T_12586; // @[Mux.scala 46:16:@9700.4]
  wire  _T_12587; // @[Mux.scala 46:19:@9701.4]
  wire [7:0] _T_12588; // @[Mux.scala 46:16:@9702.4]
  wire  _T_12589; // @[Mux.scala 46:19:@9703.4]
  wire [7:0] _T_12590; // @[Mux.scala 46:16:@9704.4]
  wire  _T_12591; // @[Mux.scala 46:19:@9705.4]
  wire [7:0] _T_12592; // @[Mux.scala 46:16:@9706.4]
  wire  _T_12593; // @[Mux.scala 46:19:@9707.4]
  wire [7:0] _T_12594; // @[Mux.scala 46:16:@9708.4]
  wire  _T_12623; // @[Mux.scala 46:19:@9710.4]
  wire [7:0] _T_12624; // @[Mux.scala 46:16:@9711.4]
  wire  _T_12625; // @[Mux.scala 46:19:@9712.4]
  wire [7:0] _T_12626; // @[Mux.scala 46:16:@9713.4]
  wire  _T_12627; // @[Mux.scala 46:19:@9714.4]
  wire [7:0] _T_12628; // @[Mux.scala 46:16:@9715.4]
  wire  _T_12629; // @[Mux.scala 46:19:@9716.4]
  wire [7:0] _T_12630; // @[Mux.scala 46:16:@9717.4]
  wire  _T_12631; // @[Mux.scala 46:19:@9718.4]
  wire [7:0] _T_12632; // @[Mux.scala 46:16:@9719.4]
  wire  _T_12633; // @[Mux.scala 46:19:@9720.4]
  wire [7:0] _T_12634; // @[Mux.scala 46:16:@9721.4]
  wire  _T_12635; // @[Mux.scala 46:19:@9722.4]
  wire [7:0] _T_12636; // @[Mux.scala 46:16:@9723.4]
  wire  _T_12637; // @[Mux.scala 46:19:@9724.4]
  wire [7:0] _T_12638; // @[Mux.scala 46:16:@9725.4]
  wire  _T_12639; // @[Mux.scala 46:19:@9726.4]
  wire [7:0] _T_12640; // @[Mux.scala 46:16:@9727.4]
  wire  _T_12641; // @[Mux.scala 46:19:@9728.4]
  wire [7:0] _T_12642; // @[Mux.scala 46:16:@9729.4]
  wire  _T_12643; // @[Mux.scala 46:19:@9730.4]
  wire [7:0] _T_12644; // @[Mux.scala 46:16:@9731.4]
  wire  _T_12645; // @[Mux.scala 46:19:@9732.4]
  wire [7:0] _T_12646; // @[Mux.scala 46:16:@9733.4]
  wire  _T_12647; // @[Mux.scala 46:19:@9734.4]
  wire [7:0] _T_12648; // @[Mux.scala 46:16:@9735.4]
  wire  _T_12649; // @[Mux.scala 46:19:@9736.4]
  wire [7:0] _T_12650; // @[Mux.scala 46:16:@9737.4]
  wire  _T_12651; // @[Mux.scala 46:19:@9738.4]
  wire [7:0] _T_12652; // @[Mux.scala 46:16:@9739.4]
  wire  _T_12653; // @[Mux.scala 46:19:@9740.4]
  wire [7:0] _T_12654; // @[Mux.scala 46:16:@9741.4]
  wire  _T_12655; // @[Mux.scala 46:19:@9742.4]
  wire [7:0] _T_12656; // @[Mux.scala 46:16:@9743.4]
  wire  _T_12657; // @[Mux.scala 46:19:@9744.4]
  wire [7:0] _T_12658; // @[Mux.scala 46:16:@9745.4]
  wire  _T_12659; // @[Mux.scala 46:19:@9746.4]
  wire [7:0] _T_12660; // @[Mux.scala 46:16:@9747.4]
  wire  _T_12661; // @[Mux.scala 46:19:@9748.4]
  wire [7:0] _T_12662; // @[Mux.scala 46:16:@9749.4]
  wire  _T_12663; // @[Mux.scala 46:19:@9750.4]
  wire [7:0] _T_12664; // @[Mux.scala 46:16:@9751.4]
  wire  _T_12665; // @[Mux.scala 46:19:@9752.4]
  wire [7:0] _T_12666; // @[Mux.scala 46:16:@9753.4]
  wire  _T_12667; // @[Mux.scala 46:19:@9754.4]
  wire [7:0] _T_12668; // @[Mux.scala 46:16:@9755.4]
  wire  _T_12669; // @[Mux.scala 46:19:@9756.4]
  wire [7:0] _T_12670; // @[Mux.scala 46:16:@9757.4]
  wire  _T_12671; // @[Mux.scala 46:19:@9758.4]
  wire [7:0] _T_12672; // @[Mux.scala 46:16:@9759.4]
  wire  _T_12673; // @[Mux.scala 46:19:@9760.4]
  wire [7:0] _T_12674; // @[Mux.scala 46:16:@9761.4]
  wire  _T_12675; // @[Mux.scala 46:19:@9762.4]
  wire [7:0] _T_12676; // @[Mux.scala 46:16:@9763.4]
  wire  _T_12706; // @[Mux.scala 46:19:@9765.4]
  wire [7:0] _T_12707; // @[Mux.scala 46:16:@9766.4]
  wire  _T_12708; // @[Mux.scala 46:19:@9767.4]
  wire [7:0] _T_12709; // @[Mux.scala 46:16:@9768.4]
  wire  _T_12710; // @[Mux.scala 46:19:@9769.4]
  wire [7:0] _T_12711; // @[Mux.scala 46:16:@9770.4]
  wire  _T_12712; // @[Mux.scala 46:19:@9771.4]
  wire [7:0] _T_12713; // @[Mux.scala 46:16:@9772.4]
  wire  _T_12714; // @[Mux.scala 46:19:@9773.4]
  wire [7:0] _T_12715; // @[Mux.scala 46:16:@9774.4]
  wire  _T_12716; // @[Mux.scala 46:19:@9775.4]
  wire [7:0] _T_12717; // @[Mux.scala 46:16:@9776.4]
  wire  _T_12718; // @[Mux.scala 46:19:@9777.4]
  wire [7:0] _T_12719; // @[Mux.scala 46:16:@9778.4]
  wire  _T_12720; // @[Mux.scala 46:19:@9779.4]
  wire [7:0] _T_12721; // @[Mux.scala 46:16:@9780.4]
  wire  _T_12722; // @[Mux.scala 46:19:@9781.4]
  wire [7:0] _T_12723; // @[Mux.scala 46:16:@9782.4]
  wire  _T_12724; // @[Mux.scala 46:19:@9783.4]
  wire [7:0] _T_12725; // @[Mux.scala 46:16:@9784.4]
  wire  _T_12726; // @[Mux.scala 46:19:@9785.4]
  wire [7:0] _T_12727; // @[Mux.scala 46:16:@9786.4]
  wire  _T_12728; // @[Mux.scala 46:19:@9787.4]
  wire [7:0] _T_12729; // @[Mux.scala 46:16:@9788.4]
  wire  _T_12730; // @[Mux.scala 46:19:@9789.4]
  wire [7:0] _T_12731; // @[Mux.scala 46:16:@9790.4]
  wire  _T_12732; // @[Mux.scala 46:19:@9791.4]
  wire [7:0] _T_12733; // @[Mux.scala 46:16:@9792.4]
  wire  _T_12734; // @[Mux.scala 46:19:@9793.4]
  wire [7:0] _T_12735; // @[Mux.scala 46:16:@9794.4]
  wire  _T_12736; // @[Mux.scala 46:19:@9795.4]
  wire [7:0] _T_12737; // @[Mux.scala 46:16:@9796.4]
  wire  _T_12738; // @[Mux.scala 46:19:@9797.4]
  wire [7:0] _T_12739; // @[Mux.scala 46:16:@9798.4]
  wire  _T_12740; // @[Mux.scala 46:19:@9799.4]
  wire [7:0] _T_12741; // @[Mux.scala 46:16:@9800.4]
  wire  _T_12742; // @[Mux.scala 46:19:@9801.4]
  wire [7:0] _T_12743; // @[Mux.scala 46:16:@9802.4]
  wire  _T_12744; // @[Mux.scala 46:19:@9803.4]
  wire [7:0] _T_12745; // @[Mux.scala 46:16:@9804.4]
  wire  _T_12746; // @[Mux.scala 46:19:@9805.4]
  wire [7:0] _T_12747; // @[Mux.scala 46:16:@9806.4]
  wire  _T_12748; // @[Mux.scala 46:19:@9807.4]
  wire [7:0] _T_12749; // @[Mux.scala 46:16:@9808.4]
  wire  _T_12750; // @[Mux.scala 46:19:@9809.4]
  wire [7:0] _T_12751; // @[Mux.scala 46:16:@9810.4]
  wire  _T_12752; // @[Mux.scala 46:19:@9811.4]
  wire [7:0] _T_12753; // @[Mux.scala 46:16:@9812.4]
  wire  _T_12754; // @[Mux.scala 46:19:@9813.4]
  wire [7:0] _T_12755; // @[Mux.scala 46:16:@9814.4]
  wire  _T_12756; // @[Mux.scala 46:19:@9815.4]
  wire [7:0] _T_12757; // @[Mux.scala 46:16:@9816.4]
  wire  _T_12758; // @[Mux.scala 46:19:@9817.4]
  wire [7:0] _T_12759; // @[Mux.scala 46:16:@9818.4]
  wire  _T_12760; // @[Mux.scala 46:19:@9819.4]
  wire [7:0] _T_12761; // @[Mux.scala 46:16:@9820.4]
  wire  _T_12792; // @[Mux.scala 46:19:@9822.4]
  wire [7:0] _T_12793; // @[Mux.scala 46:16:@9823.4]
  wire  _T_12794; // @[Mux.scala 46:19:@9824.4]
  wire [7:0] _T_12795; // @[Mux.scala 46:16:@9825.4]
  wire  _T_12796; // @[Mux.scala 46:19:@9826.4]
  wire [7:0] _T_12797; // @[Mux.scala 46:16:@9827.4]
  wire  _T_12798; // @[Mux.scala 46:19:@9828.4]
  wire [7:0] _T_12799; // @[Mux.scala 46:16:@9829.4]
  wire  _T_12800; // @[Mux.scala 46:19:@9830.4]
  wire [7:0] _T_12801; // @[Mux.scala 46:16:@9831.4]
  wire  _T_12802; // @[Mux.scala 46:19:@9832.4]
  wire [7:0] _T_12803; // @[Mux.scala 46:16:@9833.4]
  wire  _T_12804; // @[Mux.scala 46:19:@9834.4]
  wire [7:0] _T_12805; // @[Mux.scala 46:16:@9835.4]
  wire  _T_12806; // @[Mux.scala 46:19:@9836.4]
  wire [7:0] _T_12807; // @[Mux.scala 46:16:@9837.4]
  wire  _T_12808; // @[Mux.scala 46:19:@9838.4]
  wire [7:0] _T_12809; // @[Mux.scala 46:16:@9839.4]
  wire  _T_12810; // @[Mux.scala 46:19:@9840.4]
  wire [7:0] _T_12811; // @[Mux.scala 46:16:@9841.4]
  wire  _T_12812; // @[Mux.scala 46:19:@9842.4]
  wire [7:0] _T_12813; // @[Mux.scala 46:16:@9843.4]
  wire  _T_12814; // @[Mux.scala 46:19:@9844.4]
  wire [7:0] _T_12815; // @[Mux.scala 46:16:@9845.4]
  wire  _T_12816; // @[Mux.scala 46:19:@9846.4]
  wire [7:0] _T_12817; // @[Mux.scala 46:16:@9847.4]
  wire  _T_12818; // @[Mux.scala 46:19:@9848.4]
  wire [7:0] _T_12819; // @[Mux.scala 46:16:@9849.4]
  wire  _T_12820; // @[Mux.scala 46:19:@9850.4]
  wire [7:0] _T_12821; // @[Mux.scala 46:16:@9851.4]
  wire  _T_12822; // @[Mux.scala 46:19:@9852.4]
  wire [7:0] _T_12823; // @[Mux.scala 46:16:@9853.4]
  wire  _T_12824; // @[Mux.scala 46:19:@9854.4]
  wire [7:0] _T_12825; // @[Mux.scala 46:16:@9855.4]
  wire  _T_12826; // @[Mux.scala 46:19:@9856.4]
  wire [7:0] _T_12827; // @[Mux.scala 46:16:@9857.4]
  wire  _T_12828; // @[Mux.scala 46:19:@9858.4]
  wire [7:0] _T_12829; // @[Mux.scala 46:16:@9859.4]
  wire  _T_12830; // @[Mux.scala 46:19:@9860.4]
  wire [7:0] _T_12831; // @[Mux.scala 46:16:@9861.4]
  wire  _T_12832; // @[Mux.scala 46:19:@9862.4]
  wire [7:0] _T_12833; // @[Mux.scala 46:16:@9863.4]
  wire  _T_12834; // @[Mux.scala 46:19:@9864.4]
  wire [7:0] _T_12835; // @[Mux.scala 46:16:@9865.4]
  wire  _T_12836; // @[Mux.scala 46:19:@9866.4]
  wire [7:0] _T_12837; // @[Mux.scala 46:16:@9867.4]
  wire  _T_12838; // @[Mux.scala 46:19:@9868.4]
  wire [7:0] _T_12839; // @[Mux.scala 46:16:@9869.4]
  wire  _T_12840; // @[Mux.scala 46:19:@9870.4]
  wire [7:0] _T_12841; // @[Mux.scala 46:16:@9871.4]
  wire  _T_12842; // @[Mux.scala 46:19:@9872.4]
  wire [7:0] _T_12843; // @[Mux.scala 46:16:@9873.4]
  wire  _T_12844; // @[Mux.scala 46:19:@9874.4]
  wire [7:0] _T_12845; // @[Mux.scala 46:16:@9875.4]
  wire  _T_12846; // @[Mux.scala 46:19:@9876.4]
  wire [7:0] _T_12847; // @[Mux.scala 46:16:@9877.4]
  wire  _T_12848; // @[Mux.scala 46:19:@9878.4]
  wire [7:0] _T_12849; // @[Mux.scala 46:16:@9879.4]
  wire  _T_12881; // @[Mux.scala 46:19:@9881.4]
  wire [7:0] _T_12882; // @[Mux.scala 46:16:@9882.4]
  wire  _T_12883; // @[Mux.scala 46:19:@9883.4]
  wire [7:0] _T_12884; // @[Mux.scala 46:16:@9884.4]
  wire  _T_12885; // @[Mux.scala 46:19:@9885.4]
  wire [7:0] _T_12886; // @[Mux.scala 46:16:@9886.4]
  wire  _T_12887; // @[Mux.scala 46:19:@9887.4]
  wire [7:0] _T_12888; // @[Mux.scala 46:16:@9888.4]
  wire  _T_12889; // @[Mux.scala 46:19:@9889.4]
  wire [7:0] _T_12890; // @[Mux.scala 46:16:@9890.4]
  wire  _T_12891; // @[Mux.scala 46:19:@9891.4]
  wire [7:0] _T_12892; // @[Mux.scala 46:16:@9892.4]
  wire  _T_12893; // @[Mux.scala 46:19:@9893.4]
  wire [7:0] _T_12894; // @[Mux.scala 46:16:@9894.4]
  wire  _T_12895; // @[Mux.scala 46:19:@9895.4]
  wire [7:0] _T_12896; // @[Mux.scala 46:16:@9896.4]
  wire  _T_12897; // @[Mux.scala 46:19:@9897.4]
  wire [7:0] _T_12898; // @[Mux.scala 46:16:@9898.4]
  wire  _T_12899; // @[Mux.scala 46:19:@9899.4]
  wire [7:0] _T_12900; // @[Mux.scala 46:16:@9900.4]
  wire  _T_12901; // @[Mux.scala 46:19:@9901.4]
  wire [7:0] _T_12902; // @[Mux.scala 46:16:@9902.4]
  wire  _T_12903; // @[Mux.scala 46:19:@9903.4]
  wire [7:0] _T_12904; // @[Mux.scala 46:16:@9904.4]
  wire  _T_12905; // @[Mux.scala 46:19:@9905.4]
  wire [7:0] _T_12906; // @[Mux.scala 46:16:@9906.4]
  wire  _T_12907; // @[Mux.scala 46:19:@9907.4]
  wire [7:0] _T_12908; // @[Mux.scala 46:16:@9908.4]
  wire  _T_12909; // @[Mux.scala 46:19:@9909.4]
  wire [7:0] _T_12910; // @[Mux.scala 46:16:@9910.4]
  wire  _T_12911; // @[Mux.scala 46:19:@9911.4]
  wire [7:0] _T_12912; // @[Mux.scala 46:16:@9912.4]
  wire  _T_12913; // @[Mux.scala 46:19:@9913.4]
  wire [7:0] _T_12914; // @[Mux.scala 46:16:@9914.4]
  wire  _T_12915; // @[Mux.scala 46:19:@9915.4]
  wire [7:0] _T_12916; // @[Mux.scala 46:16:@9916.4]
  wire  _T_12917; // @[Mux.scala 46:19:@9917.4]
  wire [7:0] _T_12918; // @[Mux.scala 46:16:@9918.4]
  wire  _T_12919; // @[Mux.scala 46:19:@9919.4]
  wire [7:0] _T_12920; // @[Mux.scala 46:16:@9920.4]
  wire  _T_12921; // @[Mux.scala 46:19:@9921.4]
  wire [7:0] _T_12922; // @[Mux.scala 46:16:@9922.4]
  wire  _T_12923; // @[Mux.scala 46:19:@9923.4]
  wire [7:0] _T_12924; // @[Mux.scala 46:16:@9924.4]
  wire  _T_12925; // @[Mux.scala 46:19:@9925.4]
  wire [7:0] _T_12926; // @[Mux.scala 46:16:@9926.4]
  wire  _T_12927; // @[Mux.scala 46:19:@9927.4]
  wire [7:0] _T_12928; // @[Mux.scala 46:16:@9928.4]
  wire  _T_12929; // @[Mux.scala 46:19:@9929.4]
  wire [7:0] _T_12930; // @[Mux.scala 46:16:@9930.4]
  wire  _T_12931; // @[Mux.scala 46:19:@9931.4]
  wire [7:0] _T_12932; // @[Mux.scala 46:16:@9932.4]
  wire  _T_12933; // @[Mux.scala 46:19:@9933.4]
  wire [7:0] _T_12934; // @[Mux.scala 46:16:@9934.4]
  wire  _T_12935; // @[Mux.scala 46:19:@9935.4]
  wire [7:0] _T_12936; // @[Mux.scala 46:16:@9936.4]
  wire  _T_12937; // @[Mux.scala 46:19:@9937.4]
  wire [7:0] _T_12938; // @[Mux.scala 46:16:@9938.4]
  wire  _T_12939; // @[Mux.scala 46:19:@9939.4]
  wire [7:0] _T_12940; // @[Mux.scala 46:16:@9940.4]
  wire  _T_12973; // @[Mux.scala 46:19:@9942.4]
  wire [7:0] _T_12974; // @[Mux.scala 46:16:@9943.4]
  wire  _T_12975; // @[Mux.scala 46:19:@9944.4]
  wire [7:0] _T_12976; // @[Mux.scala 46:16:@9945.4]
  wire  _T_12977; // @[Mux.scala 46:19:@9946.4]
  wire [7:0] _T_12978; // @[Mux.scala 46:16:@9947.4]
  wire  _T_12979; // @[Mux.scala 46:19:@9948.4]
  wire [7:0] _T_12980; // @[Mux.scala 46:16:@9949.4]
  wire  _T_12981; // @[Mux.scala 46:19:@9950.4]
  wire [7:0] _T_12982; // @[Mux.scala 46:16:@9951.4]
  wire  _T_12983; // @[Mux.scala 46:19:@9952.4]
  wire [7:0] _T_12984; // @[Mux.scala 46:16:@9953.4]
  wire  _T_12985; // @[Mux.scala 46:19:@9954.4]
  wire [7:0] _T_12986; // @[Mux.scala 46:16:@9955.4]
  wire  _T_12987; // @[Mux.scala 46:19:@9956.4]
  wire [7:0] _T_12988; // @[Mux.scala 46:16:@9957.4]
  wire  _T_12989; // @[Mux.scala 46:19:@9958.4]
  wire [7:0] _T_12990; // @[Mux.scala 46:16:@9959.4]
  wire  _T_12991; // @[Mux.scala 46:19:@9960.4]
  wire [7:0] _T_12992; // @[Mux.scala 46:16:@9961.4]
  wire  _T_12993; // @[Mux.scala 46:19:@9962.4]
  wire [7:0] _T_12994; // @[Mux.scala 46:16:@9963.4]
  wire  _T_12995; // @[Mux.scala 46:19:@9964.4]
  wire [7:0] _T_12996; // @[Mux.scala 46:16:@9965.4]
  wire  _T_12997; // @[Mux.scala 46:19:@9966.4]
  wire [7:0] _T_12998; // @[Mux.scala 46:16:@9967.4]
  wire  _T_12999; // @[Mux.scala 46:19:@9968.4]
  wire [7:0] _T_13000; // @[Mux.scala 46:16:@9969.4]
  wire  _T_13001; // @[Mux.scala 46:19:@9970.4]
  wire [7:0] _T_13002; // @[Mux.scala 46:16:@9971.4]
  wire  _T_13003; // @[Mux.scala 46:19:@9972.4]
  wire [7:0] _T_13004; // @[Mux.scala 46:16:@9973.4]
  wire  _T_13005; // @[Mux.scala 46:19:@9974.4]
  wire [7:0] _T_13006; // @[Mux.scala 46:16:@9975.4]
  wire  _T_13007; // @[Mux.scala 46:19:@9976.4]
  wire [7:0] _T_13008; // @[Mux.scala 46:16:@9977.4]
  wire  _T_13009; // @[Mux.scala 46:19:@9978.4]
  wire [7:0] _T_13010; // @[Mux.scala 46:16:@9979.4]
  wire  _T_13011; // @[Mux.scala 46:19:@9980.4]
  wire [7:0] _T_13012; // @[Mux.scala 46:16:@9981.4]
  wire  _T_13013; // @[Mux.scala 46:19:@9982.4]
  wire [7:0] _T_13014; // @[Mux.scala 46:16:@9983.4]
  wire  _T_13015; // @[Mux.scala 46:19:@9984.4]
  wire [7:0] _T_13016; // @[Mux.scala 46:16:@9985.4]
  wire  _T_13017; // @[Mux.scala 46:19:@9986.4]
  wire [7:0] _T_13018; // @[Mux.scala 46:16:@9987.4]
  wire  _T_13019; // @[Mux.scala 46:19:@9988.4]
  wire [7:0] _T_13020; // @[Mux.scala 46:16:@9989.4]
  wire  _T_13021; // @[Mux.scala 46:19:@9990.4]
  wire [7:0] _T_13022; // @[Mux.scala 46:16:@9991.4]
  wire  _T_13023; // @[Mux.scala 46:19:@9992.4]
  wire [7:0] _T_13024; // @[Mux.scala 46:16:@9993.4]
  wire  _T_13025; // @[Mux.scala 46:19:@9994.4]
  wire [7:0] _T_13026; // @[Mux.scala 46:16:@9995.4]
  wire  _T_13027; // @[Mux.scala 46:19:@9996.4]
  wire [7:0] _T_13028; // @[Mux.scala 46:16:@9997.4]
  wire  _T_13029; // @[Mux.scala 46:19:@9998.4]
  wire [7:0] _T_13030; // @[Mux.scala 46:16:@9999.4]
  wire  _T_13031; // @[Mux.scala 46:19:@10000.4]
  wire [7:0] _T_13032; // @[Mux.scala 46:16:@10001.4]
  wire  _T_13033; // @[Mux.scala 46:19:@10002.4]
  wire [7:0] _T_13034; // @[Mux.scala 46:16:@10003.4]
  wire  _T_13068; // @[Mux.scala 46:19:@10005.4]
  wire [7:0] _T_13069; // @[Mux.scala 46:16:@10006.4]
  wire  _T_13070; // @[Mux.scala 46:19:@10007.4]
  wire [7:0] _T_13071; // @[Mux.scala 46:16:@10008.4]
  wire  _T_13072; // @[Mux.scala 46:19:@10009.4]
  wire [7:0] _T_13073; // @[Mux.scala 46:16:@10010.4]
  wire  _T_13074; // @[Mux.scala 46:19:@10011.4]
  wire [7:0] _T_13075; // @[Mux.scala 46:16:@10012.4]
  wire  _T_13076; // @[Mux.scala 46:19:@10013.4]
  wire [7:0] _T_13077; // @[Mux.scala 46:16:@10014.4]
  wire  _T_13078; // @[Mux.scala 46:19:@10015.4]
  wire [7:0] _T_13079; // @[Mux.scala 46:16:@10016.4]
  wire  _T_13080; // @[Mux.scala 46:19:@10017.4]
  wire [7:0] _T_13081; // @[Mux.scala 46:16:@10018.4]
  wire  _T_13082; // @[Mux.scala 46:19:@10019.4]
  wire [7:0] _T_13083; // @[Mux.scala 46:16:@10020.4]
  wire  _T_13084; // @[Mux.scala 46:19:@10021.4]
  wire [7:0] _T_13085; // @[Mux.scala 46:16:@10022.4]
  wire  _T_13086; // @[Mux.scala 46:19:@10023.4]
  wire [7:0] _T_13087; // @[Mux.scala 46:16:@10024.4]
  wire  _T_13088; // @[Mux.scala 46:19:@10025.4]
  wire [7:0] _T_13089; // @[Mux.scala 46:16:@10026.4]
  wire  _T_13090; // @[Mux.scala 46:19:@10027.4]
  wire [7:0] _T_13091; // @[Mux.scala 46:16:@10028.4]
  wire  _T_13092; // @[Mux.scala 46:19:@10029.4]
  wire [7:0] _T_13093; // @[Mux.scala 46:16:@10030.4]
  wire  _T_13094; // @[Mux.scala 46:19:@10031.4]
  wire [7:0] _T_13095; // @[Mux.scala 46:16:@10032.4]
  wire  _T_13096; // @[Mux.scala 46:19:@10033.4]
  wire [7:0] _T_13097; // @[Mux.scala 46:16:@10034.4]
  wire  _T_13098; // @[Mux.scala 46:19:@10035.4]
  wire [7:0] _T_13099; // @[Mux.scala 46:16:@10036.4]
  wire  _T_13100; // @[Mux.scala 46:19:@10037.4]
  wire [7:0] _T_13101; // @[Mux.scala 46:16:@10038.4]
  wire  _T_13102; // @[Mux.scala 46:19:@10039.4]
  wire [7:0] _T_13103; // @[Mux.scala 46:16:@10040.4]
  wire  _T_13104; // @[Mux.scala 46:19:@10041.4]
  wire [7:0] _T_13105; // @[Mux.scala 46:16:@10042.4]
  wire  _T_13106; // @[Mux.scala 46:19:@10043.4]
  wire [7:0] _T_13107; // @[Mux.scala 46:16:@10044.4]
  wire  _T_13108; // @[Mux.scala 46:19:@10045.4]
  wire [7:0] _T_13109; // @[Mux.scala 46:16:@10046.4]
  wire  _T_13110; // @[Mux.scala 46:19:@10047.4]
  wire [7:0] _T_13111; // @[Mux.scala 46:16:@10048.4]
  wire  _T_13112; // @[Mux.scala 46:19:@10049.4]
  wire [7:0] _T_13113; // @[Mux.scala 46:16:@10050.4]
  wire  _T_13114; // @[Mux.scala 46:19:@10051.4]
  wire [7:0] _T_13115; // @[Mux.scala 46:16:@10052.4]
  wire  _T_13116; // @[Mux.scala 46:19:@10053.4]
  wire [7:0] _T_13117; // @[Mux.scala 46:16:@10054.4]
  wire  _T_13118; // @[Mux.scala 46:19:@10055.4]
  wire [7:0] _T_13119; // @[Mux.scala 46:16:@10056.4]
  wire  _T_13120; // @[Mux.scala 46:19:@10057.4]
  wire [7:0] _T_13121; // @[Mux.scala 46:16:@10058.4]
  wire  _T_13122; // @[Mux.scala 46:19:@10059.4]
  wire [7:0] _T_13123; // @[Mux.scala 46:16:@10060.4]
  wire  _T_13124; // @[Mux.scala 46:19:@10061.4]
  wire [7:0] _T_13125; // @[Mux.scala 46:16:@10062.4]
  wire  _T_13126; // @[Mux.scala 46:19:@10063.4]
  wire [7:0] _T_13127; // @[Mux.scala 46:16:@10064.4]
  wire  _T_13128; // @[Mux.scala 46:19:@10065.4]
  wire [7:0] _T_13129; // @[Mux.scala 46:16:@10066.4]
  wire  _T_13130; // @[Mux.scala 46:19:@10067.4]
  wire [7:0] _T_13131; // @[Mux.scala 46:16:@10068.4]
  wire  _T_13166; // @[Mux.scala 46:19:@10070.4]
  wire [7:0] _T_13167; // @[Mux.scala 46:16:@10071.4]
  wire  _T_13168; // @[Mux.scala 46:19:@10072.4]
  wire [7:0] _T_13169; // @[Mux.scala 46:16:@10073.4]
  wire  _T_13170; // @[Mux.scala 46:19:@10074.4]
  wire [7:0] _T_13171; // @[Mux.scala 46:16:@10075.4]
  wire  _T_13172; // @[Mux.scala 46:19:@10076.4]
  wire [7:0] _T_13173; // @[Mux.scala 46:16:@10077.4]
  wire  _T_13174; // @[Mux.scala 46:19:@10078.4]
  wire [7:0] _T_13175; // @[Mux.scala 46:16:@10079.4]
  wire  _T_13176; // @[Mux.scala 46:19:@10080.4]
  wire [7:0] _T_13177; // @[Mux.scala 46:16:@10081.4]
  wire  _T_13178; // @[Mux.scala 46:19:@10082.4]
  wire [7:0] _T_13179; // @[Mux.scala 46:16:@10083.4]
  wire  _T_13180; // @[Mux.scala 46:19:@10084.4]
  wire [7:0] _T_13181; // @[Mux.scala 46:16:@10085.4]
  wire  _T_13182; // @[Mux.scala 46:19:@10086.4]
  wire [7:0] _T_13183; // @[Mux.scala 46:16:@10087.4]
  wire  _T_13184; // @[Mux.scala 46:19:@10088.4]
  wire [7:0] _T_13185; // @[Mux.scala 46:16:@10089.4]
  wire  _T_13186; // @[Mux.scala 46:19:@10090.4]
  wire [7:0] _T_13187; // @[Mux.scala 46:16:@10091.4]
  wire  _T_13188; // @[Mux.scala 46:19:@10092.4]
  wire [7:0] _T_13189; // @[Mux.scala 46:16:@10093.4]
  wire  _T_13190; // @[Mux.scala 46:19:@10094.4]
  wire [7:0] _T_13191; // @[Mux.scala 46:16:@10095.4]
  wire  _T_13192; // @[Mux.scala 46:19:@10096.4]
  wire [7:0] _T_13193; // @[Mux.scala 46:16:@10097.4]
  wire  _T_13194; // @[Mux.scala 46:19:@10098.4]
  wire [7:0] _T_13195; // @[Mux.scala 46:16:@10099.4]
  wire  _T_13196; // @[Mux.scala 46:19:@10100.4]
  wire [7:0] _T_13197; // @[Mux.scala 46:16:@10101.4]
  wire  _T_13198; // @[Mux.scala 46:19:@10102.4]
  wire [7:0] _T_13199; // @[Mux.scala 46:16:@10103.4]
  wire  _T_13200; // @[Mux.scala 46:19:@10104.4]
  wire [7:0] _T_13201; // @[Mux.scala 46:16:@10105.4]
  wire  _T_13202; // @[Mux.scala 46:19:@10106.4]
  wire [7:0] _T_13203; // @[Mux.scala 46:16:@10107.4]
  wire  _T_13204; // @[Mux.scala 46:19:@10108.4]
  wire [7:0] _T_13205; // @[Mux.scala 46:16:@10109.4]
  wire  _T_13206; // @[Mux.scala 46:19:@10110.4]
  wire [7:0] _T_13207; // @[Mux.scala 46:16:@10111.4]
  wire  _T_13208; // @[Mux.scala 46:19:@10112.4]
  wire [7:0] _T_13209; // @[Mux.scala 46:16:@10113.4]
  wire  _T_13210; // @[Mux.scala 46:19:@10114.4]
  wire [7:0] _T_13211; // @[Mux.scala 46:16:@10115.4]
  wire  _T_13212; // @[Mux.scala 46:19:@10116.4]
  wire [7:0] _T_13213; // @[Mux.scala 46:16:@10117.4]
  wire  _T_13214; // @[Mux.scala 46:19:@10118.4]
  wire [7:0] _T_13215; // @[Mux.scala 46:16:@10119.4]
  wire  _T_13216; // @[Mux.scala 46:19:@10120.4]
  wire [7:0] _T_13217; // @[Mux.scala 46:16:@10121.4]
  wire  _T_13218; // @[Mux.scala 46:19:@10122.4]
  wire [7:0] _T_13219; // @[Mux.scala 46:16:@10123.4]
  wire  _T_13220; // @[Mux.scala 46:19:@10124.4]
  wire [7:0] _T_13221; // @[Mux.scala 46:16:@10125.4]
  wire  _T_13222; // @[Mux.scala 46:19:@10126.4]
  wire [7:0] _T_13223; // @[Mux.scala 46:16:@10127.4]
  wire  _T_13224; // @[Mux.scala 46:19:@10128.4]
  wire [7:0] _T_13225; // @[Mux.scala 46:16:@10129.4]
  wire  _T_13226; // @[Mux.scala 46:19:@10130.4]
  wire [7:0] _T_13227; // @[Mux.scala 46:16:@10131.4]
  wire  _T_13228; // @[Mux.scala 46:19:@10132.4]
  wire [7:0] _T_13229; // @[Mux.scala 46:16:@10133.4]
  wire  _T_13230; // @[Mux.scala 46:19:@10134.4]
  wire [7:0] _T_13231; // @[Mux.scala 46:16:@10135.4]
  wire  _T_13267; // @[Mux.scala 46:19:@10137.4]
  wire [7:0] _T_13268; // @[Mux.scala 46:16:@10138.4]
  wire  _T_13269; // @[Mux.scala 46:19:@10139.4]
  wire [7:0] _T_13270; // @[Mux.scala 46:16:@10140.4]
  wire  _T_13271; // @[Mux.scala 46:19:@10141.4]
  wire [7:0] _T_13272; // @[Mux.scala 46:16:@10142.4]
  wire  _T_13273; // @[Mux.scala 46:19:@10143.4]
  wire [7:0] _T_13274; // @[Mux.scala 46:16:@10144.4]
  wire  _T_13275; // @[Mux.scala 46:19:@10145.4]
  wire [7:0] _T_13276; // @[Mux.scala 46:16:@10146.4]
  wire  _T_13277; // @[Mux.scala 46:19:@10147.4]
  wire [7:0] _T_13278; // @[Mux.scala 46:16:@10148.4]
  wire  _T_13279; // @[Mux.scala 46:19:@10149.4]
  wire [7:0] _T_13280; // @[Mux.scala 46:16:@10150.4]
  wire  _T_13281; // @[Mux.scala 46:19:@10151.4]
  wire [7:0] _T_13282; // @[Mux.scala 46:16:@10152.4]
  wire  _T_13283; // @[Mux.scala 46:19:@10153.4]
  wire [7:0] _T_13284; // @[Mux.scala 46:16:@10154.4]
  wire  _T_13285; // @[Mux.scala 46:19:@10155.4]
  wire [7:0] _T_13286; // @[Mux.scala 46:16:@10156.4]
  wire  _T_13287; // @[Mux.scala 46:19:@10157.4]
  wire [7:0] _T_13288; // @[Mux.scala 46:16:@10158.4]
  wire  _T_13289; // @[Mux.scala 46:19:@10159.4]
  wire [7:0] _T_13290; // @[Mux.scala 46:16:@10160.4]
  wire  _T_13291; // @[Mux.scala 46:19:@10161.4]
  wire [7:0] _T_13292; // @[Mux.scala 46:16:@10162.4]
  wire  _T_13293; // @[Mux.scala 46:19:@10163.4]
  wire [7:0] _T_13294; // @[Mux.scala 46:16:@10164.4]
  wire  _T_13295; // @[Mux.scala 46:19:@10165.4]
  wire [7:0] _T_13296; // @[Mux.scala 46:16:@10166.4]
  wire  _T_13297; // @[Mux.scala 46:19:@10167.4]
  wire [7:0] _T_13298; // @[Mux.scala 46:16:@10168.4]
  wire  _T_13299; // @[Mux.scala 46:19:@10169.4]
  wire [7:0] _T_13300; // @[Mux.scala 46:16:@10170.4]
  wire  _T_13301; // @[Mux.scala 46:19:@10171.4]
  wire [7:0] _T_13302; // @[Mux.scala 46:16:@10172.4]
  wire  _T_13303; // @[Mux.scala 46:19:@10173.4]
  wire [7:0] _T_13304; // @[Mux.scala 46:16:@10174.4]
  wire  _T_13305; // @[Mux.scala 46:19:@10175.4]
  wire [7:0] _T_13306; // @[Mux.scala 46:16:@10176.4]
  wire  _T_13307; // @[Mux.scala 46:19:@10177.4]
  wire [7:0] _T_13308; // @[Mux.scala 46:16:@10178.4]
  wire  _T_13309; // @[Mux.scala 46:19:@10179.4]
  wire [7:0] _T_13310; // @[Mux.scala 46:16:@10180.4]
  wire  _T_13311; // @[Mux.scala 46:19:@10181.4]
  wire [7:0] _T_13312; // @[Mux.scala 46:16:@10182.4]
  wire  _T_13313; // @[Mux.scala 46:19:@10183.4]
  wire [7:0] _T_13314; // @[Mux.scala 46:16:@10184.4]
  wire  _T_13315; // @[Mux.scala 46:19:@10185.4]
  wire [7:0] _T_13316; // @[Mux.scala 46:16:@10186.4]
  wire  _T_13317; // @[Mux.scala 46:19:@10187.4]
  wire [7:0] _T_13318; // @[Mux.scala 46:16:@10188.4]
  wire  _T_13319; // @[Mux.scala 46:19:@10189.4]
  wire [7:0] _T_13320; // @[Mux.scala 46:16:@10190.4]
  wire  _T_13321; // @[Mux.scala 46:19:@10191.4]
  wire [7:0] _T_13322; // @[Mux.scala 46:16:@10192.4]
  wire  _T_13323; // @[Mux.scala 46:19:@10193.4]
  wire [7:0] _T_13324; // @[Mux.scala 46:16:@10194.4]
  wire  _T_13325; // @[Mux.scala 46:19:@10195.4]
  wire [7:0] _T_13326; // @[Mux.scala 46:16:@10196.4]
  wire  _T_13327; // @[Mux.scala 46:19:@10197.4]
  wire [7:0] _T_13328; // @[Mux.scala 46:16:@10198.4]
  wire  _T_13329; // @[Mux.scala 46:19:@10199.4]
  wire [7:0] _T_13330; // @[Mux.scala 46:16:@10200.4]
  wire  _T_13331; // @[Mux.scala 46:19:@10201.4]
  wire [7:0] _T_13332; // @[Mux.scala 46:16:@10202.4]
  wire  _T_13333; // @[Mux.scala 46:19:@10203.4]
  wire [7:0] _T_13334; // @[Mux.scala 46:16:@10204.4]
  wire  _T_13371; // @[Mux.scala 46:19:@10206.4]
  wire [7:0] _T_13372; // @[Mux.scala 46:16:@10207.4]
  wire  _T_13373; // @[Mux.scala 46:19:@10208.4]
  wire [7:0] _T_13374; // @[Mux.scala 46:16:@10209.4]
  wire  _T_13375; // @[Mux.scala 46:19:@10210.4]
  wire [7:0] _T_13376; // @[Mux.scala 46:16:@10211.4]
  wire  _T_13377; // @[Mux.scala 46:19:@10212.4]
  wire [7:0] _T_13378; // @[Mux.scala 46:16:@10213.4]
  wire  _T_13379; // @[Mux.scala 46:19:@10214.4]
  wire [7:0] _T_13380; // @[Mux.scala 46:16:@10215.4]
  wire  _T_13381; // @[Mux.scala 46:19:@10216.4]
  wire [7:0] _T_13382; // @[Mux.scala 46:16:@10217.4]
  wire  _T_13383; // @[Mux.scala 46:19:@10218.4]
  wire [7:0] _T_13384; // @[Mux.scala 46:16:@10219.4]
  wire  _T_13385; // @[Mux.scala 46:19:@10220.4]
  wire [7:0] _T_13386; // @[Mux.scala 46:16:@10221.4]
  wire  _T_13387; // @[Mux.scala 46:19:@10222.4]
  wire [7:0] _T_13388; // @[Mux.scala 46:16:@10223.4]
  wire  _T_13389; // @[Mux.scala 46:19:@10224.4]
  wire [7:0] _T_13390; // @[Mux.scala 46:16:@10225.4]
  wire  _T_13391; // @[Mux.scala 46:19:@10226.4]
  wire [7:0] _T_13392; // @[Mux.scala 46:16:@10227.4]
  wire  _T_13393; // @[Mux.scala 46:19:@10228.4]
  wire [7:0] _T_13394; // @[Mux.scala 46:16:@10229.4]
  wire  _T_13395; // @[Mux.scala 46:19:@10230.4]
  wire [7:0] _T_13396; // @[Mux.scala 46:16:@10231.4]
  wire  _T_13397; // @[Mux.scala 46:19:@10232.4]
  wire [7:0] _T_13398; // @[Mux.scala 46:16:@10233.4]
  wire  _T_13399; // @[Mux.scala 46:19:@10234.4]
  wire [7:0] _T_13400; // @[Mux.scala 46:16:@10235.4]
  wire  _T_13401; // @[Mux.scala 46:19:@10236.4]
  wire [7:0] _T_13402; // @[Mux.scala 46:16:@10237.4]
  wire  _T_13403; // @[Mux.scala 46:19:@10238.4]
  wire [7:0] _T_13404; // @[Mux.scala 46:16:@10239.4]
  wire  _T_13405; // @[Mux.scala 46:19:@10240.4]
  wire [7:0] _T_13406; // @[Mux.scala 46:16:@10241.4]
  wire  _T_13407; // @[Mux.scala 46:19:@10242.4]
  wire [7:0] _T_13408; // @[Mux.scala 46:16:@10243.4]
  wire  _T_13409; // @[Mux.scala 46:19:@10244.4]
  wire [7:0] _T_13410; // @[Mux.scala 46:16:@10245.4]
  wire  _T_13411; // @[Mux.scala 46:19:@10246.4]
  wire [7:0] _T_13412; // @[Mux.scala 46:16:@10247.4]
  wire  _T_13413; // @[Mux.scala 46:19:@10248.4]
  wire [7:0] _T_13414; // @[Mux.scala 46:16:@10249.4]
  wire  _T_13415; // @[Mux.scala 46:19:@10250.4]
  wire [7:0] _T_13416; // @[Mux.scala 46:16:@10251.4]
  wire  _T_13417; // @[Mux.scala 46:19:@10252.4]
  wire [7:0] _T_13418; // @[Mux.scala 46:16:@10253.4]
  wire  _T_13419; // @[Mux.scala 46:19:@10254.4]
  wire [7:0] _T_13420; // @[Mux.scala 46:16:@10255.4]
  wire  _T_13421; // @[Mux.scala 46:19:@10256.4]
  wire [7:0] _T_13422; // @[Mux.scala 46:16:@10257.4]
  wire  _T_13423; // @[Mux.scala 46:19:@10258.4]
  wire [7:0] _T_13424; // @[Mux.scala 46:16:@10259.4]
  wire  _T_13425; // @[Mux.scala 46:19:@10260.4]
  wire [7:0] _T_13426; // @[Mux.scala 46:16:@10261.4]
  wire  _T_13427; // @[Mux.scala 46:19:@10262.4]
  wire [7:0] _T_13428; // @[Mux.scala 46:16:@10263.4]
  wire  _T_13429; // @[Mux.scala 46:19:@10264.4]
  wire [7:0] _T_13430; // @[Mux.scala 46:16:@10265.4]
  wire  _T_13431; // @[Mux.scala 46:19:@10266.4]
  wire [7:0] _T_13432; // @[Mux.scala 46:16:@10267.4]
  wire  _T_13433; // @[Mux.scala 46:19:@10268.4]
  wire [7:0] _T_13434; // @[Mux.scala 46:16:@10269.4]
  wire  _T_13435; // @[Mux.scala 46:19:@10270.4]
  wire [7:0] _T_13436; // @[Mux.scala 46:16:@10271.4]
  wire  _T_13437; // @[Mux.scala 46:19:@10272.4]
  wire [7:0] _T_13438; // @[Mux.scala 46:16:@10273.4]
  wire  _T_13439; // @[Mux.scala 46:19:@10274.4]
  wire [7:0] _T_13440; // @[Mux.scala 46:16:@10275.4]
  wire  _T_13478; // @[Mux.scala 46:19:@10277.4]
  wire [7:0] _T_13479; // @[Mux.scala 46:16:@10278.4]
  wire  _T_13480; // @[Mux.scala 46:19:@10279.4]
  wire [7:0] _T_13481; // @[Mux.scala 46:16:@10280.4]
  wire  _T_13482; // @[Mux.scala 46:19:@10281.4]
  wire [7:0] _T_13483; // @[Mux.scala 46:16:@10282.4]
  wire  _T_13484; // @[Mux.scala 46:19:@10283.4]
  wire [7:0] _T_13485; // @[Mux.scala 46:16:@10284.4]
  wire  _T_13486; // @[Mux.scala 46:19:@10285.4]
  wire [7:0] _T_13487; // @[Mux.scala 46:16:@10286.4]
  wire  _T_13488; // @[Mux.scala 46:19:@10287.4]
  wire [7:0] _T_13489; // @[Mux.scala 46:16:@10288.4]
  wire  _T_13490; // @[Mux.scala 46:19:@10289.4]
  wire [7:0] _T_13491; // @[Mux.scala 46:16:@10290.4]
  wire  _T_13492; // @[Mux.scala 46:19:@10291.4]
  wire [7:0] _T_13493; // @[Mux.scala 46:16:@10292.4]
  wire  _T_13494; // @[Mux.scala 46:19:@10293.4]
  wire [7:0] _T_13495; // @[Mux.scala 46:16:@10294.4]
  wire  _T_13496; // @[Mux.scala 46:19:@10295.4]
  wire [7:0] _T_13497; // @[Mux.scala 46:16:@10296.4]
  wire  _T_13498; // @[Mux.scala 46:19:@10297.4]
  wire [7:0] _T_13499; // @[Mux.scala 46:16:@10298.4]
  wire  _T_13500; // @[Mux.scala 46:19:@10299.4]
  wire [7:0] _T_13501; // @[Mux.scala 46:16:@10300.4]
  wire  _T_13502; // @[Mux.scala 46:19:@10301.4]
  wire [7:0] _T_13503; // @[Mux.scala 46:16:@10302.4]
  wire  _T_13504; // @[Mux.scala 46:19:@10303.4]
  wire [7:0] _T_13505; // @[Mux.scala 46:16:@10304.4]
  wire  _T_13506; // @[Mux.scala 46:19:@10305.4]
  wire [7:0] _T_13507; // @[Mux.scala 46:16:@10306.4]
  wire  _T_13508; // @[Mux.scala 46:19:@10307.4]
  wire [7:0] _T_13509; // @[Mux.scala 46:16:@10308.4]
  wire  _T_13510; // @[Mux.scala 46:19:@10309.4]
  wire [7:0] _T_13511; // @[Mux.scala 46:16:@10310.4]
  wire  _T_13512; // @[Mux.scala 46:19:@10311.4]
  wire [7:0] _T_13513; // @[Mux.scala 46:16:@10312.4]
  wire  _T_13514; // @[Mux.scala 46:19:@10313.4]
  wire [7:0] _T_13515; // @[Mux.scala 46:16:@10314.4]
  wire  _T_13516; // @[Mux.scala 46:19:@10315.4]
  wire [7:0] _T_13517; // @[Mux.scala 46:16:@10316.4]
  wire  _T_13518; // @[Mux.scala 46:19:@10317.4]
  wire [7:0] _T_13519; // @[Mux.scala 46:16:@10318.4]
  wire  _T_13520; // @[Mux.scala 46:19:@10319.4]
  wire [7:0] _T_13521; // @[Mux.scala 46:16:@10320.4]
  wire  _T_13522; // @[Mux.scala 46:19:@10321.4]
  wire [7:0] _T_13523; // @[Mux.scala 46:16:@10322.4]
  wire  _T_13524; // @[Mux.scala 46:19:@10323.4]
  wire [7:0] _T_13525; // @[Mux.scala 46:16:@10324.4]
  wire  _T_13526; // @[Mux.scala 46:19:@10325.4]
  wire [7:0] _T_13527; // @[Mux.scala 46:16:@10326.4]
  wire  _T_13528; // @[Mux.scala 46:19:@10327.4]
  wire [7:0] _T_13529; // @[Mux.scala 46:16:@10328.4]
  wire  _T_13530; // @[Mux.scala 46:19:@10329.4]
  wire [7:0] _T_13531; // @[Mux.scala 46:16:@10330.4]
  wire  _T_13532; // @[Mux.scala 46:19:@10331.4]
  wire [7:0] _T_13533; // @[Mux.scala 46:16:@10332.4]
  wire  _T_13534; // @[Mux.scala 46:19:@10333.4]
  wire [7:0] _T_13535; // @[Mux.scala 46:16:@10334.4]
  wire  _T_13536; // @[Mux.scala 46:19:@10335.4]
  wire [7:0] _T_13537; // @[Mux.scala 46:16:@10336.4]
  wire  _T_13538; // @[Mux.scala 46:19:@10337.4]
  wire [7:0] _T_13539; // @[Mux.scala 46:16:@10338.4]
  wire  _T_13540; // @[Mux.scala 46:19:@10339.4]
  wire [7:0] _T_13541; // @[Mux.scala 46:16:@10340.4]
  wire  _T_13542; // @[Mux.scala 46:19:@10341.4]
  wire [7:0] _T_13543; // @[Mux.scala 46:16:@10342.4]
  wire  _T_13544; // @[Mux.scala 46:19:@10343.4]
  wire [7:0] _T_13545; // @[Mux.scala 46:16:@10344.4]
  wire  _T_13546; // @[Mux.scala 46:19:@10345.4]
  wire [7:0] _T_13547; // @[Mux.scala 46:16:@10346.4]
  wire  _T_13548; // @[Mux.scala 46:19:@10347.4]
  wire [7:0] _T_13549; // @[Mux.scala 46:16:@10348.4]
  wire  _T_13588; // @[Mux.scala 46:19:@10350.4]
  wire [7:0] _T_13589; // @[Mux.scala 46:16:@10351.4]
  wire  _T_13590; // @[Mux.scala 46:19:@10352.4]
  wire [7:0] _T_13591; // @[Mux.scala 46:16:@10353.4]
  wire  _T_13592; // @[Mux.scala 46:19:@10354.4]
  wire [7:0] _T_13593; // @[Mux.scala 46:16:@10355.4]
  wire  _T_13594; // @[Mux.scala 46:19:@10356.4]
  wire [7:0] _T_13595; // @[Mux.scala 46:16:@10357.4]
  wire  _T_13596; // @[Mux.scala 46:19:@10358.4]
  wire [7:0] _T_13597; // @[Mux.scala 46:16:@10359.4]
  wire  _T_13598; // @[Mux.scala 46:19:@10360.4]
  wire [7:0] _T_13599; // @[Mux.scala 46:16:@10361.4]
  wire  _T_13600; // @[Mux.scala 46:19:@10362.4]
  wire [7:0] _T_13601; // @[Mux.scala 46:16:@10363.4]
  wire  _T_13602; // @[Mux.scala 46:19:@10364.4]
  wire [7:0] _T_13603; // @[Mux.scala 46:16:@10365.4]
  wire  _T_13604; // @[Mux.scala 46:19:@10366.4]
  wire [7:0] _T_13605; // @[Mux.scala 46:16:@10367.4]
  wire  _T_13606; // @[Mux.scala 46:19:@10368.4]
  wire [7:0] _T_13607; // @[Mux.scala 46:16:@10369.4]
  wire  _T_13608; // @[Mux.scala 46:19:@10370.4]
  wire [7:0] _T_13609; // @[Mux.scala 46:16:@10371.4]
  wire  _T_13610; // @[Mux.scala 46:19:@10372.4]
  wire [7:0] _T_13611; // @[Mux.scala 46:16:@10373.4]
  wire  _T_13612; // @[Mux.scala 46:19:@10374.4]
  wire [7:0] _T_13613; // @[Mux.scala 46:16:@10375.4]
  wire  _T_13614; // @[Mux.scala 46:19:@10376.4]
  wire [7:0] _T_13615; // @[Mux.scala 46:16:@10377.4]
  wire  _T_13616; // @[Mux.scala 46:19:@10378.4]
  wire [7:0] _T_13617; // @[Mux.scala 46:16:@10379.4]
  wire  _T_13618; // @[Mux.scala 46:19:@10380.4]
  wire [7:0] _T_13619; // @[Mux.scala 46:16:@10381.4]
  wire  _T_13620; // @[Mux.scala 46:19:@10382.4]
  wire [7:0] _T_13621; // @[Mux.scala 46:16:@10383.4]
  wire  _T_13622; // @[Mux.scala 46:19:@10384.4]
  wire [7:0] _T_13623; // @[Mux.scala 46:16:@10385.4]
  wire  _T_13624; // @[Mux.scala 46:19:@10386.4]
  wire [7:0] _T_13625; // @[Mux.scala 46:16:@10387.4]
  wire  _T_13626; // @[Mux.scala 46:19:@10388.4]
  wire [7:0] _T_13627; // @[Mux.scala 46:16:@10389.4]
  wire  _T_13628; // @[Mux.scala 46:19:@10390.4]
  wire [7:0] _T_13629; // @[Mux.scala 46:16:@10391.4]
  wire  _T_13630; // @[Mux.scala 46:19:@10392.4]
  wire [7:0] _T_13631; // @[Mux.scala 46:16:@10393.4]
  wire  _T_13632; // @[Mux.scala 46:19:@10394.4]
  wire [7:0] _T_13633; // @[Mux.scala 46:16:@10395.4]
  wire  _T_13634; // @[Mux.scala 46:19:@10396.4]
  wire [7:0] _T_13635; // @[Mux.scala 46:16:@10397.4]
  wire  _T_13636; // @[Mux.scala 46:19:@10398.4]
  wire [7:0] _T_13637; // @[Mux.scala 46:16:@10399.4]
  wire  _T_13638; // @[Mux.scala 46:19:@10400.4]
  wire [7:0] _T_13639; // @[Mux.scala 46:16:@10401.4]
  wire  _T_13640; // @[Mux.scala 46:19:@10402.4]
  wire [7:0] _T_13641; // @[Mux.scala 46:16:@10403.4]
  wire  _T_13642; // @[Mux.scala 46:19:@10404.4]
  wire [7:0] _T_13643; // @[Mux.scala 46:16:@10405.4]
  wire  _T_13644; // @[Mux.scala 46:19:@10406.4]
  wire [7:0] _T_13645; // @[Mux.scala 46:16:@10407.4]
  wire  _T_13646; // @[Mux.scala 46:19:@10408.4]
  wire [7:0] _T_13647; // @[Mux.scala 46:16:@10409.4]
  wire  _T_13648; // @[Mux.scala 46:19:@10410.4]
  wire [7:0] _T_13649; // @[Mux.scala 46:16:@10411.4]
  wire  _T_13650; // @[Mux.scala 46:19:@10412.4]
  wire [7:0] _T_13651; // @[Mux.scala 46:16:@10413.4]
  wire  _T_13652; // @[Mux.scala 46:19:@10414.4]
  wire [7:0] _T_13653; // @[Mux.scala 46:16:@10415.4]
  wire  _T_13654; // @[Mux.scala 46:19:@10416.4]
  wire [7:0] _T_13655; // @[Mux.scala 46:16:@10417.4]
  wire  _T_13656; // @[Mux.scala 46:19:@10418.4]
  wire [7:0] _T_13657; // @[Mux.scala 46:16:@10419.4]
  wire  _T_13658; // @[Mux.scala 46:19:@10420.4]
  wire [7:0] _T_13659; // @[Mux.scala 46:16:@10421.4]
  wire  _T_13660; // @[Mux.scala 46:19:@10422.4]
  wire [7:0] _T_13661; // @[Mux.scala 46:16:@10423.4]
  wire  _T_13701; // @[Mux.scala 46:19:@10425.4]
  wire [7:0] _T_13702; // @[Mux.scala 46:16:@10426.4]
  wire  _T_13703; // @[Mux.scala 46:19:@10427.4]
  wire [7:0] _T_13704; // @[Mux.scala 46:16:@10428.4]
  wire  _T_13705; // @[Mux.scala 46:19:@10429.4]
  wire [7:0] _T_13706; // @[Mux.scala 46:16:@10430.4]
  wire  _T_13707; // @[Mux.scala 46:19:@10431.4]
  wire [7:0] _T_13708; // @[Mux.scala 46:16:@10432.4]
  wire  _T_13709; // @[Mux.scala 46:19:@10433.4]
  wire [7:0] _T_13710; // @[Mux.scala 46:16:@10434.4]
  wire  _T_13711; // @[Mux.scala 46:19:@10435.4]
  wire [7:0] _T_13712; // @[Mux.scala 46:16:@10436.4]
  wire  _T_13713; // @[Mux.scala 46:19:@10437.4]
  wire [7:0] _T_13714; // @[Mux.scala 46:16:@10438.4]
  wire  _T_13715; // @[Mux.scala 46:19:@10439.4]
  wire [7:0] _T_13716; // @[Mux.scala 46:16:@10440.4]
  wire  _T_13717; // @[Mux.scala 46:19:@10441.4]
  wire [7:0] _T_13718; // @[Mux.scala 46:16:@10442.4]
  wire  _T_13719; // @[Mux.scala 46:19:@10443.4]
  wire [7:0] _T_13720; // @[Mux.scala 46:16:@10444.4]
  wire  _T_13721; // @[Mux.scala 46:19:@10445.4]
  wire [7:0] _T_13722; // @[Mux.scala 46:16:@10446.4]
  wire  _T_13723; // @[Mux.scala 46:19:@10447.4]
  wire [7:0] _T_13724; // @[Mux.scala 46:16:@10448.4]
  wire  _T_13725; // @[Mux.scala 46:19:@10449.4]
  wire [7:0] _T_13726; // @[Mux.scala 46:16:@10450.4]
  wire  _T_13727; // @[Mux.scala 46:19:@10451.4]
  wire [7:0] _T_13728; // @[Mux.scala 46:16:@10452.4]
  wire  _T_13729; // @[Mux.scala 46:19:@10453.4]
  wire [7:0] _T_13730; // @[Mux.scala 46:16:@10454.4]
  wire  _T_13731; // @[Mux.scala 46:19:@10455.4]
  wire [7:0] _T_13732; // @[Mux.scala 46:16:@10456.4]
  wire  _T_13733; // @[Mux.scala 46:19:@10457.4]
  wire [7:0] _T_13734; // @[Mux.scala 46:16:@10458.4]
  wire  _T_13735; // @[Mux.scala 46:19:@10459.4]
  wire [7:0] _T_13736; // @[Mux.scala 46:16:@10460.4]
  wire  _T_13737; // @[Mux.scala 46:19:@10461.4]
  wire [7:0] _T_13738; // @[Mux.scala 46:16:@10462.4]
  wire  _T_13739; // @[Mux.scala 46:19:@10463.4]
  wire [7:0] _T_13740; // @[Mux.scala 46:16:@10464.4]
  wire  _T_13741; // @[Mux.scala 46:19:@10465.4]
  wire [7:0] _T_13742; // @[Mux.scala 46:16:@10466.4]
  wire  _T_13743; // @[Mux.scala 46:19:@10467.4]
  wire [7:0] _T_13744; // @[Mux.scala 46:16:@10468.4]
  wire  _T_13745; // @[Mux.scala 46:19:@10469.4]
  wire [7:0] _T_13746; // @[Mux.scala 46:16:@10470.4]
  wire  _T_13747; // @[Mux.scala 46:19:@10471.4]
  wire [7:0] _T_13748; // @[Mux.scala 46:16:@10472.4]
  wire  _T_13749; // @[Mux.scala 46:19:@10473.4]
  wire [7:0] _T_13750; // @[Mux.scala 46:16:@10474.4]
  wire  _T_13751; // @[Mux.scala 46:19:@10475.4]
  wire [7:0] _T_13752; // @[Mux.scala 46:16:@10476.4]
  wire  _T_13753; // @[Mux.scala 46:19:@10477.4]
  wire [7:0] _T_13754; // @[Mux.scala 46:16:@10478.4]
  wire  _T_13755; // @[Mux.scala 46:19:@10479.4]
  wire [7:0] _T_13756; // @[Mux.scala 46:16:@10480.4]
  wire  _T_13757; // @[Mux.scala 46:19:@10481.4]
  wire [7:0] _T_13758; // @[Mux.scala 46:16:@10482.4]
  wire  _T_13759; // @[Mux.scala 46:19:@10483.4]
  wire [7:0] _T_13760; // @[Mux.scala 46:16:@10484.4]
  wire  _T_13761; // @[Mux.scala 46:19:@10485.4]
  wire [7:0] _T_13762; // @[Mux.scala 46:16:@10486.4]
  wire  _T_13763; // @[Mux.scala 46:19:@10487.4]
  wire [7:0] _T_13764; // @[Mux.scala 46:16:@10488.4]
  wire  _T_13765; // @[Mux.scala 46:19:@10489.4]
  wire [7:0] _T_13766; // @[Mux.scala 46:16:@10490.4]
  wire  _T_13767; // @[Mux.scala 46:19:@10491.4]
  wire [7:0] _T_13768; // @[Mux.scala 46:16:@10492.4]
  wire  _T_13769; // @[Mux.scala 46:19:@10493.4]
  wire [7:0] _T_13770; // @[Mux.scala 46:16:@10494.4]
  wire  _T_13771; // @[Mux.scala 46:19:@10495.4]
  wire [7:0] _T_13772; // @[Mux.scala 46:16:@10496.4]
  wire  _T_13773; // @[Mux.scala 46:19:@10497.4]
  wire [7:0] _T_13774; // @[Mux.scala 46:16:@10498.4]
  wire  _T_13775; // @[Mux.scala 46:19:@10499.4]
  wire [7:0] _T_13776; // @[Mux.scala 46:16:@10500.4]
  wire  _T_13817; // @[Mux.scala 46:19:@10502.4]
  wire [7:0] _T_13818; // @[Mux.scala 46:16:@10503.4]
  wire  _T_13819; // @[Mux.scala 46:19:@10504.4]
  wire [7:0] _T_13820; // @[Mux.scala 46:16:@10505.4]
  wire  _T_13821; // @[Mux.scala 46:19:@10506.4]
  wire [7:0] _T_13822; // @[Mux.scala 46:16:@10507.4]
  wire  _T_13823; // @[Mux.scala 46:19:@10508.4]
  wire [7:0] _T_13824; // @[Mux.scala 46:16:@10509.4]
  wire  _T_13825; // @[Mux.scala 46:19:@10510.4]
  wire [7:0] _T_13826; // @[Mux.scala 46:16:@10511.4]
  wire  _T_13827; // @[Mux.scala 46:19:@10512.4]
  wire [7:0] _T_13828; // @[Mux.scala 46:16:@10513.4]
  wire  _T_13829; // @[Mux.scala 46:19:@10514.4]
  wire [7:0] _T_13830; // @[Mux.scala 46:16:@10515.4]
  wire  _T_13831; // @[Mux.scala 46:19:@10516.4]
  wire [7:0] _T_13832; // @[Mux.scala 46:16:@10517.4]
  wire  _T_13833; // @[Mux.scala 46:19:@10518.4]
  wire [7:0] _T_13834; // @[Mux.scala 46:16:@10519.4]
  wire  _T_13835; // @[Mux.scala 46:19:@10520.4]
  wire [7:0] _T_13836; // @[Mux.scala 46:16:@10521.4]
  wire  _T_13837; // @[Mux.scala 46:19:@10522.4]
  wire [7:0] _T_13838; // @[Mux.scala 46:16:@10523.4]
  wire  _T_13839; // @[Mux.scala 46:19:@10524.4]
  wire [7:0] _T_13840; // @[Mux.scala 46:16:@10525.4]
  wire  _T_13841; // @[Mux.scala 46:19:@10526.4]
  wire [7:0] _T_13842; // @[Mux.scala 46:16:@10527.4]
  wire  _T_13843; // @[Mux.scala 46:19:@10528.4]
  wire [7:0] _T_13844; // @[Mux.scala 46:16:@10529.4]
  wire  _T_13845; // @[Mux.scala 46:19:@10530.4]
  wire [7:0] _T_13846; // @[Mux.scala 46:16:@10531.4]
  wire  _T_13847; // @[Mux.scala 46:19:@10532.4]
  wire [7:0] _T_13848; // @[Mux.scala 46:16:@10533.4]
  wire  _T_13849; // @[Mux.scala 46:19:@10534.4]
  wire [7:0] _T_13850; // @[Mux.scala 46:16:@10535.4]
  wire  _T_13851; // @[Mux.scala 46:19:@10536.4]
  wire [7:0] _T_13852; // @[Mux.scala 46:16:@10537.4]
  wire  _T_13853; // @[Mux.scala 46:19:@10538.4]
  wire [7:0] _T_13854; // @[Mux.scala 46:16:@10539.4]
  wire  _T_13855; // @[Mux.scala 46:19:@10540.4]
  wire [7:0] _T_13856; // @[Mux.scala 46:16:@10541.4]
  wire  _T_13857; // @[Mux.scala 46:19:@10542.4]
  wire [7:0] _T_13858; // @[Mux.scala 46:16:@10543.4]
  wire  _T_13859; // @[Mux.scala 46:19:@10544.4]
  wire [7:0] _T_13860; // @[Mux.scala 46:16:@10545.4]
  wire  _T_13861; // @[Mux.scala 46:19:@10546.4]
  wire [7:0] _T_13862; // @[Mux.scala 46:16:@10547.4]
  wire  _T_13863; // @[Mux.scala 46:19:@10548.4]
  wire [7:0] _T_13864; // @[Mux.scala 46:16:@10549.4]
  wire  _T_13865; // @[Mux.scala 46:19:@10550.4]
  wire [7:0] _T_13866; // @[Mux.scala 46:16:@10551.4]
  wire  _T_13867; // @[Mux.scala 46:19:@10552.4]
  wire [7:0] _T_13868; // @[Mux.scala 46:16:@10553.4]
  wire  _T_13869; // @[Mux.scala 46:19:@10554.4]
  wire [7:0] _T_13870; // @[Mux.scala 46:16:@10555.4]
  wire  _T_13871; // @[Mux.scala 46:19:@10556.4]
  wire [7:0] _T_13872; // @[Mux.scala 46:16:@10557.4]
  wire  _T_13873; // @[Mux.scala 46:19:@10558.4]
  wire [7:0] _T_13874; // @[Mux.scala 46:16:@10559.4]
  wire  _T_13875; // @[Mux.scala 46:19:@10560.4]
  wire [7:0] _T_13876; // @[Mux.scala 46:16:@10561.4]
  wire  _T_13877; // @[Mux.scala 46:19:@10562.4]
  wire [7:0] _T_13878; // @[Mux.scala 46:16:@10563.4]
  wire  _T_13879; // @[Mux.scala 46:19:@10564.4]
  wire [7:0] _T_13880; // @[Mux.scala 46:16:@10565.4]
  wire  _T_13881; // @[Mux.scala 46:19:@10566.4]
  wire [7:0] _T_13882; // @[Mux.scala 46:16:@10567.4]
  wire  _T_13883; // @[Mux.scala 46:19:@10568.4]
  wire [7:0] _T_13884; // @[Mux.scala 46:16:@10569.4]
  wire  _T_13885; // @[Mux.scala 46:19:@10570.4]
  wire [7:0] _T_13886; // @[Mux.scala 46:16:@10571.4]
  wire  _T_13887; // @[Mux.scala 46:19:@10572.4]
  wire [7:0] _T_13888; // @[Mux.scala 46:16:@10573.4]
  wire  _T_13889; // @[Mux.scala 46:19:@10574.4]
  wire [7:0] _T_13890; // @[Mux.scala 46:16:@10575.4]
  wire  _T_13891; // @[Mux.scala 46:19:@10576.4]
  wire [7:0] _T_13892; // @[Mux.scala 46:16:@10577.4]
  wire  _T_13893; // @[Mux.scala 46:19:@10578.4]
  wire [7:0] _T_13894; // @[Mux.scala 46:16:@10579.4]
  wire  _T_13936; // @[Mux.scala 46:19:@10581.4]
  wire [7:0] _T_13937; // @[Mux.scala 46:16:@10582.4]
  wire  _T_13938; // @[Mux.scala 46:19:@10583.4]
  wire [7:0] _T_13939; // @[Mux.scala 46:16:@10584.4]
  wire  _T_13940; // @[Mux.scala 46:19:@10585.4]
  wire [7:0] _T_13941; // @[Mux.scala 46:16:@10586.4]
  wire  _T_13942; // @[Mux.scala 46:19:@10587.4]
  wire [7:0] _T_13943; // @[Mux.scala 46:16:@10588.4]
  wire  _T_13944; // @[Mux.scala 46:19:@10589.4]
  wire [7:0] _T_13945; // @[Mux.scala 46:16:@10590.4]
  wire  _T_13946; // @[Mux.scala 46:19:@10591.4]
  wire [7:0] _T_13947; // @[Mux.scala 46:16:@10592.4]
  wire  _T_13948; // @[Mux.scala 46:19:@10593.4]
  wire [7:0] _T_13949; // @[Mux.scala 46:16:@10594.4]
  wire  _T_13950; // @[Mux.scala 46:19:@10595.4]
  wire [7:0] _T_13951; // @[Mux.scala 46:16:@10596.4]
  wire  _T_13952; // @[Mux.scala 46:19:@10597.4]
  wire [7:0] _T_13953; // @[Mux.scala 46:16:@10598.4]
  wire  _T_13954; // @[Mux.scala 46:19:@10599.4]
  wire [7:0] _T_13955; // @[Mux.scala 46:16:@10600.4]
  wire  _T_13956; // @[Mux.scala 46:19:@10601.4]
  wire [7:0] _T_13957; // @[Mux.scala 46:16:@10602.4]
  wire  _T_13958; // @[Mux.scala 46:19:@10603.4]
  wire [7:0] _T_13959; // @[Mux.scala 46:16:@10604.4]
  wire  _T_13960; // @[Mux.scala 46:19:@10605.4]
  wire [7:0] _T_13961; // @[Mux.scala 46:16:@10606.4]
  wire  _T_13962; // @[Mux.scala 46:19:@10607.4]
  wire [7:0] _T_13963; // @[Mux.scala 46:16:@10608.4]
  wire  _T_13964; // @[Mux.scala 46:19:@10609.4]
  wire [7:0] _T_13965; // @[Mux.scala 46:16:@10610.4]
  wire  _T_13966; // @[Mux.scala 46:19:@10611.4]
  wire [7:0] _T_13967; // @[Mux.scala 46:16:@10612.4]
  wire  _T_13968; // @[Mux.scala 46:19:@10613.4]
  wire [7:0] _T_13969; // @[Mux.scala 46:16:@10614.4]
  wire  _T_13970; // @[Mux.scala 46:19:@10615.4]
  wire [7:0] _T_13971; // @[Mux.scala 46:16:@10616.4]
  wire  _T_13972; // @[Mux.scala 46:19:@10617.4]
  wire [7:0] _T_13973; // @[Mux.scala 46:16:@10618.4]
  wire  _T_13974; // @[Mux.scala 46:19:@10619.4]
  wire [7:0] _T_13975; // @[Mux.scala 46:16:@10620.4]
  wire  _T_13976; // @[Mux.scala 46:19:@10621.4]
  wire [7:0] _T_13977; // @[Mux.scala 46:16:@10622.4]
  wire  _T_13978; // @[Mux.scala 46:19:@10623.4]
  wire [7:0] _T_13979; // @[Mux.scala 46:16:@10624.4]
  wire  _T_13980; // @[Mux.scala 46:19:@10625.4]
  wire [7:0] _T_13981; // @[Mux.scala 46:16:@10626.4]
  wire  _T_13982; // @[Mux.scala 46:19:@10627.4]
  wire [7:0] _T_13983; // @[Mux.scala 46:16:@10628.4]
  wire  _T_13984; // @[Mux.scala 46:19:@10629.4]
  wire [7:0] _T_13985; // @[Mux.scala 46:16:@10630.4]
  wire  _T_13986; // @[Mux.scala 46:19:@10631.4]
  wire [7:0] _T_13987; // @[Mux.scala 46:16:@10632.4]
  wire  _T_13988; // @[Mux.scala 46:19:@10633.4]
  wire [7:0] _T_13989; // @[Mux.scala 46:16:@10634.4]
  wire  _T_13990; // @[Mux.scala 46:19:@10635.4]
  wire [7:0] _T_13991; // @[Mux.scala 46:16:@10636.4]
  wire  _T_13992; // @[Mux.scala 46:19:@10637.4]
  wire [7:0] _T_13993; // @[Mux.scala 46:16:@10638.4]
  wire  _T_13994; // @[Mux.scala 46:19:@10639.4]
  wire [7:0] _T_13995; // @[Mux.scala 46:16:@10640.4]
  wire  _T_13996; // @[Mux.scala 46:19:@10641.4]
  wire [7:0] _T_13997; // @[Mux.scala 46:16:@10642.4]
  wire  _T_13998; // @[Mux.scala 46:19:@10643.4]
  wire [7:0] _T_13999; // @[Mux.scala 46:16:@10644.4]
  wire  _T_14000; // @[Mux.scala 46:19:@10645.4]
  wire [7:0] _T_14001; // @[Mux.scala 46:16:@10646.4]
  wire  _T_14002; // @[Mux.scala 46:19:@10647.4]
  wire [7:0] _T_14003; // @[Mux.scala 46:16:@10648.4]
  wire  _T_14004; // @[Mux.scala 46:19:@10649.4]
  wire [7:0] _T_14005; // @[Mux.scala 46:16:@10650.4]
  wire  _T_14006; // @[Mux.scala 46:19:@10651.4]
  wire [7:0] _T_14007; // @[Mux.scala 46:16:@10652.4]
  wire  _T_14008; // @[Mux.scala 46:19:@10653.4]
  wire [7:0] _T_14009; // @[Mux.scala 46:16:@10654.4]
  wire  _T_14010; // @[Mux.scala 46:19:@10655.4]
  wire [7:0] _T_14011; // @[Mux.scala 46:16:@10656.4]
  wire  _T_14012; // @[Mux.scala 46:19:@10657.4]
  wire [7:0] _T_14013; // @[Mux.scala 46:16:@10658.4]
  wire  _T_14014; // @[Mux.scala 46:19:@10659.4]
  wire [7:0] _T_14015; // @[Mux.scala 46:16:@10660.4]
  wire  _T_14058; // @[Mux.scala 46:19:@10662.4]
  wire [7:0] _T_14059; // @[Mux.scala 46:16:@10663.4]
  wire  _T_14060; // @[Mux.scala 46:19:@10664.4]
  wire [7:0] _T_14061; // @[Mux.scala 46:16:@10665.4]
  wire  _T_14062; // @[Mux.scala 46:19:@10666.4]
  wire [7:0] _T_14063; // @[Mux.scala 46:16:@10667.4]
  wire  _T_14064; // @[Mux.scala 46:19:@10668.4]
  wire [7:0] _T_14065; // @[Mux.scala 46:16:@10669.4]
  wire  _T_14066; // @[Mux.scala 46:19:@10670.4]
  wire [7:0] _T_14067; // @[Mux.scala 46:16:@10671.4]
  wire  _T_14068; // @[Mux.scala 46:19:@10672.4]
  wire [7:0] _T_14069; // @[Mux.scala 46:16:@10673.4]
  wire  _T_14070; // @[Mux.scala 46:19:@10674.4]
  wire [7:0] _T_14071; // @[Mux.scala 46:16:@10675.4]
  wire  _T_14072; // @[Mux.scala 46:19:@10676.4]
  wire [7:0] _T_14073; // @[Mux.scala 46:16:@10677.4]
  wire  _T_14074; // @[Mux.scala 46:19:@10678.4]
  wire [7:0] _T_14075; // @[Mux.scala 46:16:@10679.4]
  wire  _T_14076; // @[Mux.scala 46:19:@10680.4]
  wire [7:0] _T_14077; // @[Mux.scala 46:16:@10681.4]
  wire  _T_14078; // @[Mux.scala 46:19:@10682.4]
  wire [7:0] _T_14079; // @[Mux.scala 46:16:@10683.4]
  wire  _T_14080; // @[Mux.scala 46:19:@10684.4]
  wire [7:0] _T_14081; // @[Mux.scala 46:16:@10685.4]
  wire  _T_14082; // @[Mux.scala 46:19:@10686.4]
  wire [7:0] _T_14083; // @[Mux.scala 46:16:@10687.4]
  wire  _T_14084; // @[Mux.scala 46:19:@10688.4]
  wire [7:0] _T_14085; // @[Mux.scala 46:16:@10689.4]
  wire  _T_14086; // @[Mux.scala 46:19:@10690.4]
  wire [7:0] _T_14087; // @[Mux.scala 46:16:@10691.4]
  wire  _T_14088; // @[Mux.scala 46:19:@10692.4]
  wire [7:0] _T_14089; // @[Mux.scala 46:16:@10693.4]
  wire  _T_14090; // @[Mux.scala 46:19:@10694.4]
  wire [7:0] _T_14091; // @[Mux.scala 46:16:@10695.4]
  wire  _T_14092; // @[Mux.scala 46:19:@10696.4]
  wire [7:0] _T_14093; // @[Mux.scala 46:16:@10697.4]
  wire  _T_14094; // @[Mux.scala 46:19:@10698.4]
  wire [7:0] _T_14095; // @[Mux.scala 46:16:@10699.4]
  wire  _T_14096; // @[Mux.scala 46:19:@10700.4]
  wire [7:0] _T_14097; // @[Mux.scala 46:16:@10701.4]
  wire  _T_14098; // @[Mux.scala 46:19:@10702.4]
  wire [7:0] _T_14099; // @[Mux.scala 46:16:@10703.4]
  wire  _T_14100; // @[Mux.scala 46:19:@10704.4]
  wire [7:0] _T_14101; // @[Mux.scala 46:16:@10705.4]
  wire  _T_14102; // @[Mux.scala 46:19:@10706.4]
  wire [7:0] _T_14103; // @[Mux.scala 46:16:@10707.4]
  wire  _T_14104; // @[Mux.scala 46:19:@10708.4]
  wire [7:0] _T_14105; // @[Mux.scala 46:16:@10709.4]
  wire  _T_14106; // @[Mux.scala 46:19:@10710.4]
  wire [7:0] _T_14107; // @[Mux.scala 46:16:@10711.4]
  wire  _T_14108; // @[Mux.scala 46:19:@10712.4]
  wire [7:0] _T_14109; // @[Mux.scala 46:16:@10713.4]
  wire  _T_14110; // @[Mux.scala 46:19:@10714.4]
  wire [7:0] _T_14111; // @[Mux.scala 46:16:@10715.4]
  wire  _T_14112; // @[Mux.scala 46:19:@10716.4]
  wire [7:0] _T_14113; // @[Mux.scala 46:16:@10717.4]
  wire  _T_14114; // @[Mux.scala 46:19:@10718.4]
  wire [7:0] _T_14115; // @[Mux.scala 46:16:@10719.4]
  wire  _T_14116; // @[Mux.scala 46:19:@10720.4]
  wire [7:0] _T_14117; // @[Mux.scala 46:16:@10721.4]
  wire  _T_14118; // @[Mux.scala 46:19:@10722.4]
  wire [7:0] _T_14119; // @[Mux.scala 46:16:@10723.4]
  wire  _T_14120; // @[Mux.scala 46:19:@10724.4]
  wire [7:0] _T_14121; // @[Mux.scala 46:16:@10725.4]
  wire  _T_14122; // @[Mux.scala 46:19:@10726.4]
  wire [7:0] _T_14123; // @[Mux.scala 46:16:@10727.4]
  wire  _T_14124; // @[Mux.scala 46:19:@10728.4]
  wire [7:0] _T_14125; // @[Mux.scala 46:16:@10729.4]
  wire  _T_14126; // @[Mux.scala 46:19:@10730.4]
  wire [7:0] _T_14127; // @[Mux.scala 46:16:@10731.4]
  wire  _T_14128; // @[Mux.scala 46:19:@10732.4]
  wire [7:0] _T_14129; // @[Mux.scala 46:16:@10733.4]
  wire  _T_14130; // @[Mux.scala 46:19:@10734.4]
  wire [7:0] _T_14131; // @[Mux.scala 46:16:@10735.4]
  wire  _T_14132; // @[Mux.scala 46:19:@10736.4]
  wire [7:0] _T_14133; // @[Mux.scala 46:16:@10737.4]
  wire  _T_14134; // @[Mux.scala 46:19:@10738.4]
  wire [7:0] _T_14135; // @[Mux.scala 46:16:@10739.4]
  wire  _T_14136; // @[Mux.scala 46:19:@10740.4]
  wire [7:0] _T_14137; // @[Mux.scala 46:16:@10741.4]
  wire  _T_14138; // @[Mux.scala 46:19:@10742.4]
  wire [7:0] _T_14139; // @[Mux.scala 46:16:@10743.4]
  wire  _T_14183; // @[Mux.scala 46:19:@10745.4]
  wire [7:0] _T_14184; // @[Mux.scala 46:16:@10746.4]
  wire  _T_14185; // @[Mux.scala 46:19:@10747.4]
  wire [7:0] _T_14186; // @[Mux.scala 46:16:@10748.4]
  wire  _T_14187; // @[Mux.scala 46:19:@10749.4]
  wire [7:0] _T_14188; // @[Mux.scala 46:16:@10750.4]
  wire  _T_14189; // @[Mux.scala 46:19:@10751.4]
  wire [7:0] _T_14190; // @[Mux.scala 46:16:@10752.4]
  wire  _T_14191; // @[Mux.scala 46:19:@10753.4]
  wire [7:0] _T_14192; // @[Mux.scala 46:16:@10754.4]
  wire  _T_14193; // @[Mux.scala 46:19:@10755.4]
  wire [7:0] _T_14194; // @[Mux.scala 46:16:@10756.4]
  wire  _T_14195; // @[Mux.scala 46:19:@10757.4]
  wire [7:0] _T_14196; // @[Mux.scala 46:16:@10758.4]
  wire  _T_14197; // @[Mux.scala 46:19:@10759.4]
  wire [7:0] _T_14198; // @[Mux.scala 46:16:@10760.4]
  wire  _T_14199; // @[Mux.scala 46:19:@10761.4]
  wire [7:0] _T_14200; // @[Mux.scala 46:16:@10762.4]
  wire  _T_14201; // @[Mux.scala 46:19:@10763.4]
  wire [7:0] _T_14202; // @[Mux.scala 46:16:@10764.4]
  wire  _T_14203; // @[Mux.scala 46:19:@10765.4]
  wire [7:0] _T_14204; // @[Mux.scala 46:16:@10766.4]
  wire  _T_14205; // @[Mux.scala 46:19:@10767.4]
  wire [7:0] _T_14206; // @[Mux.scala 46:16:@10768.4]
  wire  _T_14207; // @[Mux.scala 46:19:@10769.4]
  wire [7:0] _T_14208; // @[Mux.scala 46:16:@10770.4]
  wire  _T_14209; // @[Mux.scala 46:19:@10771.4]
  wire [7:0] _T_14210; // @[Mux.scala 46:16:@10772.4]
  wire  _T_14211; // @[Mux.scala 46:19:@10773.4]
  wire [7:0] _T_14212; // @[Mux.scala 46:16:@10774.4]
  wire  _T_14213; // @[Mux.scala 46:19:@10775.4]
  wire [7:0] _T_14214; // @[Mux.scala 46:16:@10776.4]
  wire  _T_14215; // @[Mux.scala 46:19:@10777.4]
  wire [7:0] _T_14216; // @[Mux.scala 46:16:@10778.4]
  wire  _T_14217; // @[Mux.scala 46:19:@10779.4]
  wire [7:0] _T_14218; // @[Mux.scala 46:16:@10780.4]
  wire  _T_14219; // @[Mux.scala 46:19:@10781.4]
  wire [7:0] _T_14220; // @[Mux.scala 46:16:@10782.4]
  wire  _T_14221; // @[Mux.scala 46:19:@10783.4]
  wire [7:0] _T_14222; // @[Mux.scala 46:16:@10784.4]
  wire  _T_14223; // @[Mux.scala 46:19:@10785.4]
  wire [7:0] _T_14224; // @[Mux.scala 46:16:@10786.4]
  wire  _T_14225; // @[Mux.scala 46:19:@10787.4]
  wire [7:0] _T_14226; // @[Mux.scala 46:16:@10788.4]
  wire  _T_14227; // @[Mux.scala 46:19:@10789.4]
  wire [7:0] _T_14228; // @[Mux.scala 46:16:@10790.4]
  wire  _T_14229; // @[Mux.scala 46:19:@10791.4]
  wire [7:0] _T_14230; // @[Mux.scala 46:16:@10792.4]
  wire  _T_14231; // @[Mux.scala 46:19:@10793.4]
  wire [7:0] _T_14232; // @[Mux.scala 46:16:@10794.4]
  wire  _T_14233; // @[Mux.scala 46:19:@10795.4]
  wire [7:0] _T_14234; // @[Mux.scala 46:16:@10796.4]
  wire  _T_14235; // @[Mux.scala 46:19:@10797.4]
  wire [7:0] _T_14236; // @[Mux.scala 46:16:@10798.4]
  wire  _T_14237; // @[Mux.scala 46:19:@10799.4]
  wire [7:0] _T_14238; // @[Mux.scala 46:16:@10800.4]
  wire  _T_14239; // @[Mux.scala 46:19:@10801.4]
  wire [7:0] _T_14240; // @[Mux.scala 46:16:@10802.4]
  wire  _T_14241; // @[Mux.scala 46:19:@10803.4]
  wire [7:0] _T_14242; // @[Mux.scala 46:16:@10804.4]
  wire  _T_14243; // @[Mux.scala 46:19:@10805.4]
  wire [7:0] _T_14244; // @[Mux.scala 46:16:@10806.4]
  wire  _T_14245; // @[Mux.scala 46:19:@10807.4]
  wire [7:0] _T_14246; // @[Mux.scala 46:16:@10808.4]
  wire  _T_14247; // @[Mux.scala 46:19:@10809.4]
  wire [7:0] _T_14248; // @[Mux.scala 46:16:@10810.4]
  wire  _T_14249; // @[Mux.scala 46:19:@10811.4]
  wire [7:0] _T_14250; // @[Mux.scala 46:16:@10812.4]
  wire  _T_14251; // @[Mux.scala 46:19:@10813.4]
  wire [7:0] _T_14252; // @[Mux.scala 46:16:@10814.4]
  wire  _T_14253; // @[Mux.scala 46:19:@10815.4]
  wire [7:0] _T_14254; // @[Mux.scala 46:16:@10816.4]
  wire  _T_14255; // @[Mux.scala 46:19:@10817.4]
  wire [7:0] _T_14256; // @[Mux.scala 46:16:@10818.4]
  wire  _T_14257; // @[Mux.scala 46:19:@10819.4]
  wire [7:0] _T_14258; // @[Mux.scala 46:16:@10820.4]
  wire  _T_14259; // @[Mux.scala 46:19:@10821.4]
  wire [7:0] _T_14260; // @[Mux.scala 46:16:@10822.4]
  wire  _T_14261; // @[Mux.scala 46:19:@10823.4]
  wire [7:0] _T_14262; // @[Mux.scala 46:16:@10824.4]
  wire  _T_14263; // @[Mux.scala 46:19:@10825.4]
  wire [7:0] _T_14264; // @[Mux.scala 46:16:@10826.4]
  wire  _T_14265; // @[Mux.scala 46:19:@10827.4]
  wire [7:0] _T_14266; // @[Mux.scala 46:16:@10828.4]
  wire  _T_14311; // @[Mux.scala 46:19:@10830.4]
  wire [7:0] _T_14312; // @[Mux.scala 46:16:@10831.4]
  wire  _T_14313; // @[Mux.scala 46:19:@10832.4]
  wire [7:0] _T_14314; // @[Mux.scala 46:16:@10833.4]
  wire  _T_14315; // @[Mux.scala 46:19:@10834.4]
  wire [7:0] _T_14316; // @[Mux.scala 46:16:@10835.4]
  wire  _T_14317; // @[Mux.scala 46:19:@10836.4]
  wire [7:0] _T_14318; // @[Mux.scala 46:16:@10837.4]
  wire  _T_14319; // @[Mux.scala 46:19:@10838.4]
  wire [7:0] _T_14320; // @[Mux.scala 46:16:@10839.4]
  wire  _T_14321; // @[Mux.scala 46:19:@10840.4]
  wire [7:0] _T_14322; // @[Mux.scala 46:16:@10841.4]
  wire  _T_14323; // @[Mux.scala 46:19:@10842.4]
  wire [7:0] _T_14324; // @[Mux.scala 46:16:@10843.4]
  wire  _T_14325; // @[Mux.scala 46:19:@10844.4]
  wire [7:0] _T_14326; // @[Mux.scala 46:16:@10845.4]
  wire  _T_14327; // @[Mux.scala 46:19:@10846.4]
  wire [7:0] _T_14328; // @[Mux.scala 46:16:@10847.4]
  wire  _T_14329; // @[Mux.scala 46:19:@10848.4]
  wire [7:0] _T_14330; // @[Mux.scala 46:16:@10849.4]
  wire  _T_14331; // @[Mux.scala 46:19:@10850.4]
  wire [7:0] _T_14332; // @[Mux.scala 46:16:@10851.4]
  wire  _T_14333; // @[Mux.scala 46:19:@10852.4]
  wire [7:0] _T_14334; // @[Mux.scala 46:16:@10853.4]
  wire  _T_14335; // @[Mux.scala 46:19:@10854.4]
  wire [7:0] _T_14336; // @[Mux.scala 46:16:@10855.4]
  wire  _T_14337; // @[Mux.scala 46:19:@10856.4]
  wire [7:0] _T_14338; // @[Mux.scala 46:16:@10857.4]
  wire  _T_14339; // @[Mux.scala 46:19:@10858.4]
  wire [7:0] _T_14340; // @[Mux.scala 46:16:@10859.4]
  wire  _T_14341; // @[Mux.scala 46:19:@10860.4]
  wire [7:0] _T_14342; // @[Mux.scala 46:16:@10861.4]
  wire  _T_14343; // @[Mux.scala 46:19:@10862.4]
  wire [7:0] _T_14344; // @[Mux.scala 46:16:@10863.4]
  wire  _T_14345; // @[Mux.scala 46:19:@10864.4]
  wire [7:0] _T_14346; // @[Mux.scala 46:16:@10865.4]
  wire  _T_14347; // @[Mux.scala 46:19:@10866.4]
  wire [7:0] _T_14348; // @[Mux.scala 46:16:@10867.4]
  wire  _T_14349; // @[Mux.scala 46:19:@10868.4]
  wire [7:0] _T_14350; // @[Mux.scala 46:16:@10869.4]
  wire  _T_14351; // @[Mux.scala 46:19:@10870.4]
  wire [7:0] _T_14352; // @[Mux.scala 46:16:@10871.4]
  wire  _T_14353; // @[Mux.scala 46:19:@10872.4]
  wire [7:0] _T_14354; // @[Mux.scala 46:16:@10873.4]
  wire  _T_14355; // @[Mux.scala 46:19:@10874.4]
  wire [7:0] _T_14356; // @[Mux.scala 46:16:@10875.4]
  wire  _T_14357; // @[Mux.scala 46:19:@10876.4]
  wire [7:0] _T_14358; // @[Mux.scala 46:16:@10877.4]
  wire  _T_14359; // @[Mux.scala 46:19:@10878.4]
  wire [7:0] _T_14360; // @[Mux.scala 46:16:@10879.4]
  wire  _T_14361; // @[Mux.scala 46:19:@10880.4]
  wire [7:0] _T_14362; // @[Mux.scala 46:16:@10881.4]
  wire  _T_14363; // @[Mux.scala 46:19:@10882.4]
  wire [7:0] _T_14364; // @[Mux.scala 46:16:@10883.4]
  wire  _T_14365; // @[Mux.scala 46:19:@10884.4]
  wire [7:0] _T_14366; // @[Mux.scala 46:16:@10885.4]
  wire  _T_14367; // @[Mux.scala 46:19:@10886.4]
  wire [7:0] _T_14368; // @[Mux.scala 46:16:@10887.4]
  wire  _T_14369; // @[Mux.scala 46:19:@10888.4]
  wire [7:0] _T_14370; // @[Mux.scala 46:16:@10889.4]
  wire  _T_14371; // @[Mux.scala 46:19:@10890.4]
  wire [7:0] _T_14372; // @[Mux.scala 46:16:@10891.4]
  wire  _T_14373; // @[Mux.scala 46:19:@10892.4]
  wire [7:0] _T_14374; // @[Mux.scala 46:16:@10893.4]
  wire  _T_14375; // @[Mux.scala 46:19:@10894.4]
  wire [7:0] _T_14376; // @[Mux.scala 46:16:@10895.4]
  wire  _T_14377; // @[Mux.scala 46:19:@10896.4]
  wire [7:0] _T_14378; // @[Mux.scala 46:16:@10897.4]
  wire  _T_14379; // @[Mux.scala 46:19:@10898.4]
  wire [7:0] _T_14380; // @[Mux.scala 46:16:@10899.4]
  wire  _T_14381; // @[Mux.scala 46:19:@10900.4]
  wire [7:0] _T_14382; // @[Mux.scala 46:16:@10901.4]
  wire  _T_14383; // @[Mux.scala 46:19:@10902.4]
  wire [7:0] _T_14384; // @[Mux.scala 46:16:@10903.4]
  wire  _T_14385; // @[Mux.scala 46:19:@10904.4]
  wire [7:0] _T_14386; // @[Mux.scala 46:16:@10905.4]
  wire  _T_14387; // @[Mux.scala 46:19:@10906.4]
  wire [7:0] _T_14388; // @[Mux.scala 46:16:@10907.4]
  wire  _T_14389; // @[Mux.scala 46:19:@10908.4]
  wire [7:0] _T_14390; // @[Mux.scala 46:16:@10909.4]
  wire  _T_14391; // @[Mux.scala 46:19:@10910.4]
  wire [7:0] _T_14392; // @[Mux.scala 46:16:@10911.4]
  wire  _T_14393; // @[Mux.scala 46:19:@10912.4]
  wire [7:0] _T_14394; // @[Mux.scala 46:16:@10913.4]
  wire  _T_14395; // @[Mux.scala 46:19:@10914.4]
  wire [7:0] _T_14396; // @[Mux.scala 46:16:@10915.4]
  wire  _T_14442; // @[Mux.scala 46:19:@10917.4]
  wire [7:0] _T_14443; // @[Mux.scala 46:16:@10918.4]
  wire  _T_14444; // @[Mux.scala 46:19:@10919.4]
  wire [7:0] _T_14445; // @[Mux.scala 46:16:@10920.4]
  wire  _T_14446; // @[Mux.scala 46:19:@10921.4]
  wire [7:0] _T_14447; // @[Mux.scala 46:16:@10922.4]
  wire  _T_14448; // @[Mux.scala 46:19:@10923.4]
  wire [7:0] _T_14449; // @[Mux.scala 46:16:@10924.4]
  wire  _T_14450; // @[Mux.scala 46:19:@10925.4]
  wire [7:0] _T_14451; // @[Mux.scala 46:16:@10926.4]
  wire  _T_14452; // @[Mux.scala 46:19:@10927.4]
  wire [7:0] _T_14453; // @[Mux.scala 46:16:@10928.4]
  wire  _T_14454; // @[Mux.scala 46:19:@10929.4]
  wire [7:0] _T_14455; // @[Mux.scala 46:16:@10930.4]
  wire  _T_14456; // @[Mux.scala 46:19:@10931.4]
  wire [7:0] _T_14457; // @[Mux.scala 46:16:@10932.4]
  wire  _T_14458; // @[Mux.scala 46:19:@10933.4]
  wire [7:0] _T_14459; // @[Mux.scala 46:16:@10934.4]
  wire  _T_14460; // @[Mux.scala 46:19:@10935.4]
  wire [7:0] _T_14461; // @[Mux.scala 46:16:@10936.4]
  wire  _T_14462; // @[Mux.scala 46:19:@10937.4]
  wire [7:0] _T_14463; // @[Mux.scala 46:16:@10938.4]
  wire  _T_14464; // @[Mux.scala 46:19:@10939.4]
  wire [7:0] _T_14465; // @[Mux.scala 46:16:@10940.4]
  wire  _T_14466; // @[Mux.scala 46:19:@10941.4]
  wire [7:0] _T_14467; // @[Mux.scala 46:16:@10942.4]
  wire  _T_14468; // @[Mux.scala 46:19:@10943.4]
  wire [7:0] _T_14469; // @[Mux.scala 46:16:@10944.4]
  wire  _T_14470; // @[Mux.scala 46:19:@10945.4]
  wire [7:0] _T_14471; // @[Mux.scala 46:16:@10946.4]
  wire  _T_14472; // @[Mux.scala 46:19:@10947.4]
  wire [7:0] _T_14473; // @[Mux.scala 46:16:@10948.4]
  wire  _T_14474; // @[Mux.scala 46:19:@10949.4]
  wire [7:0] _T_14475; // @[Mux.scala 46:16:@10950.4]
  wire  _T_14476; // @[Mux.scala 46:19:@10951.4]
  wire [7:0] _T_14477; // @[Mux.scala 46:16:@10952.4]
  wire  _T_14478; // @[Mux.scala 46:19:@10953.4]
  wire [7:0] _T_14479; // @[Mux.scala 46:16:@10954.4]
  wire  _T_14480; // @[Mux.scala 46:19:@10955.4]
  wire [7:0] _T_14481; // @[Mux.scala 46:16:@10956.4]
  wire  _T_14482; // @[Mux.scala 46:19:@10957.4]
  wire [7:0] _T_14483; // @[Mux.scala 46:16:@10958.4]
  wire  _T_14484; // @[Mux.scala 46:19:@10959.4]
  wire [7:0] _T_14485; // @[Mux.scala 46:16:@10960.4]
  wire  _T_14486; // @[Mux.scala 46:19:@10961.4]
  wire [7:0] _T_14487; // @[Mux.scala 46:16:@10962.4]
  wire  _T_14488; // @[Mux.scala 46:19:@10963.4]
  wire [7:0] _T_14489; // @[Mux.scala 46:16:@10964.4]
  wire  _T_14490; // @[Mux.scala 46:19:@10965.4]
  wire [7:0] _T_14491; // @[Mux.scala 46:16:@10966.4]
  wire  _T_14492; // @[Mux.scala 46:19:@10967.4]
  wire [7:0] _T_14493; // @[Mux.scala 46:16:@10968.4]
  wire  _T_14494; // @[Mux.scala 46:19:@10969.4]
  wire [7:0] _T_14495; // @[Mux.scala 46:16:@10970.4]
  wire  _T_14496; // @[Mux.scala 46:19:@10971.4]
  wire [7:0] _T_14497; // @[Mux.scala 46:16:@10972.4]
  wire  _T_14498; // @[Mux.scala 46:19:@10973.4]
  wire [7:0] _T_14499; // @[Mux.scala 46:16:@10974.4]
  wire  _T_14500; // @[Mux.scala 46:19:@10975.4]
  wire [7:0] _T_14501; // @[Mux.scala 46:16:@10976.4]
  wire  _T_14502; // @[Mux.scala 46:19:@10977.4]
  wire [7:0] _T_14503; // @[Mux.scala 46:16:@10978.4]
  wire  _T_14504; // @[Mux.scala 46:19:@10979.4]
  wire [7:0] _T_14505; // @[Mux.scala 46:16:@10980.4]
  wire  _T_14506; // @[Mux.scala 46:19:@10981.4]
  wire [7:0] _T_14507; // @[Mux.scala 46:16:@10982.4]
  wire  _T_14508; // @[Mux.scala 46:19:@10983.4]
  wire [7:0] _T_14509; // @[Mux.scala 46:16:@10984.4]
  wire  _T_14510; // @[Mux.scala 46:19:@10985.4]
  wire [7:0] _T_14511; // @[Mux.scala 46:16:@10986.4]
  wire  _T_14512; // @[Mux.scala 46:19:@10987.4]
  wire [7:0] _T_14513; // @[Mux.scala 46:16:@10988.4]
  wire  _T_14514; // @[Mux.scala 46:19:@10989.4]
  wire [7:0] _T_14515; // @[Mux.scala 46:16:@10990.4]
  wire  _T_14516; // @[Mux.scala 46:19:@10991.4]
  wire [7:0] _T_14517; // @[Mux.scala 46:16:@10992.4]
  wire  _T_14518; // @[Mux.scala 46:19:@10993.4]
  wire [7:0] _T_14519; // @[Mux.scala 46:16:@10994.4]
  wire  _T_14520; // @[Mux.scala 46:19:@10995.4]
  wire [7:0] _T_14521; // @[Mux.scala 46:16:@10996.4]
  wire  _T_14522; // @[Mux.scala 46:19:@10997.4]
  wire [7:0] _T_14523; // @[Mux.scala 46:16:@10998.4]
  wire  _T_14524; // @[Mux.scala 46:19:@10999.4]
  wire [7:0] _T_14525; // @[Mux.scala 46:16:@11000.4]
  wire  _T_14526; // @[Mux.scala 46:19:@11001.4]
  wire [7:0] _T_14527; // @[Mux.scala 46:16:@11002.4]
  wire  _T_14528; // @[Mux.scala 46:19:@11003.4]
  wire [7:0] _T_14529; // @[Mux.scala 46:16:@11004.4]
  wire  _T_14576; // @[Mux.scala 46:19:@11006.4]
  wire [7:0] _T_14577; // @[Mux.scala 46:16:@11007.4]
  wire  _T_14578; // @[Mux.scala 46:19:@11008.4]
  wire [7:0] _T_14579; // @[Mux.scala 46:16:@11009.4]
  wire  _T_14580; // @[Mux.scala 46:19:@11010.4]
  wire [7:0] _T_14581; // @[Mux.scala 46:16:@11011.4]
  wire  _T_14582; // @[Mux.scala 46:19:@11012.4]
  wire [7:0] _T_14583; // @[Mux.scala 46:16:@11013.4]
  wire  _T_14584; // @[Mux.scala 46:19:@11014.4]
  wire [7:0] _T_14585; // @[Mux.scala 46:16:@11015.4]
  wire  _T_14586; // @[Mux.scala 46:19:@11016.4]
  wire [7:0] _T_14587; // @[Mux.scala 46:16:@11017.4]
  wire  _T_14588; // @[Mux.scala 46:19:@11018.4]
  wire [7:0] _T_14589; // @[Mux.scala 46:16:@11019.4]
  wire  _T_14590; // @[Mux.scala 46:19:@11020.4]
  wire [7:0] _T_14591; // @[Mux.scala 46:16:@11021.4]
  wire  _T_14592; // @[Mux.scala 46:19:@11022.4]
  wire [7:0] _T_14593; // @[Mux.scala 46:16:@11023.4]
  wire  _T_14594; // @[Mux.scala 46:19:@11024.4]
  wire [7:0] _T_14595; // @[Mux.scala 46:16:@11025.4]
  wire  _T_14596; // @[Mux.scala 46:19:@11026.4]
  wire [7:0] _T_14597; // @[Mux.scala 46:16:@11027.4]
  wire  _T_14598; // @[Mux.scala 46:19:@11028.4]
  wire [7:0] _T_14599; // @[Mux.scala 46:16:@11029.4]
  wire  _T_14600; // @[Mux.scala 46:19:@11030.4]
  wire [7:0] _T_14601; // @[Mux.scala 46:16:@11031.4]
  wire  _T_14602; // @[Mux.scala 46:19:@11032.4]
  wire [7:0] _T_14603; // @[Mux.scala 46:16:@11033.4]
  wire  _T_14604; // @[Mux.scala 46:19:@11034.4]
  wire [7:0] _T_14605; // @[Mux.scala 46:16:@11035.4]
  wire  _T_14606; // @[Mux.scala 46:19:@11036.4]
  wire [7:0] _T_14607; // @[Mux.scala 46:16:@11037.4]
  wire  _T_14608; // @[Mux.scala 46:19:@11038.4]
  wire [7:0] _T_14609; // @[Mux.scala 46:16:@11039.4]
  wire  _T_14610; // @[Mux.scala 46:19:@11040.4]
  wire [7:0] _T_14611; // @[Mux.scala 46:16:@11041.4]
  wire  _T_14612; // @[Mux.scala 46:19:@11042.4]
  wire [7:0] _T_14613; // @[Mux.scala 46:16:@11043.4]
  wire  _T_14614; // @[Mux.scala 46:19:@11044.4]
  wire [7:0] _T_14615; // @[Mux.scala 46:16:@11045.4]
  wire  _T_14616; // @[Mux.scala 46:19:@11046.4]
  wire [7:0] _T_14617; // @[Mux.scala 46:16:@11047.4]
  wire  _T_14618; // @[Mux.scala 46:19:@11048.4]
  wire [7:0] _T_14619; // @[Mux.scala 46:16:@11049.4]
  wire  _T_14620; // @[Mux.scala 46:19:@11050.4]
  wire [7:0] _T_14621; // @[Mux.scala 46:16:@11051.4]
  wire  _T_14622; // @[Mux.scala 46:19:@11052.4]
  wire [7:0] _T_14623; // @[Mux.scala 46:16:@11053.4]
  wire  _T_14624; // @[Mux.scala 46:19:@11054.4]
  wire [7:0] _T_14625; // @[Mux.scala 46:16:@11055.4]
  wire  _T_14626; // @[Mux.scala 46:19:@11056.4]
  wire [7:0] _T_14627; // @[Mux.scala 46:16:@11057.4]
  wire  _T_14628; // @[Mux.scala 46:19:@11058.4]
  wire [7:0] _T_14629; // @[Mux.scala 46:16:@11059.4]
  wire  _T_14630; // @[Mux.scala 46:19:@11060.4]
  wire [7:0] _T_14631; // @[Mux.scala 46:16:@11061.4]
  wire  _T_14632; // @[Mux.scala 46:19:@11062.4]
  wire [7:0] _T_14633; // @[Mux.scala 46:16:@11063.4]
  wire  _T_14634; // @[Mux.scala 46:19:@11064.4]
  wire [7:0] _T_14635; // @[Mux.scala 46:16:@11065.4]
  wire  _T_14636; // @[Mux.scala 46:19:@11066.4]
  wire [7:0] _T_14637; // @[Mux.scala 46:16:@11067.4]
  wire  _T_14638; // @[Mux.scala 46:19:@11068.4]
  wire [7:0] _T_14639; // @[Mux.scala 46:16:@11069.4]
  wire  _T_14640; // @[Mux.scala 46:19:@11070.4]
  wire [7:0] _T_14641; // @[Mux.scala 46:16:@11071.4]
  wire  _T_14642; // @[Mux.scala 46:19:@11072.4]
  wire [7:0] _T_14643; // @[Mux.scala 46:16:@11073.4]
  wire  _T_14644; // @[Mux.scala 46:19:@11074.4]
  wire [7:0] _T_14645; // @[Mux.scala 46:16:@11075.4]
  wire  _T_14646; // @[Mux.scala 46:19:@11076.4]
  wire [7:0] _T_14647; // @[Mux.scala 46:16:@11077.4]
  wire  _T_14648; // @[Mux.scala 46:19:@11078.4]
  wire [7:0] _T_14649; // @[Mux.scala 46:16:@11079.4]
  wire  _T_14650; // @[Mux.scala 46:19:@11080.4]
  wire [7:0] _T_14651; // @[Mux.scala 46:16:@11081.4]
  wire  _T_14652; // @[Mux.scala 46:19:@11082.4]
  wire [7:0] _T_14653; // @[Mux.scala 46:16:@11083.4]
  wire  _T_14654; // @[Mux.scala 46:19:@11084.4]
  wire [7:0] _T_14655; // @[Mux.scala 46:16:@11085.4]
  wire  _T_14656; // @[Mux.scala 46:19:@11086.4]
  wire [7:0] _T_14657; // @[Mux.scala 46:16:@11087.4]
  wire  _T_14658; // @[Mux.scala 46:19:@11088.4]
  wire [7:0] _T_14659; // @[Mux.scala 46:16:@11089.4]
  wire  _T_14660; // @[Mux.scala 46:19:@11090.4]
  wire [7:0] _T_14661; // @[Mux.scala 46:16:@11091.4]
  wire  _T_14662; // @[Mux.scala 46:19:@11092.4]
  wire [7:0] _T_14663; // @[Mux.scala 46:16:@11093.4]
  wire  _T_14664; // @[Mux.scala 46:19:@11094.4]
  wire [7:0] _T_14665; // @[Mux.scala 46:16:@11095.4]
  wire  _T_14713; // @[Mux.scala 46:19:@11097.4]
  wire [7:0] _T_14714; // @[Mux.scala 46:16:@11098.4]
  wire  _T_14715; // @[Mux.scala 46:19:@11099.4]
  wire [7:0] _T_14716; // @[Mux.scala 46:16:@11100.4]
  wire  _T_14717; // @[Mux.scala 46:19:@11101.4]
  wire [7:0] _T_14718; // @[Mux.scala 46:16:@11102.4]
  wire  _T_14719; // @[Mux.scala 46:19:@11103.4]
  wire [7:0] _T_14720; // @[Mux.scala 46:16:@11104.4]
  wire  _T_14721; // @[Mux.scala 46:19:@11105.4]
  wire [7:0] _T_14722; // @[Mux.scala 46:16:@11106.4]
  wire  _T_14723; // @[Mux.scala 46:19:@11107.4]
  wire [7:0] _T_14724; // @[Mux.scala 46:16:@11108.4]
  wire  _T_14725; // @[Mux.scala 46:19:@11109.4]
  wire [7:0] _T_14726; // @[Mux.scala 46:16:@11110.4]
  wire  _T_14727; // @[Mux.scala 46:19:@11111.4]
  wire [7:0] _T_14728; // @[Mux.scala 46:16:@11112.4]
  wire  _T_14729; // @[Mux.scala 46:19:@11113.4]
  wire [7:0] _T_14730; // @[Mux.scala 46:16:@11114.4]
  wire  _T_14731; // @[Mux.scala 46:19:@11115.4]
  wire [7:0] _T_14732; // @[Mux.scala 46:16:@11116.4]
  wire  _T_14733; // @[Mux.scala 46:19:@11117.4]
  wire [7:0] _T_14734; // @[Mux.scala 46:16:@11118.4]
  wire  _T_14735; // @[Mux.scala 46:19:@11119.4]
  wire [7:0] _T_14736; // @[Mux.scala 46:16:@11120.4]
  wire  _T_14737; // @[Mux.scala 46:19:@11121.4]
  wire [7:0] _T_14738; // @[Mux.scala 46:16:@11122.4]
  wire  _T_14739; // @[Mux.scala 46:19:@11123.4]
  wire [7:0] _T_14740; // @[Mux.scala 46:16:@11124.4]
  wire  _T_14741; // @[Mux.scala 46:19:@11125.4]
  wire [7:0] _T_14742; // @[Mux.scala 46:16:@11126.4]
  wire  _T_14743; // @[Mux.scala 46:19:@11127.4]
  wire [7:0] _T_14744; // @[Mux.scala 46:16:@11128.4]
  wire  _T_14745; // @[Mux.scala 46:19:@11129.4]
  wire [7:0] _T_14746; // @[Mux.scala 46:16:@11130.4]
  wire  _T_14747; // @[Mux.scala 46:19:@11131.4]
  wire [7:0] _T_14748; // @[Mux.scala 46:16:@11132.4]
  wire  _T_14749; // @[Mux.scala 46:19:@11133.4]
  wire [7:0] _T_14750; // @[Mux.scala 46:16:@11134.4]
  wire  _T_14751; // @[Mux.scala 46:19:@11135.4]
  wire [7:0] _T_14752; // @[Mux.scala 46:16:@11136.4]
  wire  _T_14753; // @[Mux.scala 46:19:@11137.4]
  wire [7:0] _T_14754; // @[Mux.scala 46:16:@11138.4]
  wire  _T_14755; // @[Mux.scala 46:19:@11139.4]
  wire [7:0] _T_14756; // @[Mux.scala 46:16:@11140.4]
  wire  _T_14757; // @[Mux.scala 46:19:@11141.4]
  wire [7:0] _T_14758; // @[Mux.scala 46:16:@11142.4]
  wire  _T_14759; // @[Mux.scala 46:19:@11143.4]
  wire [7:0] _T_14760; // @[Mux.scala 46:16:@11144.4]
  wire  _T_14761; // @[Mux.scala 46:19:@11145.4]
  wire [7:0] _T_14762; // @[Mux.scala 46:16:@11146.4]
  wire  _T_14763; // @[Mux.scala 46:19:@11147.4]
  wire [7:0] _T_14764; // @[Mux.scala 46:16:@11148.4]
  wire  _T_14765; // @[Mux.scala 46:19:@11149.4]
  wire [7:0] _T_14766; // @[Mux.scala 46:16:@11150.4]
  wire  _T_14767; // @[Mux.scala 46:19:@11151.4]
  wire [7:0] _T_14768; // @[Mux.scala 46:16:@11152.4]
  wire  _T_14769; // @[Mux.scala 46:19:@11153.4]
  wire [7:0] _T_14770; // @[Mux.scala 46:16:@11154.4]
  wire  _T_14771; // @[Mux.scala 46:19:@11155.4]
  wire [7:0] _T_14772; // @[Mux.scala 46:16:@11156.4]
  wire  _T_14773; // @[Mux.scala 46:19:@11157.4]
  wire [7:0] _T_14774; // @[Mux.scala 46:16:@11158.4]
  wire  _T_14775; // @[Mux.scala 46:19:@11159.4]
  wire [7:0] _T_14776; // @[Mux.scala 46:16:@11160.4]
  wire  _T_14777; // @[Mux.scala 46:19:@11161.4]
  wire [7:0] _T_14778; // @[Mux.scala 46:16:@11162.4]
  wire  _T_14779; // @[Mux.scala 46:19:@11163.4]
  wire [7:0] _T_14780; // @[Mux.scala 46:16:@11164.4]
  wire  _T_14781; // @[Mux.scala 46:19:@11165.4]
  wire [7:0] _T_14782; // @[Mux.scala 46:16:@11166.4]
  wire  _T_14783; // @[Mux.scala 46:19:@11167.4]
  wire [7:0] _T_14784; // @[Mux.scala 46:16:@11168.4]
  wire  _T_14785; // @[Mux.scala 46:19:@11169.4]
  wire [7:0] _T_14786; // @[Mux.scala 46:16:@11170.4]
  wire  _T_14787; // @[Mux.scala 46:19:@11171.4]
  wire [7:0] _T_14788; // @[Mux.scala 46:16:@11172.4]
  wire  _T_14789; // @[Mux.scala 46:19:@11173.4]
  wire [7:0] _T_14790; // @[Mux.scala 46:16:@11174.4]
  wire  _T_14791; // @[Mux.scala 46:19:@11175.4]
  wire [7:0] _T_14792; // @[Mux.scala 46:16:@11176.4]
  wire  _T_14793; // @[Mux.scala 46:19:@11177.4]
  wire [7:0] _T_14794; // @[Mux.scala 46:16:@11178.4]
  wire  _T_14795; // @[Mux.scala 46:19:@11179.4]
  wire [7:0] _T_14796; // @[Mux.scala 46:16:@11180.4]
  wire  _T_14797; // @[Mux.scala 46:19:@11181.4]
  wire [7:0] _T_14798; // @[Mux.scala 46:16:@11182.4]
  wire  _T_14799; // @[Mux.scala 46:19:@11183.4]
  wire [7:0] _T_14800; // @[Mux.scala 46:16:@11184.4]
  wire  _T_14801; // @[Mux.scala 46:19:@11185.4]
  wire [7:0] _T_14802; // @[Mux.scala 46:16:@11186.4]
  wire  _T_14803; // @[Mux.scala 46:19:@11187.4]
  wire [7:0] _T_14804; // @[Mux.scala 46:16:@11188.4]
  wire  _T_14853; // @[Mux.scala 46:19:@11190.4]
  wire [7:0] _T_14854; // @[Mux.scala 46:16:@11191.4]
  wire  _T_14855; // @[Mux.scala 46:19:@11192.4]
  wire [7:0] _T_14856; // @[Mux.scala 46:16:@11193.4]
  wire  _T_14857; // @[Mux.scala 46:19:@11194.4]
  wire [7:0] _T_14858; // @[Mux.scala 46:16:@11195.4]
  wire  _T_14859; // @[Mux.scala 46:19:@11196.4]
  wire [7:0] _T_14860; // @[Mux.scala 46:16:@11197.4]
  wire  _T_14861; // @[Mux.scala 46:19:@11198.4]
  wire [7:0] _T_14862; // @[Mux.scala 46:16:@11199.4]
  wire  _T_14863; // @[Mux.scala 46:19:@11200.4]
  wire [7:0] _T_14864; // @[Mux.scala 46:16:@11201.4]
  wire  _T_14865; // @[Mux.scala 46:19:@11202.4]
  wire [7:0] _T_14866; // @[Mux.scala 46:16:@11203.4]
  wire  _T_14867; // @[Mux.scala 46:19:@11204.4]
  wire [7:0] _T_14868; // @[Mux.scala 46:16:@11205.4]
  wire  _T_14869; // @[Mux.scala 46:19:@11206.4]
  wire [7:0] _T_14870; // @[Mux.scala 46:16:@11207.4]
  wire  _T_14871; // @[Mux.scala 46:19:@11208.4]
  wire [7:0] _T_14872; // @[Mux.scala 46:16:@11209.4]
  wire  _T_14873; // @[Mux.scala 46:19:@11210.4]
  wire [7:0] _T_14874; // @[Mux.scala 46:16:@11211.4]
  wire  _T_14875; // @[Mux.scala 46:19:@11212.4]
  wire [7:0] _T_14876; // @[Mux.scala 46:16:@11213.4]
  wire  _T_14877; // @[Mux.scala 46:19:@11214.4]
  wire [7:0] _T_14878; // @[Mux.scala 46:16:@11215.4]
  wire  _T_14879; // @[Mux.scala 46:19:@11216.4]
  wire [7:0] _T_14880; // @[Mux.scala 46:16:@11217.4]
  wire  _T_14881; // @[Mux.scala 46:19:@11218.4]
  wire [7:0] _T_14882; // @[Mux.scala 46:16:@11219.4]
  wire  _T_14883; // @[Mux.scala 46:19:@11220.4]
  wire [7:0] _T_14884; // @[Mux.scala 46:16:@11221.4]
  wire  _T_14885; // @[Mux.scala 46:19:@11222.4]
  wire [7:0] _T_14886; // @[Mux.scala 46:16:@11223.4]
  wire  _T_14887; // @[Mux.scala 46:19:@11224.4]
  wire [7:0] _T_14888; // @[Mux.scala 46:16:@11225.4]
  wire  _T_14889; // @[Mux.scala 46:19:@11226.4]
  wire [7:0] _T_14890; // @[Mux.scala 46:16:@11227.4]
  wire  _T_14891; // @[Mux.scala 46:19:@11228.4]
  wire [7:0] _T_14892; // @[Mux.scala 46:16:@11229.4]
  wire  _T_14893; // @[Mux.scala 46:19:@11230.4]
  wire [7:0] _T_14894; // @[Mux.scala 46:16:@11231.4]
  wire  _T_14895; // @[Mux.scala 46:19:@11232.4]
  wire [7:0] _T_14896; // @[Mux.scala 46:16:@11233.4]
  wire  _T_14897; // @[Mux.scala 46:19:@11234.4]
  wire [7:0] _T_14898; // @[Mux.scala 46:16:@11235.4]
  wire  _T_14899; // @[Mux.scala 46:19:@11236.4]
  wire [7:0] _T_14900; // @[Mux.scala 46:16:@11237.4]
  wire  _T_14901; // @[Mux.scala 46:19:@11238.4]
  wire [7:0] _T_14902; // @[Mux.scala 46:16:@11239.4]
  wire  _T_14903; // @[Mux.scala 46:19:@11240.4]
  wire [7:0] _T_14904; // @[Mux.scala 46:16:@11241.4]
  wire  _T_14905; // @[Mux.scala 46:19:@11242.4]
  wire [7:0] _T_14906; // @[Mux.scala 46:16:@11243.4]
  wire  _T_14907; // @[Mux.scala 46:19:@11244.4]
  wire [7:0] _T_14908; // @[Mux.scala 46:16:@11245.4]
  wire  _T_14909; // @[Mux.scala 46:19:@11246.4]
  wire [7:0] _T_14910; // @[Mux.scala 46:16:@11247.4]
  wire  _T_14911; // @[Mux.scala 46:19:@11248.4]
  wire [7:0] _T_14912; // @[Mux.scala 46:16:@11249.4]
  wire  _T_14913; // @[Mux.scala 46:19:@11250.4]
  wire [7:0] _T_14914; // @[Mux.scala 46:16:@11251.4]
  wire  _T_14915; // @[Mux.scala 46:19:@11252.4]
  wire [7:0] _T_14916; // @[Mux.scala 46:16:@11253.4]
  wire  _T_14917; // @[Mux.scala 46:19:@11254.4]
  wire [7:0] _T_14918; // @[Mux.scala 46:16:@11255.4]
  wire  _T_14919; // @[Mux.scala 46:19:@11256.4]
  wire [7:0] _T_14920; // @[Mux.scala 46:16:@11257.4]
  wire  _T_14921; // @[Mux.scala 46:19:@11258.4]
  wire [7:0] _T_14922; // @[Mux.scala 46:16:@11259.4]
  wire  _T_14923; // @[Mux.scala 46:19:@11260.4]
  wire [7:0] _T_14924; // @[Mux.scala 46:16:@11261.4]
  wire  _T_14925; // @[Mux.scala 46:19:@11262.4]
  wire [7:0] _T_14926; // @[Mux.scala 46:16:@11263.4]
  wire  _T_14927; // @[Mux.scala 46:19:@11264.4]
  wire [7:0] _T_14928; // @[Mux.scala 46:16:@11265.4]
  wire  _T_14929; // @[Mux.scala 46:19:@11266.4]
  wire [7:0] _T_14930; // @[Mux.scala 46:16:@11267.4]
  wire  _T_14931; // @[Mux.scala 46:19:@11268.4]
  wire [7:0] _T_14932; // @[Mux.scala 46:16:@11269.4]
  wire  _T_14933; // @[Mux.scala 46:19:@11270.4]
  wire [7:0] _T_14934; // @[Mux.scala 46:16:@11271.4]
  wire  _T_14935; // @[Mux.scala 46:19:@11272.4]
  wire [7:0] _T_14936; // @[Mux.scala 46:16:@11273.4]
  wire  _T_14937; // @[Mux.scala 46:19:@11274.4]
  wire [7:0] _T_14938; // @[Mux.scala 46:16:@11275.4]
  wire  _T_14939; // @[Mux.scala 46:19:@11276.4]
  wire [7:0] _T_14940; // @[Mux.scala 46:16:@11277.4]
  wire  _T_14941; // @[Mux.scala 46:19:@11278.4]
  wire [7:0] _T_14942; // @[Mux.scala 46:16:@11279.4]
  wire  _T_14943; // @[Mux.scala 46:19:@11280.4]
  wire [7:0] _T_14944; // @[Mux.scala 46:16:@11281.4]
  wire  _T_14945; // @[Mux.scala 46:19:@11282.4]
  wire [7:0] _T_14946; // @[Mux.scala 46:16:@11283.4]
  wire  _T_14996; // @[Mux.scala 46:19:@11285.4]
  wire [7:0] _T_14997; // @[Mux.scala 46:16:@11286.4]
  wire  _T_14998; // @[Mux.scala 46:19:@11287.4]
  wire [7:0] _T_14999; // @[Mux.scala 46:16:@11288.4]
  wire  _T_15000; // @[Mux.scala 46:19:@11289.4]
  wire [7:0] _T_15001; // @[Mux.scala 46:16:@11290.4]
  wire  _T_15002; // @[Mux.scala 46:19:@11291.4]
  wire [7:0] _T_15003; // @[Mux.scala 46:16:@11292.4]
  wire  _T_15004; // @[Mux.scala 46:19:@11293.4]
  wire [7:0] _T_15005; // @[Mux.scala 46:16:@11294.4]
  wire  _T_15006; // @[Mux.scala 46:19:@11295.4]
  wire [7:0] _T_15007; // @[Mux.scala 46:16:@11296.4]
  wire  _T_15008; // @[Mux.scala 46:19:@11297.4]
  wire [7:0] _T_15009; // @[Mux.scala 46:16:@11298.4]
  wire  _T_15010; // @[Mux.scala 46:19:@11299.4]
  wire [7:0] _T_15011; // @[Mux.scala 46:16:@11300.4]
  wire  _T_15012; // @[Mux.scala 46:19:@11301.4]
  wire [7:0] _T_15013; // @[Mux.scala 46:16:@11302.4]
  wire  _T_15014; // @[Mux.scala 46:19:@11303.4]
  wire [7:0] _T_15015; // @[Mux.scala 46:16:@11304.4]
  wire  _T_15016; // @[Mux.scala 46:19:@11305.4]
  wire [7:0] _T_15017; // @[Mux.scala 46:16:@11306.4]
  wire  _T_15018; // @[Mux.scala 46:19:@11307.4]
  wire [7:0] _T_15019; // @[Mux.scala 46:16:@11308.4]
  wire  _T_15020; // @[Mux.scala 46:19:@11309.4]
  wire [7:0] _T_15021; // @[Mux.scala 46:16:@11310.4]
  wire  _T_15022; // @[Mux.scala 46:19:@11311.4]
  wire [7:0] _T_15023; // @[Mux.scala 46:16:@11312.4]
  wire  _T_15024; // @[Mux.scala 46:19:@11313.4]
  wire [7:0] _T_15025; // @[Mux.scala 46:16:@11314.4]
  wire  _T_15026; // @[Mux.scala 46:19:@11315.4]
  wire [7:0] _T_15027; // @[Mux.scala 46:16:@11316.4]
  wire  _T_15028; // @[Mux.scala 46:19:@11317.4]
  wire [7:0] _T_15029; // @[Mux.scala 46:16:@11318.4]
  wire  _T_15030; // @[Mux.scala 46:19:@11319.4]
  wire [7:0] _T_15031; // @[Mux.scala 46:16:@11320.4]
  wire  _T_15032; // @[Mux.scala 46:19:@11321.4]
  wire [7:0] _T_15033; // @[Mux.scala 46:16:@11322.4]
  wire  _T_15034; // @[Mux.scala 46:19:@11323.4]
  wire [7:0] _T_15035; // @[Mux.scala 46:16:@11324.4]
  wire  _T_15036; // @[Mux.scala 46:19:@11325.4]
  wire [7:0] _T_15037; // @[Mux.scala 46:16:@11326.4]
  wire  _T_15038; // @[Mux.scala 46:19:@11327.4]
  wire [7:0] _T_15039; // @[Mux.scala 46:16:@11328.4]
  wire  _T_15040; // @[Mux.scala 46:19:@11329.4]
  wire [7:0] _T_15041; // @[Mux.scala 46:16:@11330.4]
  wire  _T_15042; // @[Mux.scala 46:19:@11331.4]
  wire [7:0] _T_15043; // @[Mux.scala 46:16:@11332.4]
  wire  _T_15044; // @[Mux.scala 46:19:@11333.4]
  wire [7:0] _T_15045; // @[Mux.scala 46:16:@11334.4]
  wire  _T_15046; // @[Mux.scala 46:19:@11335.4]
  wire [7:0] _T_15047; // @[Mux.scala 46:16:@11336.4]
  wire  _T_15048; // @[Mux.scala 46:19:@11337.4]
  wire [7:0] _T_15049; // @[Mux.scala 46:16:@11338.4]
  wire  _T_15050; // @[Mux.scala 46:19:@11339.4]
  wire [7:0] _T_15051; // @[Mux.scala 46:16:@11340.4]
  wire  _T_15052; // @[Mux.scala 46:19:@11341.4]
  wire [7:0] _T_15053; // @[Mux.scala 46:16:@11342.4]
  wire  _T_15054; // @[Mux.scala 46:19:@11343.4]
  wire [7:0] _T_15055; // @[Mux.scala 46:16:@11344.4]
  wire  _T_15056; // @[Mux.scala 46:19:@11345.4]
  wire [7:0] _T_15057; // @[Mux.scala 46:16:@11346.4]
  wire  _T_15058; // @[Mux.scala 46:19:@11347.4]
  wire [7:0] _T_15059; // @[Mux.scala 46:16:@11348.4]
  wire  _T_15060; // @[Mux.scala 46:19:@11349.4]
  wire [7:0] _T_15061; // @[Mux.scala 46:16:@11350.4]
  wire  _T_15062; // @[Mux.scala 46:19:@11351.4]
  wire [7:0] _T_15063; // @[Mux.scala 46:16:@11352.4]
  wire  _T_15064; // @[Mux.scala 46:19:@11353.4]
  wire [7:0] _T_15065; // @[Mux.scala 46:16:@11354.4]
  wire  _T_15066; // @[Mux.scala 46:19:@11355.4]
  wire [7:0] _T_15067; // @[Mux.scala 46:16:@11356.4]
  wire  _T_15068; // @[Mux.scala 46:19:@11357.4]
  wire [7:0] _T_15069; // @[Mux.scala 46:16:@11358.4]
  wire  _T_15070; // @[Mux.scala 46:19:@11359.4]
  wire [7:0] _T_15071; // @[Mux.scala 46:16:@11360.4]
  wire  _T_15072; // @[Mux.scala 46:19:@11361.4]
  wire [7:0] _T_15073; // @[Mux.scala 46:16:@11362.4]
  wire  _T_15074; // @[Mux.scala 46:19:@11363.4]
  wire [7:0] _T_15075; // @[Mux.scala 46:16:@11364.4]
  wire  _T_15076; // @[Mux.scala 46:19:@11365.4]
  wire [7:0] _T_15077; // @[Mux.scala 46:16:@11366.4]
  wire  _T_15078; // @[Mux.scala 46:19:@11367.4]
  wire [7:0] _T_15079; // @[Mux.scala 46:16:@11368.4]
  wire  _T_15080; // @[Mux.scala 46:19:@11369.4]
  wire [7:0] _T_15081; // @[Mux.scala 46:16:@11370.4]
  wire  _T_15082; // @[Mux.scala 46:19:@11371.4]
  wire [7:0] _T_15083; // @[Mux.scala 46:16:@11372.4]
  wire  _T_15084; // @[Mux.scala 46:19:@11373.4]
  wire [7:0] _T_15085; // @[Mux.scala 46:16:@11374.4]
  wire  _T_15086; // @[Mux.scala 46:19:@11375.4]
  wire [7:0] _T_15087; // @[Mux.scala 46:16:@11376.4]
  wire  _T_15088; // @[Mux.scala 46:19:@11377.4]
  wire [7:0] _T_15089; // @[Mux.scala 46:16:@11378.4]
  wire  _T_15090; // @[Mux.scala 46:19:@11379.4]
  wire [7:0] _T_15091; // @[Mux.scala 46:16:@11380.4]
  wire  _T_15142; // @[Mux.scala 46:19:@11382.4]
  wire [7:0] _T_15143; // @[Mux.scala 46:16:@11383.4]
  wire  _T_15144; // @[Mux.scala 46:19:@11384.4]
  wire [7:0] _T_15145; // @[Mux.scala 46:16:@11385.4]
  wire  _T_15146; // @[Mux.scala 46:19:@11386.4]
  wire [7:0] _T_15147; // @[Mux.scala 46:16:@11387.4]
  wire  _T_15148; // @[Mux.scala 46:19:@11388.4]
  wire [7:0] _T_15149; // @[Mux.scala 46:16:@11389.4]
  wire  _T_15150; // @[Mux.scala 46:19:@11390.4]
  wire [7:0] _T_15151; // @[Mux.scala 46:16:@11391.4]
  wire  _T_15152; // @[Mux.scala 46:19:@11392.4]
  wire [7:0] _T_15153; // @[Mux.scala 46:16:@11393.4]
  wire  _T_15154; // @[Mux.scala 46:19:@11394.4]
  wire [7:0] _T_15155; // @[Mux.scala 46:16:@11395.4]
  wire  _T_15156; // @[Mux.scala 46:19:@11396.4]
  wire [7:0] _T_15157; // @[Mux.scala 46:16:@11397.4]
  wire  _T_15158; // @[Mux.scala 46:19:@11398.4]
  wire [7:0] _T_15159; // @[Mux.scala 46:16:@11399.4]
  wire  _T_15160; // @[Mux.scala 46:19:@11400.4]
  wire [7:0] _T_15161; // @[Mux.scala 46:16:@11401.4]
  wire  _T_15162; // @[Mux.scala 46:19:@11402.4]
  wire [7:0] _T_15163; // @[Mux.scala 46:16:@11403.4]
  wire  _T_15164; // @[Mux.scala 46:19:@11404.4]
  wire [7:0] _T_15165; // @[Mux.scala 46:16:@11405.4]
  wire  _T_15166; // @[Mux.scala 46:19:@11406.4]
  wire [7:0] _T_15167; // @[Mux.scala 46:16:@11407.4]
  wire  _T_15168; // @[Mux.scala 46:19:@11408.4]
  wire [7:0] _T_15169; // @[Mux.scala 46:16:@11409.4]
  wire  _T_15170; // @[Mux.scala 46:19:@11410.4]
  wire [7:0] _T_15171; // @[Mux.scala 46:16:@11411.4]
  wire  _T_15172; // @[Mux.scala 46:19:@11412.4]
  wire [7:0] _T_15173; // @[Mux.scala 46:16:@11413.4]
  wire  _T_15174; // @[Mux.scala 46:19:@11414.4]
  wire [7:0] _T_15175; // @[Mux.scala 46:16:@11415.4]
  wire  _T_15176; // @[Mux.scala 46:19:@11416.4]
  wire [7:0] _T_15177; // @[Mux.scala 46:16:@11417.4]
  wire  _T_15178; // @[Mux.scala 46:19:@11418.4]
  wire [7:0] _T_15179; // @[Mux.scala 46:16:@11419.4]
  wire  _T_15180; // @[Mux.scala 46:19:@11420.4]
  wire [7:0] _T_15181; // @[Mux.scala 46:16:@11421.4]
  wire  _T_15182; // @[Mux.scala 46:19:@11422.4]
  wire [7:0] _T_15183; // @[Mux.scala 46:16:@11423.4]
  wire  _T_15184; // @[Mux.scala 46:19:@11424.4]
  wire [7:0] _T_15185; // @[Mux.scala 46:16:@11425.4]
  wire  _T_15186; // @[Mux.scala 46:19:@11426.4]
  wire [7:0] _T_15187; // @[Mux.scala 46:16:@11427.4]
  wire  _T_15188; // @[Mux.scala 46:19:@11428.4]
  wire [7:0] _T_15189; // @[Mux.scala 46:16:@11429.4]
  wire  _T_15190; // @[Mux.scala 46:19:@11430.4]
  wire [7:0] _T_15191; // @[Mux.scala 46:16:@11431.4]
  wire  _T_15192; // @[Mux.scala 46:19:@11432.4]
  wire [7:0] _T_15193; // @[Mux.scala 46:16:@11433.4]
  wire  _T_15194; // @[Mux.scala 46:19:@11434.4]
  wire [7:0] _T_15195; // @[Mux.scala 46:16:@11435.4]
  wire  _T_15196; // @[Mux.scala 46:19:@11436.4]
  wire [7:0] _T_15197; // @[Mux.scala 46:16:@11437.4]
  wire  _T_15198; // @[Mux.scala 46:19:@11438.4]
  wire [7:0] _T_15199; // @[Mux.scala 46:16:@11439.4]
  wire  _T_15200; // @[Mux.scala 46:19:@11440.4]
  wire [7:0] _T_15201; // @[Mux.scala 46:16:@11441.4]
  wire  _T_15202; // @[Mux.scala 46:19:@11442.4]
  wire [7:0] _T_15203; // @[Mux.scala 46:16:@11443.4]
  wire  _T_15204; // @[Mux.scala 46:19:@11444.4]
  wire [7:0] _T_15205; // @[Mux.scala 46:16:@11445.4]
  wire  _T_15206; // @[Mux.scala 46:19:@11446.4]
  wire [7:0] _T_15207; // @[Mux.scala 46:16:@11447.4]
  wire  _T_15208; // @[Mux.scala 46:19:@11448.4]
  wire [7:0] _T_15209; // @[Mux.scala 46:16:@11449.4]
  wire  _T_15210; // @[Mux.scala 46:19:@11450.4]
  wire [7:0] _T_15211; // @[Mux.scala 46:16:@11451.4]
  wire  _T_15212; // @[Mux.scala 46:19:@11452.4]
  wire [7:0] _T_15213; // @[Mux.scala 46:16:@11453.4]
  wire  _T_15214; // @[Mux.scala 46:19:@11454.4]
  wire [7:0] _T_15215; // @[Mux.scala 46:16:@11455.4]
  wire  _T_15216; // @[Mux.scala 46:19:@11456.4]
  wire [7:0] _T_15217; // @[Mux.scala 46:16:@11457.4]
  wire  _T_15218; // @[Mux.scala 46:19:@11458.4]
  wire [7:0] _T_15219; // @[Mux.scala 46:16:@11459.4]
  wire  _T_15220; // @[Mux.scala 46:19:@11460.4]
  wire [7:0] _T_15221; // @[Mux.scala 46:16:@11461.4]
  wire  _T_15222; // @[Mux.scala 46:19:@11462.4]
  wire [7:0] _T_15223; // @[Mux.scala 46:16:@11463.4]
  wire  _T_15224; // @[Mux.scala 46:19:@11464.4]
  wire [7:0] _T_15225; // @[Mux.scala 46:16:@11465.4]
  wire  _T_15226; // @[Mux.scala 46:19:@11466.4]
  wire [7:0] _T_15227; // @[Mux.scala 46:16:@11467.4]
  wire  _T_15228; // @[Mux.scala 46:19:@11468.4]
  wire [7:0] _T_15229; // @[Mux.scala 46:16:@11469.4]
  wire  _T_15230; // @[Mux.scala 46:19:@11470.4]
  wire [7:0] _T_15231; // @[Mux.scala 46:16:@11471.4]
  wire  _T_15232; // @[Mux.scala 46:19:@11472.4]
  wire [7:0] _T_15233; // @[Mux.scala 46:16:@11473.4]
  wire  _T_15234; // @[Mux.scala 46:19:@11474.4]
  wire [7:0] _T_15235; // @[Mux.scala 46:16:@11475.4]
  wire  _T_15236; // @[Mux.scala 46:19:@11476.4]
  wire [7:0] _T_15237; // @[Mux.scala 46:16:@11477.4]
  wire  _T_15238; // @[Mux.scala 46:19:@11478.4]
  wire [7:0] _T_15239; // @[Mux.scala 46:16:@11479.4]
  wire  _T_15291; // @[Mux.scala 46:19:@11481.4]
  wire [7:0] _T_15292; // @[Mux.scala 46:16:@11482.4]
  wire  _T_15293; // @[Mux.scala 46:19:@11483.4]
  wire [7:0] _T_15294; // @[Mux.scala 46:16:@11484.4]
  wire  _T_15295; // @[Mux.scala 46:19:@11485.4]
  wire [7:0] _T_15296; // @[Mux.scala 46:16:@11486.4]
  wire  _T_15297; // @[Mux.scala 46:19:@11487.4]
  wire [7:0] _T_15298; // @[Mux.scala 46:16:@11488.4]
  wire  _T_15299; // @[Mux.scala 46:19:@11489.4]
  wire [7:0] _T_15300; // @[Mux.scala 46:16:@11490.4]
  wire  _T_15301; // @[Mux.scala 46:19:@11491.4]
  wire [7:0] _T_15302; // @[Mux.scala 46:16:@11492.4]
  wire  _T_15303; // @[Mux.scala 46:19:@11493.4]
  wire [7:0] _T_15304; // @[Mux.scala 46:16:@11494.4]
  wire  _T_15305; // @[Mux.scala 46:19:@11495.4]
  wire [7:0] _T_15306; // @[Mux.scala 46:16:@11496.4]
  wire  _T_15307; // @[Mux.scala 46:19:@11497.4]
  wire [7:0] _T_15308; // @[Mux.scala 46:16:@11498.4]
  wire  _T_15309; // @[Mux.scala 46:19:@11499.4]
  wire [7:0] _T_15310; // @[Mux.scala 46:16:@11500.4]
  wire  _T_15311; // @[Mux.scala 46:19:@11501.4]
  wire [7:0] _T_15312; // @[Mux.scala 46:16:@11502.4]
  wire  _T_15313; // @[Mux.scala 46:19:@11503.4]
  wire [7:0] _T_15314; // @[Mux.scala 46:16:@11504.4]
  wire  _T_15315; // @[Mux.scala 46:19:@11505.4]
  wire [7:0] _T_15316; // @[Mux.scala 46:16:@11506.4]
  wire  _T_15317; // @[Mux.scala 46:19:@11507.4]
  wire [7:0] _T_15318; // @[Mux.scala 46:16:@11508.4]
  wire  _T_15319; // @[Mux.scala 46:19:@11509.4]
  wire [7:0] _T_15320; // @[Mux.scala 46:16:@11510.4]
  wire  _T_15321; // @[Mux.scala 46:19:@11511.4]
  wire [7:0] _T_15322; // @[Mux.scala 46:16:@11512.4]
  wire  _T_15323; // @[Mux.scala 46:19:@11513.4]
  wire [7:0] _T_15324; // @[Mux.scala 46:16:@11514.4]
  wire  _T_15325; // @[Mux.scala 46:19:@11515.4]
  wire [7:0] _T_15326; // @[Mux.scala 46:16:@11516.4]
  wire  _T_15327; // @[Mux.scala 46:19:@11517.4]
  wire [7:0] _T_15328; // @[Mux.scala 46:16:@11518.4]
  wire  _T_15329; // @[Mux.scala 46:19:@11519.4]
  wire [7:0] _T_15330; // @[Mux.scala 46:16:@11520.4]
  wire  _T_15331; // @[Mux.scala 46:19:@11521.4]
  wire [7:0] _T_15332; // @[Mux.scala 46:16:@11522.4]
  wire  _T_15333; // @[Mux.scala 46:19:@11523.4]
  wire [7:0] _T_15334; // @[Mux.scala 46:16:@11524.4]
  wire  _T_15335; // @[Mux.scala 46:19:@11525.4]
  wire [7:0] _T_15336; // @[Mux.scala 46:16:@11526.4]
  wire  _T_15337; // @[Mux.scala 46:19:@11527.4]
  wire [7:0] _T_15338; // @[Mux.scala 46:16:@11528.4]
  wire  _T_15339; // @[Mux.scala 46:19:@11529.4]
  wire [7:0] _T_15340; // @[Mux.scala 46:16:@11530.4]
  wire  _T_15341; // @[Mux.scala 46:19:@11531.4]
  wire [7:0] _T_15342; // @[Mux.scala 46:16:@11532.4]
  wire  _T_15343; // @[Mux.scala 46:19:@11533.4]
  wire [7:0] _T_15344; // @[Mux.scala 46:16:@11534.4]
  wire  _T_15345; // @[Mux.scala 46:19:@11535.4]
  wire [7:0] _T_15346; // @[Mux.scala 46:16:@11536.4]
  wire  _T_15347; // @[Mux.scala 46:19:@11537.4]
  wire [7:0] _T_15348; // @[Mux.scala 46:16:@11538.4]
  wire  _T_15349; // @[Mux.scala 46:19:@11539.4]
  wire [7:0] _T_15350; // @[Mux.scala 46:16:@11540.4]
  wire  _T_15351; // @[Mux.scala 46:19:@11541.4]
  wire [7:0] _T_15352; // @[Mux.scala 46:16:@11542.4]
  wire  _T_15353; // @[Mux.scala 46:19:@11543.4]
  wire [7:0] _T_15354; // @[Mux.scala 46:16:@11544.4]
  wire  _T_15355; // @[Mux.scala 46:19:@11545.4]
  wire [7:0] _T_15356; // @[Mux.scala 46:16:@11546.4]
  wire  _T_15357; // @[Mux.scala 46:19:@11547.4]
  wire [7:0] _T_15358; // @[Mux.scala 46:16:@11548.4]
  wire  _T_15359; // @[Mux.scala 46:19:@11549.4]
  wire [7:0] _T_15360; // @[Mux.scala 46:16:@11550.4]
  wire  _T_15361; // @[Mux.scala 46:19:@11551.4]
  wire [7:0] _T_15362; // @[Mux.scala 46:16:@11552.4]
  wire  _T_15363; // @[Mux.scala 46:19:@11553.4]
  wire [7:0] _T_15364; // @[Mux.scala 46:16:@11554.4]
  wire  _T_15365; // @[Mux.scala 46:19:@11555.4]
  wire [7:0] _T_15366; // @[Mux.scala 46:16:@11556.4]
  wire  _T_15367; // @[Mux.scala 46:19:@11557.4]
  wire [7:0] _T_15368; // @[Mux.scala 46:16:@11558.4]
  wire  _T_15369; // @[Mux.scala 46:19:@11559.4]
  wire [7:0] _T_15370; // @[Mux.scala 46:16:@11560.4]
  wire  _T_15371; // @[Mux.scala 46:19:@11561.4]
  wire [7:0] _T_15372; // @[Mux.scala 46:16:@11562.4]
  wire  _T_15373; // @[Mux.scala 46:19:@11563.4]
  wire [7:0] _T_15374; // @[Mux.scala 46:16:@11564.4]
  wire  _T_15375; // @[Mux.scala 46:19:@11565.4]
  wire [7:0] _T_15376; // @[Mux.scala 46:16:@11566.4]
  wire  _T_15377; // @[Mux.scala 46:19:@11567.4]
  wire [7:0] _T_15378; // @[Mux.scala 46:16:@11568.4]
  wire  _T_15379; // @[Mux.scala 46:19:@11569.4]
  wire [7:0] _T_15380; // @[Mux.scala 46:16:@11570.4]
  wire  _T_15381; // @[Mux.scala 46:19:@11571.4]
  wire [7:0] _T_15382; // @[Mux.scala 46:16:@11572.4]
  wire  _T_15383; // @[Mux.scala 46:19:@11573.4]
  wire [7:0] _T_15384; // @[Mux.scala 46:16:@11574.4]
  wire  _T_15385; // @[Mux.scala 46:19:@11575.4]
  wire [7:0] _T_15386; // @[Mux.scala 46:16:@11576.4]
  wire  _T_15387; // @[Mux.scala 46:19:@11577.4]
  wire [7:0] _T_15388; // @[Mux.scala 46:16:@11578.4]
  wire  _T_15389; // @[Mux.scala 46:19:@11579.4]
  wire [7:0] _T_15390; // @[Mux.scala 46:16:@11580.4]
  wire  _T_15443; // @[Mux.scala 46:19:@11582.4]
  wire [7:0] _T_15444; // @[Mux.scala 46:16:@11583.4]
  wire  _T_15445; // @[Mux.scala 46:19:@11584.4]
  wire [7:0] _T_15446; // @[Mux.scala 46:16:@11585.4]
  wire  _T_15447; // @[Mux.scala 46:19:@11586.4]
  wire [7:0] _T_15448; // @[Mux.scala 46:16:@11587.4]
  wire  _T_15449; // @[Mux.scala 46:19:@11588.4]
  wire [7:0] _T_15450; // @[Mux.scala 46:16:@11589.4]
  wire  _T_15451; // @[Mux.scala 46:19:@11590.4]
  wire [7:0] _T_15452; // @[Mux.scala 46:16:@11591.4]
  wire  _T_15453; // @[Mux.scala 46:19:@11592.4]
  wire [7:0] _T_15454; // @[Mux.scala 46:16:@11593.4]
  wire  _T_15455; // @[Mux.scala 46:19:@11594.4]
  wire [7:0] _T_15456; // @[Mux.scala 46:16:@11595.4]
  wire  _T_15457; // @[Mux.scala 46:19:@11596.4]
  wire [7:0] _T_15458; // @[Mux.scala 46:16:@11597.4]
  wire  _T_15459; // @[Mux.scala 46:19:@11598.4]
  wire [7:0] _T_15460; // @[Mux.scala 46:16:@11599.4]
  wire  _T_15461; // @[Mux.scala 46:19:@11600.4]
  wire [7:0] _T_15462; // @[Mux.scala 46:16:@11601.4]
  wire  _T_15463; // @[Mux.scala 46:19:@11602.4]
  wire [7:0] _T_15464; // @[Mux.scala 46:16:@11603.4]
  wire  _T_15465; // @[Mux.scala 46:19:@11604.4]
  wire [7:0] _T_15466; // @[Mux.scala 46:16:@11605.4]
  wire  _T_15467; // @[Mux.scala 46:19:@11606.4]
  wire [7:0] _T_15468; // @[Mux.scala 46:16:@11607.4]
  wire  _T_15469; // @[Mux.scala 46:19:@11608.4]
  wire [7:0] _T_15470; // @[Mux.scala 46:16:@11609.4]
  wire  _T_15471; // @[Mux.scala 46:19:@11610.4]
  wire [7:0] _T_15472; // @[Mux.scala 46:16:@11611.4]
  wire  _T_15473; // @[Mux.scala 46:19:@11612.4]
  wire [7:0] _T_15474; // @[Mux.scala 46:16:@11613.4]
  wire  _T_15475; // @[Mux.scala 46:19:@11614.4]
  wire [7:0] _T_15476; // @[Mux.scala 46:16:@11615.4]
  wire  _T_15477; // @[Mux.scala 46:19:@11616.4]
  wire [7:0] _T_15478; // @[Mux.scala 46:16:@11617.4]
  wire  _T_15479; // @[Mux.scala 46:19:@11618.4]
  wire [7:0] _T_15480; // @[Mux.scala 46:16:@11619.4]
  wire  _T_15481; // @[Mux.scala 46:19:@11620.4]
  wire [7:0] _T_15482; // @[Mux.scala 46:16:@11621.4]
  wire  _T_15483; // @[Mux.scala 46:19:@11622.4]
  wire [7:0] _T_15484; // @[Mux.scala 46:16:@11623.4]
  wire  _T_15485; // @[Mux.scala 46:19:@11624.4]
  wire [7:0] _T_15486; // @[Mux.scala 46:16:@11625.4]
  wire  _T_15487; // @[Mux.scala 46:19:@11626.4]
  wire [7:0] _T_15488; // @[Mux.scala 46:16:@11627.4]
  wire  _T_15489; // @[Mux.scala 46:19:@11628.4]
  wire [7:0] _T_15490; // @[Mux.scala 46:16:@11629.4]
  wire  _T_15491; // @[Mux.scala 46:19:@11630.4]
  wire [7:0] _T_15492; // @[Mux.scala 46:16:@11631.4]
  wire  _T_15493; // @[Mux.scala 46:19:@11632.4]
  wire [7:0] _T_15494; // @[Mux.scala 46:16:@11633.4]
  wire  _T_15495; // @[Mux.scala 46:19:@11634.4]
  wire [7:0] _T_15496; // @[Mux.scala 46:16:@11635.4]
  wire  _T_15497; // @[Mux.scala 46:19:@11636.4]
  wire [7:0] _T_15498; // @[Mux.scala 46:16:@11637.4]
  wire  _T_15499; // @[Mux.scala 46:19:@11638.4]
  wire [7:0] _T_15500; // @[Mux.scala 46:16:@11639.4]
  wire  _T_15501; // @[Mux.scala 46:19:@11640.4]
  wire [7:0] _T_15502; // @[Mux.scala 46:16:@11641.4]
  wire  _T_15503; // @[Mux.scala 46:19:@11642.4]
  wire [7:0] _T_15504; // @[Mux.scala 46:16:@11643.4]
  wire  _T_15505; // @[Mux.scala 46:19:@11644.4]
  wire [7:0] _T_15506; // @[Mux.scala 46:16:@11645.4]
  wire  _T_15507; // @[Mux.scala 46:19:@11646.4]
  wire [7:0] _T_15508; // @[Mux.scala 46:16:@11647.4]
  wire  _T_15509; // @[Mux.scala 46:19:@11648.4]
  wire [7:0] _T_15510; // @[Mux.scala 46:16:@11649.4]
  wire  _T_15511; // @[Mux.scala 46:19:@11650.4]
  wire [7:0] _T_15512; // @[Mux.scala 46:16:@11651.4]
  wire  _T_15513; // @[Mux.scala 46:19:@11652.4]
  wire [7:0] _T_15514; // @[Mux.scala 46:16:@11653.4]
  wire  _T_15515; // @[Mux.scala 46:19:@11654.4]
  wire [7:0] _T_15516; // @[Mux.scala 46:16:@11655.4]
  wire  _T_15517; // @[Mux.scala 46:19:@11656.4]
  wire [7:0] _T_15518; // @[Mux.scala 46:16:@11657.4]
  wire  _T_15519; // @[Mux.scala 46:19:@11658.4]
  wire [7:0] _T_15520; // @[Mux.scala 46:16:@11659.4]
  wire  _T_15521; // @[Mux.scala 46:19:@11660.4]
  wire [7:0] _T_15522; // @[Mux.scala 46:16:@11661.4]
  wire  _T_15523; // @[Mux.scala 46:19:@11662.4]
  wire [7:0] _T_15524; // @[Mux.scala 46:16:@11663.4]
  wire  _T_15525; // @[Mux.scala 46:19:@11664.4]
  wire [7:0] _T_15526; // @[Mux.scala 46:16:@11665.4]
  wire  _T_15527; // @[Mux.scala 46:19:@11666.4]
  wire [7:0] _T_15528; // @[Mux.scala 46:16:@11667.4]
  wire  _T_15529; // @[Mux.scala 46:19:@11668.4]
  wire [7:0] _T_15530; // @[Mux.scala 46:16:@11669.4]
  wire  _T_15531; // @[Mux.scala 46:19:@11670.4]
  wire [7:0] _T_15532; // @[Mux.scala 46:16:@11671.4]
  wire  _T_15533; // @[Mux.scala 46:19:@11672.4]
  wire [7:0] _T_15534; // @[Mux.scala 46:16:@11673.4]
  wire  _T_15535; // @[Mux.scala 46:19:@11674.4]
  wire [7:0] _T_15536; // @[Mux.scala 46:16:@11675.4]
  wire  _T_15537; // @[Mux.scala 46:19:@11676.4]
  wire [7:0] _T_15538; // @[Mux.scala 46:16:@11677.4]
  wire  _T_15539; // @[Mux.scala 46:19:@11678.4]
  wire [7:0] _T_15540; // @[Mux.scala 46:16:@11679.4]
  wire  _T_15541; // @[Mux.scala 46:19:@11680.4]
  wire [7:0] _T_15542; // @[Mux.scala 46:16:@11681.4]
  wire  _T_15543; // @[Mux.scala 46:19:@11682.4]
  wire [7:0] _T_15544; // @[Mux.scala 46:16:@11683.4]
  wire  _T_15598; // @[Mux.scala 46:19:@11685.4]
  wire [7:0] _T_15599; // @[Mux.scala 46:16:@11686.4]
  wire  _T_15600; // @[Mux.scala 46:19:@11687.4]
  wire [7:0] _T_15601; // @[Mux.scala 46:16:@11688.4]
  wire  _T_15602; // @[Mux.scala 46:19:@11689.4]
  wire [7:0] _T_15603; // @[Mux.scala 46:16:@11690.4]
  wire  _T_15604; // @[Mux.scala 46:19:@11691.4]
  wire [7:0] _T_15605; // @[Mux.scala 46:16:@11692.4]
  wire  _T_15606; // @[Mux.scala 46:19:@11693.4]
  wire [7:0] _T_15607; // @[Mux.scala 46:16:@11694.4]
  wire  _T_15608; // @[Mux.scala 46:19:@11695.4]
  wire [7:0] _T_15609; // @[Mux.scala 46:16:@11696.4]
  wire  _T_15610; // @[Mux.scala 46:19:@11697.4]
  wire [7:0] _T_15611; // @[Mux.scala 46:16:@11698.4]
  wire  _T_15612; // @[Mux.scala 46:19:@11699.4]
  wire [7:0] _T_15613; // @[Mux.scala 46:16:@11700.4]
  wire  _T_15614; // @[Mux.scala 46:19:@11701.4]
  wire [7:0] _T_15615; // @[Mux.scala 46:16:@11702.4]
  wire  _T_15616; // @[Mux.scala 46:19:@11703.4]
  wire [7:0] _T_15617; // @[Mux.scala 46:16:@11704.4]
  wire  _T_15618; // @[Mux.scala 46:19:@11705.4]
  wire [7:0] _T_15619; // @[Mux.scala 46:16:@11706.4]
  wire  _T_15620; // @[Mux.scala 46:19:@11707.4]
  wire [7:0] _T_15621; // @[Mux.scala 46:16:@11708.4]
  wire  _T_15622; // @[Mux.scala 46:19:@11709.4]
  wire [7:0] _T_15623; // @[Mux.scala 46:16:@11710.4]
  wire  _T_15624; // @[Mux.scala 46:19:@11711.4]
  wire [7:0] _T_15625; // @[Mux.scala 46:16:@11712.4]
  wire  _T_15626; // @[Mux.scala 46:19:@11713.4]
  wire [7:0] _T_15627; // @[Mux.scala 46:16:@11714.4]
  wire  _T_15628; // @[Mux.scala 46:19:@11715.4]
  wire [7:0] _T_15629; // @[Mux.scala 46:16:@11716.4]
  wire  _T_15630; // @[Mux.scala 46:19:@11717.4]
  wire [7:0] _T_15631; // @[Mux.scala 46:16:@11718.4]
  wire  _T_15632; // @[Mux.scala 46:19:@11719.4]
  wire [7:0] _T_15633; // @[Mux.scala 46:16:@11720.4]
  wire  _T_15634; // @[Mux.scala 46:19:@11721.4]
  wire [7:0] _T_15635; // @[Mux.scala 46:16:@11722.4]
  wire  _T_15636; // @[Mux.scala 46:19:@11723.4]
  wire [7:0] _T_15637; // @[Mux.scala 46:16:@11724.4]
  wire  _T_15638; // @[Mux.scala 46:19:@11725.4]
  wire [7:0] _T_15639; // @[Mux.scala 46:16:@11726.4]
  wire  _T_15640; // @[Mux.scala 46:19:@11727.4]
  wire [7:0] _T_15641; // @[Mux.scala 46:16:@11728.4]
  wire  _T_15642; // @[Mux.scala 46:19:@11729.4]
  wire [7:0] _T_15643; // @[Mux.scala 46:16:@11730.4]
  wire  _T_15644; // @[Mux.scala 46:19:@11731.4]
  wire [7:0] _T_15645; // @[Mux.scala 46:16:@11732.4]
  wire  _T_15646; // @[Mux.scala 46:19:@11733.4]
  wire [7:0] _T_15647; // @[Mux.scala 46:16:@11734.4]
  wire  _T_15648; // @[Mux.scala 46:19:@11735.4]
  wire [7:0] _T_15649; // @[Mux.scala 46:16:@11736.4]
  wire  _T_15650; // @[Mux.scala 46:19:@11737.4]
  wire [7:0] _T_15651; // @[Mux.scala 46:16:@11738.4]
  wire  _T_15652; // @[Mux.scala 46:19:@11739.4]
  wire [7:0] _T_15653; // @[Mux.scala 46:16:@11740.4]
  wire  _T_15654; // @[Mux.scala 46:19:@11741.4]
  wire [7:0] _T_15655; // @[Mux.scala 46:16:@11742.4]
  wire  _T_15656; // @[Mux.scala 46:19:@11743.4]
  wire [7:0] _T_15657; // @[Mux.scala 46:16:@11744.4]
  wire  _T_15658; // @[Mux.scala 46:19:@11745.4]
  wire [7:0] _T_15659; // @[Mux.scala 46:16:@11746.4]
  wire  _T_15660; // @[Mux.scala 46:19:@11747.4]
  wire [7:0] _T_15661; // @[Mux.scala 46:16:@11748.4]
  wire  _T_15662; // @[Mux.scala 46:19:@11749.4]
  wire [7:0] _T_15663; // @[Mux.scala 46:16:@11750.4]
  wire  _T_15664; // @[Mux.scala 46:19:@11751.4]
  wire [7:0] _T_15665; // @[Mux.scala 46:16:@11752.4]
  wire  _T_15666; // @[Mux.scala 46:19:@11753.4]
  wire [7:0] _T_15667; // @[Mux.scala 46:16:@11754.4]
  wire  _T_15668; // @[Mux.scala 46:19:@11755.4]
  wire [7:0] _T_15669; // @[Mux.scala 46:16:@11756.4]
  wire  _T_15670; // @[Mux.scala 46:19:@11757.4]
  wire [7:0] _T_15671; // @[Mux.scala 46:16:@11758.4]
  wire  _T_15672; // @[Mux.scala 46:19:@11759.4]
  wire [7:0] _T_15673; // @[Mux.scala 46:16:@11760.4]
  wire  _T_15674; // @[Mux.scala 46:19:@11761.4]
  wire [7:0] _T_15675; // @[Mux.scala 46:16:@11762.4]
  wire  _T_15676; // @[Mux.scala 46:19:@11763.4]
  wire [7:0] _T_15677; // @[Mux.scala 46:16:@11764.4]
  wire  _T_15678; // @[Mux.scala 46:19:@11765.4]
  wire [7:0] _T_15679; // @[Mux.scala 46:16:@11766.4]
  wire  _T_15680; // @[Mux.scala 46:19:@11767.4]
  wire [7:0] _T_15681; // @[Mux.scala 46:16:@11768.4]
  wire  _T_15682; // @[Mux.scala 46:19:@11769.4]
  wire [7:0] _T_15683; // @[Mux.scala 46:16:@11770.4]
  wire  _T_15684; // @[Mux.scala 46:19:@11771.4]
  wire [7:0] _T_15685; // @[Mux.scala 46:16:@11772.4]
  wire  _T_15686; // @[Mux.scala 46:19:@11773.4]
  wire [7:0] _T_15687; // @[Mux.scala 46:16:@11774.4]
  wire  _T_15688; // @[Mux.scala 46:19:@11775.4]
  wire [7:0] _T_15689; // @[Mux.scala 46:16:@11776.4]
  wire  _T_15690; // @[Mux.scala 46:19:@11777.4]
  wire [7:0] _T_15691; // @[Mux.scala 46:16:@11778.4]
  wire  _T_15692; // @[Mux.scala 46:19:@11779.4]
  wire [7:0] _T_15693; // @[Mux.scala 46:16:@11780.4]
  wire  _T_15694; // @[Mux.scala 46:19:@11781.4]
  wire [7:0] _T_15695; // @[Mux.scala 46:16:@11782.4]
  wire  _T_15696; // @[Mux.scala 46:19:@11783.4]
  wire [7:0] _T_15697; // @[Mux.scala 46:16:@11784.4]
  wire  _T_15698; // @[Mux.scala 46:19:@11785.4]
  wire [7:0] _T_15699; // @[Mux.scala 46:16:@11786.4]
  wire  _T_15700; // @[Mux.scala 46:19:@11787.4]
  wire [7:0] _T_15701; // @[Mux.scala 46:16:@11788.4]
  wire  _T_15756; // @[Mux.scala 46:19:@11790.4]
  wire [7:0] _T_15757; // @[Mux.scala 46:16:@11791.4]
  wire  _T_15758; // @[Mux.scala 46:19:@11792.4]
  wire [7:0] _T_15759; // @[Mux.scala 46:16:@11793.4]
  wire  _T_15760; // @[Mux.scala 46:19:@11794.4]
  wire [7:0] _T_15761; // @[Mux.scala 46:16:@11795.4]
  wire  _T_15762; // @[Mux.scala 46:19:@11796.4]
  wire [7:0] _T_15763; // @[Mux.scala 46:16:@11797.4]
  wire  _T_15764; // @[Mux.scala 46:19:@11798.4]
  wire [7:0] _T_15765; // @[Mux.scala 46:16:@11799.4]
  wire  _T_15766; // @[Mux.scala 46:19:@11800.4]
  wire [7:0] _T_15767; // @[Mux.scala 46:16:@11801.4]
  wire  _T_15768; // @[Mux.scala 46:19:@11802.4]
  wire [7:0] _T_15769; // @[Mux.scala 46:16:@11803.4]
  wire  _T_15770; // @[Mux.scala 46:19:@11804.4]
  wire [7:0] _T_15771; // @[Mux.scala 46:16:@11805.4]
  wire  _T_15772; // @[Mux.scala 46:19:@11806.4]
  wire [7:0] _T_15773; // @[Mux.scala 46:16:@11807.4]
  wire  _T_15774; // @[Mux.scala 46:19:@11808.4]
  wire [7:0] _T_15775; // @[Mux.scala 46:16:@11809.4]
  wire  _T_15776; // @[Mux.scala 46:19:@11810.4]
  wire [7:0] _T_15777; // @[Mux.scala 46:16:@11811.4]
  wire  _T_15778; // @[Mux.scala 46:19:@11812.4]
  wire [7:0] _T_15779; // @[Mux.scala 46:16:@11813.4]
  wire  _T_15780; // @[Mux.scala 46:19:@11814.4]
  wire [7:0] _T_15781; // @[Mux.scala 46:16:@11815.4]
  wire  _T_15782; // @[Mux.scala 46:19:@11816.4]
  wire [7:0] _T_15783; // @[Mux.scala 46:16:@11817.4]
  wire  _T_15784; // @[Mux.scala 46:19:@11818.4]
  wire [7:0] _T_15785; // @[Mux.scala 46:16:@11819.4]
  wire  _T_15786; // @[Mux.scala 46:19:@11820.4]
  wire [7:0] _T_15787; // @[Mux.scala 46:16:@11821.4]
  wire  _T_15788; // @[Mux.scala 46:19:@11822.4]
  wire [7:0] _T_15789; // @[Mux.scala 46:16:@11823.4]
  wire  _T_15790; // @[Mux.scala 46:19:@11824.4]
  wire [7:0] _T_15791; // @[Mux.scala 46:16:@11825.4]
  wire  _T_15792; // @[Mux.scala 46:19:@11826.4]
  wire [7:0] _T_15793; // @[Mux.scala 46:16:@11827.4]
  wire  _T_15794; // @[Mux.scala 46:19:@11828.4]
  wire [7:0] _T_15795; // @[Mux.scala 46:16:@11829.4]
  wire  _T_15796; // @[Mux.scala 46:19:@11830.4]
  wire [7:0] _T_15797; // @[Mux.scala 46:16:@11831.4]
  wire  _T_15798; // @[Mux.scala 46:19:@11832.4]
  wire [7:0] _T_15799; // @[Mux.scala 46:16:@11833.4]
  wire  _T_15800; // @[Mux.scala 46:19:@11834.4]
  wire [7:0] _T_15801; // @[Mux.scala 46:16:@11835.4]
  wire  _T_15802; // @[Mux.scala 46:19:@11836.4]
  wire [7:0] _T_15803; // @[Mux.scala 46:16:@11837.4]
  wire  _T_15804; // @[Mux.scala 46:19:@11838.4]
  wire [7:0] _T_15805; // @[Mux.scala 46:16:@11839.4]
  wire  _T_15806; // @[Mux.scala 46:19:@11840.4]
  wire [7:0] _T_15807; // @[Mux.scala 46:16:@11841.4]
  wire  _T_15808; // @[Mux.scala 46:19:@11842.4]
  wire [7:0] _T_15809; // @[Mux.scala 46:16:@11843.4]
  wire  _T_15810; // @[Mux.scala 46:19:@11844.4]
  wire [7:0] _T_15811; // @[Mux.scala 46:16:@11845.4]
  wire  _T_15812; // @[Mux.scala 46:19:@11846.4]
  wire [7:0] _T_15813; // @[Mux.scala 46:16:@11847.4]
  wire  _T_15814; // @[Mux.scala 46:19:@11848.4]
  wire [7:0] _T_15815; // @[Mux.scala 46:16:@11849.4]
  wire  _T_15816; // @[Mux.scala 46:19:@11850.4]
  wire [7:0] _T_15817; // @[Mux.scala 46:16:@11851.4]
  wire  _T_15818; // @[Mux.scala 46:19:@11852.4]
  wire [7:0] _T_15819; // @[Mux.scala 46:16:@11853.4]
  wire  _T_15820; // @[Mux.scala 46:19:@11854.4]
  wire [7:0] _T_15821; // @[Mux.scala 46:16:@11855.4]
  wire  _T_15822; // @[Mux.scala 46:19:@11856.4]
  wire [7:0] _T_15823; // @[Mux.scala 46:16:@11857.4]
  wire  _T_15824; // @[Mux.scala 46:19:@11858.4]
  wire [7:0] _T_15825; // @[Mux.scala 46:16:@11859.4]
  wire  _T_15826; // @[Mux.scala 46:19:@11860.4]
  wire [7:0] _T_15827; // @[Mux.scala 46:16:@11861.4]
  wire  _T_15828; // @[Mux.scala 46:19:@11862.4]
  wire [7:0] _T_15829; // @[Mux.scala 46:16:@11863.4]
  wire  _T_15830; // @[Mux.scala 46:19:@11864.4]
  wire [7:0] _T_15831; // @[Mux.scala 46:16:@11865.4]
  wire  _T_15832; // @[Mux.scala 46:19:@11866.4]
  wire [7:0] _T_15833; // @[Mux.scala 46:16:@11867.4]
  wire  _T_15834; // @[Mux.scala 46:19:@11868.4]
  wire [7:0] _T_15835; // @[Mux.scala 46:16:@11869.4]
  wire  _T_15836; // @[Mux.scala 46:19:@11870.4]
  wire [7:0] _T_15837; // @[Mux.scala 46:16:@11871.4]
  wire  _T_15838; // @[Mux.scala 46:19:@11872.4]
  wire [7:0] _T_15839; // @[Mux.scala 46:16:@11873.4]
  wire  _T_15840; // @[Mux.scala 46:19:@11874.4]
  wire [7:0] _T_15841; // @[Mux.scala 46:16:@11875.4]
  wire  _T_15842; // @[Mux.scala 46:19:@11876.4]
  wire [7:0] _T_15843; // @[Mux.scala 46:16:@11877.4]
  wire  _T_15844; // @[Mux.scala 46:19:@11878.4]
  wire [7:0] _T_15845; // @[Mux.scala 46:16:@11879.4]
  wire  _T_15846; // @[Mux.scala 46:19:@11880.4]
  wire [7:0] _T_15847; // @[Mux.scala 46:16:@11881.4]
  wire  _T_15848; // @[Mux.scala 46:19:@11882.4]
  wire [7:0] _T_15849; // @[Mux.scala 46:16:@11883.4]
  wire  _T_15850; // @[Mux.scala 46:19:@11884.4]
  wire [7:0] _T_15851; // @[Mux.scala 46:16:@11885.4]
  wire  _T_15852; // @[Mux.scala 46:19:@11886.4]
  wire [7:0] _T_15853; // @[Mux.scala 46:16:@11887.4]
  wire  _T_15854; // @[Mux.scala 46:19:@11888.4]
  wire [7:0] _T_15855; // @[Mux.scala 46:16:@11889.4]
  wire  _T_15856; // @[Mux.scala 46:19:@11890.4]
  wire [7:0] _T_15857; // @[Mux.scala 46:16:@11891.4]
  wire  _T_15858; // @[Mux.scala 46:19:@11892.4]
  wire [7:0] _T_15859; // @[Mux.scala 46:16:@11893.4]
  wire  _T_15860; // @[Mux.scala 46:19:@11894.4]
  wire [7:0] _T_15861; // @[Mux.scala 46:16:@11895.4]
  wire  _T_15917; // @[Mux.scala 46:19:@11897.4]
  wire [7:0] _T_15918; // @[Mux.scala 46:16:@11898.4]
  wire  _T_15919; // @[Mux.scala 46:19:@11899.4]
  wire [7:0] _T_15920; // @[Mux.scala 46:16:@11900.4]
  wire  _T_15921; // @[Mux.scala 46:19:@11901.4]
  wire [7:0] _T_15922; // @[Mux.scala 46:16:@11902.4]
  wire  _T_15923; // @[Mux.scala 46:19:@11903.4]
  wire [7:0] _T_15924; // @[Mux.scala 46:16:@11904.4]
  wire  _T_15925; // @[Mux.scala 46:19:@11905.4]
  wire [7:0] _T_15926; // @[Mux.scala 46:16:@11906.4]
  wire  _T_15927; // @[Mux.scala 46:19:@11907.4]
  wire [7:0] _T_15928; // @[Mux.scala 46:16:@11908.4]
  wire  _T_15929; // @[Mux.scala 46:19:@11909.4]
  wire [7:0] _T_15930; // @[Mux.scala 46:16:@11910.4]
  wire  _T_15931; // @[Mux.scala 46:19:@11911.4]
  wire [7:0] _T_15932; // @[Mux.scala 46:16:@11912.4]
  wire  _T_15933; // @[Mux.scala 46:19:@11913.4]
  wire [7:0] _T_15934; // @[Mux.scala 46:16:@11914.4]
  wire  _T_15935; // @[Mux.scala 46:19:@11915.4]
  wire [7:0] _T_15936; // @[Mux.scala 46:16:@11916.4]
  wire  _T_15937; // @[Mux.scala 46:19:@11917.4]
  wire [7:0] _T_15938; // @[Mux.scala 46:16:@11918.4]
  wire  _T_15939; // @[Mux.scala 46:19:@11919.4]
  wire [7:0] _T_15940; // @[Mux.scala 46:16:@11920.4]
  wire  _T_15941; // @[Mux.scala 46:19:@11921.4]
  wire [7:0] _T_15942; // @[Mux.scala 46:16:@11922.4]
  wire  _T_15943; // @[Mux.scala 46:19:@11923.4]
  wire [7:0] _T_15944; // @[Mux.scala 46:16:@11924.4]
  wire  _T_15945; // @[Mux.scala 46:19:@11925.4]
  wire [7:0] _T_15946; // @[Mux.scala 46:16:@11926.4]
  wire  _T_15947; // @[Mux.scala 46:19:@11927.4]
  wire [7:0] _T_15948; // @[Mux.scala 46:16:@11928.4]
  wire  _T_15949; // @[Mux.scala 46:19:@11929.4]
  wire [7:0] _T_15950; // @[Mux.scala 46:16:@11930.4]
  wire  _T_15951; // @[Mux.scala 46:19:@11931.4]
  wire [7:0] _T_15952; // @[Mux.scala 46:16:@11932.4]
  wire  _T_15953; // @[Mux.scala 46:19:@11933.4]
  wire [7:0] _T_15954; // @[Mux.scala 46:16:@11934.4]
  wire  _T_15955; // @[Mux.scala 46:19:@11935.4]
  wire [7:0] _T_15956; // @[Mux.scala 46:16:@11936.4]
  wire  _T_15957; // @[Mux.scala 46:19:@11937.4]
  wire [7:0] _T_15958; // @[Mux.scala 46:16:@11938.4]
  wire  _T_15959; // @[Mux.scala 46:19:@11939.4]
  wire [7:0] _T_15960; // @[Mux.scala 46:16:@11940.4]
  wire  _T_15961; // @[Mux.scala 46:19:@11941.4]
  wire [7:0] _T_15962; // @[Mux.scala 46:16:@11942.4]
  wire  _T_15963; // @[Mux.scala 46:19:@11943.4]
  wire [7:0] _T_15964; // @[Mux.scala 46:16:@11944.4]
  wire  _T_15965; // @[Mux.scala 46:19:@11945.4]
  wire [7:0] _T_15966; // @[Mux.scala 46:16:@11946.4]
  wire  _T_15967; // @[Mux.scala 46:19:@11947.4]
  wire [7:0] _T_15968; // @[Mux.scala 46:16:@11948.4]
  wire  _T_15969; // @[Mux.scala 46:19:@11949.4]
  wire [7:0] _T_15970; // @[Mux.scala 46:16:@11950.4]
  wire  _T_15971; // @[Mux.scala 46:19:@11951.4]
  wire [7:0] _T_15972; // @[Mux.scala 46:16:@11952.4]
  wire  _T_15973; // @[Mux.scala 46:19:@11953.4]
  wire [7:0] _T_15974; // @[Mux.scala 46:16:@11954.4]
  wire  _T_15975; // @[Mux.scala 46:19:@11955.4]
  wire [7:0] _T_15976; // @[Mux.scala 46:16:@11956.4]
  wire  _T_15977; // @[Mux.scala 46:19:@11957.4]
  wire [7:0] _T_15978; // @[Mux.scala 46:16:@11958.4]
  wire  _T_15979; // @[Mux.scala 46:19:@11959.4]
  wire [7:0] _T_15980; // @[Mux.scala 46:16:@11960.4]
  wire  _T_15981; // @[Mux.scala 46:19:@11961.4]
  wire [7:0] _T_15982; // @[Mux.scala 46:16:@11962.4]
  wire  _T_15983; // @[Mux.scala 46:19:@11963.4]
  wire [7:0] _T_15984; // @[Mux.scala 46:16:@11964.4]
  wire  _T_15985; // @[Mux.scala 46:19:@11965.4]
  wire [7:0] _T_15986; // @[Mux.scala 46:16:@11966.4]
  wire  _T_15987; // @[Mux.scala 46:19:@11967.4]
  wire [7:0] _T_15988; // @[Mux.scala 46:16:@11968.4]
  wire  _T_15989; // @[Mux.scala 46:19:@11969.4]
  wire [7:0] _T_15990; // @[Mux.scala 46:16:@11970.4]
  wire  _T_15991; // @[Mux.scala 46:19:@11971.4]
  wire [7:0] _T_15992; // @[Mux.scala 46:16:@11972.4]
  wire  _T_15993; // @[Mux.scala 46:19:@11973.4]
  wire [7:0] _T_15994; // @[Mux.scala 46:16:@11974.4]
  wire  _T_15995; // @[Mux.scala 46:19:@11975.4]
  wire [7:0] _T_15996; // @[Mux.scala 46:16:@11976.4]
  wire  _T_15997; // @[Mux.scala 46:19:@11977.4]
  wire [7:0] _T_15998; // @[Mux.scala 46:16:@11978.4]
  wire  _T_15999; // @[Mux.scala 46:19:@11979.4]
  wire [7:0] _T_16000; // @[Mux.scala 46:16:@11980.4]
  wire  _T_16001; // @[Mux.scala 46:19:@11981.4]
  wire [7:0] _T_16002; // @[Mux.scala 46:16:@11982.4]
  wire  _T_16003; // @[Mux.scala 46:19:@11983.4]
  wire [7:0] _T_16004; // @[Mux.scala 46:16:@11984.4]
  wire  _T_16005; // @[Mux.scala 46:19:@11985.4]
  wire [7:0] _T_16006; // @[Mux.scala 46:16:@11986.4]
  wire  _T_16007; // @[Mux.scala 46:19:@11987.4]
  wire [7:0] _T_16008; // @[Mux.scala 46:16:@11988.4]
  wire  _T_16009; // @[Mux.scala 46:19:@11989.4]
  wire [7:0] _T_16010; // @[Mux.scala 46:16:@11990.4]
  wire  _T_16011; // @[Mux.scala 46:19:@11991.4]
  wire [7:0] _T_16012; // @[Mux.scala 46:16:@11992.4]
  wire  _T_16013; // @[Mux.scala 46:19:@11993.4]
  wire [7:0] _T_16014; // @[Mux.scala 46:16:@11994.4]
  wire  _T_16015; // @[Mux.scala 46:19:@11995.4]
  wire [7:0] _T_16016; // @[Mux.scala 46:16:@11996.4]
  wire  _T_16017; // @[Mux.scala 46:19:@11997.4]
  wire [7:0] _T_16018; // @[Mux.scala 46:16:@11998.4]
  wire  _T_16019; // @[Mux.scala 46:19:@11999.4]
  wire [7:0] _T_16020; // @[Mux.scala 46:16:@12000.4]
  wire  _T_16021; // @[Mux.scala 46:19:@12001.4]
  wire [7:0] _T_16022; // @[Mux.scala 46:16:@12002.4]
  wire  _T_16023; // @[Mux.scala 46:19:@12003.4]
  wire [7:0] _T_16024; // @[Mux.scala 46:16:@12004.4]
  wire  _T_16081; // @[Mux.scala 46:19:@12006.4]
  wire [7:0] _T_16082; // @[Mux.scala 46:16:@12007.4]
  wire  _T_16083; // @[Mux.scala 46:19:@12008.4]
  wire [7:0] _T_16084; // @[Mux.scala 46:16:@12009.4]
  wire  _T_16085; // @[Mux.scala 46:19:@12010.4]
  wire [7:0] _T_16086; // @[Mux.scala 46:16:@12011.4]
  wire  _T_16087; // @[Mux.scala 46:19:@12012.4]
  wire [7:0] _T_16088; // @[Mux.scala 46:16:@12013.4]
  wire  _T_16089; // @[Mux.scala 46:19:@12014.4]
  wire [7:0] _T_16090; // @[Mux.scala 46:16:@12015.4]
  wire  _T_16091; // @[Mux.scala 46:19:@12016.4]
  wire [7:0] _T_16092; // @[Mux.scala 46:16:@12017.4]
  wire  _T_16093; // @[Mux.scala 46:19:@12018.4]
  wire [7:0] _T_16094; // @[Mux.scala 46:16:@12019.4]
  wire  _T_16095; // @[Mux.scala 46:19:@12020.4]
  wire [7:0] _T_16096; // @[Mux.scala 46:16:@12021.4]
  wire  _T_16097; // @[Mux.scala 46:19:@12022.4]
  wire [7:0] _T_16098; // @[Mux.scala 46:16:@12023.4]
  wire  _T_16099; // @[Mux.scala 46:19:@12024.4]
  wire [7:0] _T_16100; // @[Mux.scala 46:16:@12025.4]
  wire  _T_16101; // @[Mux.scala 46:19:@12026.4]
  wire [7:0] _T_16102; // @[Mux.scala 46:16:@12027.4]
  wire  _T_16103; // @[Mux.scala 46:19:@12028.4]
  wire [7:0] _T_16104; // @[Mux.scala 46:16:@12029.4]
  wire  _T_16105; // @[Mux.scala 46:19:@12030.4]
  wire [7:0] _T_16106; // @[Mux.scala 46:16:@12031.4]
  wire  _T_16107; // @[Mux.scala 46:19:@12032.4]
  wire [7:0] _T_16108; // @[Mux.scala 46:16:@12033.4]
  wire  _T_16109; // @[Mux.scala 46:19:@12034.4]
  wire [7:0] _T_16110; // @[Mux.scala 46:16:@12035.4]
  wire  _T_16111; // @[Mux.scala 46:19:@12036.4]
  wire [7:0] _T_16112; // @[Mux.scala 46:16:@12037.4]
  wire  _T_16113; // @[Mux.scala 46:19:@12038.4]
  wire [7:0] _T_16114; // @[Mux.scala 46:16:@12039.4]
  wire  _T_16115; // @[Mux.scala 46:19:@12040.4]
  wire [7:0] _T_16116; // @[Mux.scala 46:16:@12041.4]
  wire  _T_16117; // @[Mux.scala 46:19:@12042.4]
  wire [7:0] _T_16118; // @[Mux.scala 46:16:@12043.4]
  wire  _T_16119; // @[Mux.scala 46:19:@12044.4]
  wire [7:0] _T_16120; // @[Mux.scala 46:16:@12045.4]
  wire  _T_16121; // @[Mux.scala 46:19:@12046.4]
  wire [7:0] _T_16122; // @[Mux.scala 46:16:@12047.4]
  wire  _T_16123; // @[Mux.scala 46:19:@12048.4]
  wire [7:0] _T_16124; // @[Mux.scala 46:16:@12049.4]
  wire  _T_16125; // @[Mux.scala 46:19:@12050.4]
  wire [7:0] _T_16126; // @[Mux.scala 46:16:@12051.4]
  wire  _T_16127; // @[Mux.scala 46:19:@12052.4]
  wire [7:0] _T_16128; // @[Mux.scala 46:16:@12053.4]
  wire  _T_16129; // @[Mux.scala 46:19:@12054.4]
  wire [7:0] _T_16130; // @[Mux.scala 46:16:@12055.4]
  wire  _T_16131; // @[Mux.scala 46:19:@12056.4]
  wire [7:0] _T_16132; // @[Mux.scala 46:16:@12057.4]
  wire  _T_16133; // @[Mux.scala 46:19:@12058.4]
  wire [7:0] _T_16134; // @[Mux.scala 46:16:@12059.4]
  wire  _T_16135; // @[Mux.scala 46:19:@12060.4]
  wire [7:0] _T_16136; // @[Mux.scala 46:16:@12061.4]
  wire  _T_16137; // @[Mux.scala 46:19:@12062.4]
  wire [7:0] _T_16138; // @[Mux.scala 46:16:@12063.4]
  wire  _T_16139; // @[Mux.scala 46:19:@12064.4]
  wire [7:0] _T_16140; // @[Mux.scala 46:16:@12065.4]
  wire  _T_16141; // @[Mux.scala 46:19:@12066.4]
  wire [7:0] _T_16142; // @[Mux.scala 46:16:@12067.4]
  wire  _T_16143; // @[Mux.scala 46:19:@12068.4]
  wire [7:0] _T_16144; // @[Mux.scala 46:16:@12069.4]
  wire  _T_16145; // @[Mux.scala 46:19:@12070.4]
  wire [7:0] _T_16146; // @[Mux.scala 46:16:@12071.4]
  wire  _T_16147; // @[Mux.scala 46:19:@12072.4]
  wire [7:0] _T_16148; // @[Mux.scala 46:16:@12073.4]
  wire  _T_16149; // @[Mux.scala 46:19:@12074.4]
  wire [7:0] _T_16150; // @[Mux.scala 46:16:@12075.4]
  wire  _T_16151; // @[Mux.scala 46:19:@12076.4]
  wire [7:0] _T_16152; // @[Mux.scala 46:16:@12077.4]
  wire  _T_16153; // @[Mux.scala 46:19:@12078.4]
  wire [7:0] _T_16154; // @[Mux.scala 46:16:@12079.4]
  wire  _T_16155; // @[Mux.scala 46:19:@12080.4]
  wire [7:0] _T_16156; // @[Mux.scala 46:16:@12081.4]
  wire  _T_16157; // @[Mux.scala 46:19:@12082.4]
  wire [7:0] _T_16158; // @[Mux.scala 46:16:@12083.4]
  wire  _T_16159; // @[Mux.scala 46:19:@12084.4]
  wire [7:0] _T_16160; // @[Mux.scala 46:16:@12085.4]
  wire  _T_16161; // @[Mux.scala 46:19:@12086.4]
  wire [7:0] _T_16162; // @[Mux.scala 46:16:@12087.4]
  wire  _T_16163; // @[Mux.scala 46:19:@12088.4]
  wire [7:0] _T_16164; // @[Mux.scala 46:16:@12089.4]
  wire  _T_16165; // @[Mux.scala 46:19:@12090.4]
  wire [7:0] _T_16166; // @[Mux.scala 46:16:@12091.4]
  wire  _T_16167; // @[Mux.scala 46:19:@12092.4]
  wire [7:0] _T_16168; // @[Mux.scala 46:16:@12093.4]
  wire  _T_16169; // @[Mux.scala 46:19:@12094.4]
  wire [7:0] _T_16170; // @[Mux.scala 46:16:@12095.4]
  wire  _T_16171; // @[Mux.scala 46:19:@12096.4]
  wire [7:0] _T_16172; // @[Mux.scala 46:16:@12097.4]
  wire  _T_16173; // @[Mux.scala 46:19:@12098.4]
  wire [7:0] _T_16174; // @[Mux.scala 46:16:@12099.4]
  wire  _T_16175; // @[Mux.scala 46:19:@12100.4]
  wire [7:0] _T_16176; // @[Mux.scala 46:16:@12101.4]
  wire  _T_16177; // @[Mux.scala 46:19:@12102.4]
  wire [7:0] _T_16178; // @[Mux.scala 46:16:@12103.4]
  wire  _T_16179; // @[Mux.scala 46:19:@12104.4]
  wire [7:0] _T_16180; // @[Mux.scala 46:16:@12105.4]
  wire  _T_16181; // @[Mux.scala 46:19:@12106.4]
  wire [7:0] _T_16182; // @[Mux.scala 46:16:@12107.4]
  wire  _T_16183; // @[Mux.scala 46:19:@12108.4]
  wire [7:0] _T_16184; // @[Mux.scala 46:16:@12109.4]
  wire  _T_16185; // @[Mux.scala 46:19:@12110.4]
  wire [7:0] _T_16186; // @[Mux.scala 46:16:@12111.4]
  wire  _T_16187; // @[Mux.scala 46:19:@12112.4]
  wire [7:0] _T_16188; // @[Mux.scala 46:16:@12113.4]
  wire  _T_16189; // @[Mux.scala 46:19:@12114.4]
  wire [7:0] _T_16190; // @[Mux.scala 46:16:@12115.4]
  wire  _T_16248; // @[Mux.scala 46:19:@12117.4]
  wire [7:0] _T_16249; // @[Mux.scala 46:16:@12118.4]
  wire  _T_16250; // @[Mux.scala 46:19:@12119.4]
  wire [7:0] _T_16251; // @[Mux.scala 46:16:@12120.4]
  wire  _T_16252; // @[Mux.scala 46:19:@12121.4]
  wire [7:0] _T_16253; // @[Mux.scala 46:16:@12122.4]
  wire  _T_16254; // @[Mux.scala 46:19:@12123.4]
  wire [7:0] _T_16255; // @[Mux.scala 46:16:@12124.4]
  wire  _T_16256; // @[Mux.scala 46:19:@12125.4]
  wire [7:0] _T_16257; // @[Mux.scala 46:16:@12126.4]
  wire  _T_16258; // @[Mux.scala 46:19:@12127.4]
  wire [7:0] _T_16259; // @[Mux.scala 46:16:@12128.4]
  wire  _T_16260; // @[Mux.scala 46:19:@12129.4]
  wire [7:0] _T_16261; // @[Mux.scala 46:16:@12130.4]
  wire  _T_16262; // @[Mux.scala 46:19:@12131.4]
  wire [7:0] _T_16263; // @[Mux.scala 46:16:@12132.4]
  wire  _T_16264; // @[Mux.scala 46:19:@12133.4]
  wire [7:0] _T_16265; // @[Mux.scala 46:16:@12134.4]
  wire  _T_16266; // @[Mux.scala 46:19:@12135.4]
  wire [7:0] _T_16267; // @[Mux.scala 46:16:@12136.4]
  wire  _T_16268; // @[Mux.scala 46:19:@12137.4]
  wire [7:0] _T_16269; // @[Mux.scala 46:16:@12138.4]
  wire  _T_16270; // @[Mux.scala 46:19:@12139.4]
  wire [7:0] _T_16271; // @[Mux.scala 46:16:@12140.4]
  wire  _T_16272; // @[Mux.scala 46:19:@12141.4]
  wire [7:0] _T_16273; // @[Mux.scala 46:16:@12142.4]
  wire  _T_16274; // @[Mux.scala 46:19:@12143.4]
  wire [7:0] _T_16275; // @[Mux.scala 46:16:@12144.4]
  wire  _T_16276; // @[Mux.scala 46:19:@12145.4]
  wire [7:0] _T_16277; // @[Mux.scala 46:16:@12146.4]
  wire  _T_16278; // @[Mux.scala 46:19:@12147.4]
  wire [7:0] _T_16279; // @[Mux.scala 46:16:@12148.4]
  wire  _T_16280; // @[Mux.scala 46:19:@12149.4]
  wire [7:0] _T_16281; // @[Mux.scala 46:16:@12150.4]
  wire  _T_16282; // @[Mux.scala 46:19:@12151.4]
  wire [7:0] _T_16283; // @[Mux.scala 46:16:@12152.4]
  wire  _T_16284; // @[Mux.scala 46:19:@12153.4]
  wire [7:0] _T_16285; // @[Mux.scala 46:16:@12154.4]
  wire  _T_16286; // @[Mux.scala 46:19:@12155.4]
  wire [7:0] _T_16287; // @[Mux.scala 46:16:@12156.4]
  wire  _T_16288; // @[Mux.scala 46:19:@12157.4]
  wire [7:0] _T_16289; // @[Mux.scala 46:16:@12158.4]
  wire  _T_16290; // @[Mux.scala 46:19:@12159.4]
  wire [7:0] _T_16291; // @[Mux.scala 46:16:@12160.4]
  wire  _T_16292; // @[Mux.scala 46:19:@12161.4]
  wire [7:0] _T_16293; // @[Mux.scala 46:16:@12162.4]
  wire  _T_16294; // @[Mux.scala 46:19:@12163.4]
  wire [7:0] _T_16295; // @[Mux.scala 46:16:@12164.4]
  wire  _T_16296; // @[Mux.scala 46:19:@12165.4]
  wire [7:0] _T_16297; // @[Mux.scala 46:16:@12166.4]
  wire  _T_16298; // @[Mux.scala 46:19:@12167.4]
  wire [7:0] _T_16299; // @[Mux.scala 46:16:@12168.4]
  wire  _T_16300; // @[Mux.scala 46:19:@12169.4]
  wire [7:0] _T_16301; // @[Mux.scala 46:16:@12170.4]
  wire  _T_16302; // @[Mux.scala 46:19:@12171.4]
  wire [7:0] _T_16303; // @[Mux.scala 46:16:@12172.4]
  wire  _T_16304; // @[Mux.scala 46:19:@12173.4]
  wire [7:0] _T_16305; // @[Mux.scala 46:16:@12174.4]
  wire  _T_16306; // @[Mux.scala 46:19:@12175.4]
  wire [7:0] _T_16307; // @[Mux.scala 46:16:@12176.4]
  wire  _T_16308; // @[Mux.scala 46:19:@12177.4]
  wire [7:0] _T_16309; // @[Mux.scala 46:16:@12178.4]
  wire  _T_16310; // @[Mux.scala 46:19:@12179.4]
  wire [7:0] _T_16311; // @[Mux.scala 46:16:@12180.4]
  wire  _T_16312; // @[Mux.scala 46:19:@12181.4]
  wire [7:0] _T_16313; // @[Mux.scala 46:16:@12182.4]
  wire  _T_16314; // @[Mux.scala 46:19:@12183.4]
  wire [7:0] _T_16315; // @[Mux.scala 46:16:@12184.4]
  wire  _T_16316; // @[Mux.scala 46:19:@12185.4]
  wire [7:0] _T_16317; // @[Mux.scala 46:16:@12186.4]
  wire  _T_16318; // @[Mux.scala 46:19:@12187.4]
  wire [7:0] _T_16319; // @[Mux.scala 46:16:@12188.4]
  wire  _T_16320; // @[Mux.scala 46:19:@12189.4]
  wire [7:0] _T_16321; // @[Mux.scala 46:16:@12190.4]
  wire  _T_16322; // @[Mux.scala 46:19:@12191.4]
  wire [7:0] _T_16323; // @[Mux.scala 46:16:@12192.4]
  wire  _T_16324; // @[Mux.scala 46:19:@12193.4]
  wire [7:0] _T_16325; // @[Mux.scala 46:16:@12194.4]
  wire  _T_16326; // @[Mux.scala 46:19:@12195.4]
  wire [7:0] _T_16327; // @[Mux.scala 46:16:@12196.4]
  wire  _T_16328; // @[Mux.scala 46:19:@12197.4]
  wire [7:0] _T_16329; // @[Mux.scala 46:16:@12198.4]
  wire  _T_16330; // @[Mux.scala 46:19:@12199.4]
  wire [7:0] _T_16331; // @[Mux.scala 46:16:@12200.4]
  wire  _T_16332; // @[Mux.scala 46:19:@12201.4]
  wire [7:0] _T_16333; // @[Mux.scala 46:16:@12202.4]
  wire  _T_16334; // @[Mux.scala 46:19:@12203.4]
  wire [7:0] _T_16335; // @[Mux.scala 46:16:@12204.4]
  wire  _T_16336; // @[Mux.scala 46:19:@12205.4]
  wire [7:0] _T_16337; // @[Mux.scala 46:16:@12206.4]
  wire  _T_16338; // @[Mux.scala 46:19:@12207.4]
  wire [7:0] _T_16339; // @[Mux.scala 46:16:@12208.4]
  wire  _T_16340; // @[Mux.scala 46:19:@12209.4]
  wire [7:0] _T_16341; // @[Mux.scala 46:16:@12210.4]
  wire  _T_16342; // @[Mux.scala 46:19:@12211.4]
  wire [7:0] _T_16343; // @[Mux.scala 46:16:@12212.4]
  wire  _T_16344; // @[Mux.scala 46:19:@12213.4]
  wire [7:0] _T_16345; // @[Mux.scala 46:16:@12214.4]
  wire  _T_16346; // @[Mux.scala 46:19:@12215.4]
  wire [7:0] _T_16347; // @[Mux.scala 46:16:@12216.4]
  wire  _T_16348; // @[Mux.scala 46:19:@12217.4]
  wire [7:0] _T_16349; // @[Mux.scala 46:16:@12218.4]
  wire  _T_16350; // @[Mux.scala 46:19:@12219.4]
  wire [7:0] _T_16351; // @[Mux.scala 46:16:@12220.4]
  wire  _T_16352; // @[Mux.scala 46:19:@12221.4]
  wire [7:0] _T_16353; // @[Mux.scala 46:16:@12222.4]
  wire  _T_16354; // @[Mux.scala 46:19:@12223.4]
  wire [7:0] _T_16355; // @[Mux.scala 46:16:@12224.4]
  wire  _T_16356; // @[Mux.scala 46:19:@12225.4]
  wire [7:0] _T_16357; // @[Mux.scala 46:16:@12226.4]
  wire  _T_16358; // @[Mux.scala 46:19:@12227.4]
  wire [7:0] _T_16359; // @[Mux.scala 46:16:@12228.4]
  wire  _T_16418; // @[Mux.scala 46:19:@12230.4]
  wire [7:0] _T_16419; // @[Mux.scala 46:16:@12231.4]
  wire  _T_16420; // @[Mux.scala 46:19:@12232.4]
  wire [7:0] _T_16421; // @[Mux.scala 46:16:@12233.4]
  wire  _T_16422; // @[Mux.scala 46:19:@12234.4]
  wire [7:0] _T_16423; // @[Mux.scala 46:16:@12235.4]
  wire  _T_16424; // @[Mux.scala 46:19:@12236.4]
  wire [7:0] _T_16425; // @[Mux.scala 46:16:@12237.4]
  wire  _T_16426; // @[Mux.scala 46:19:@12238.4]
  wire [7:0] _T_16427; // @[Mux.scala 46:16:@12239.4]
  wire  _T_16428; // @[Mux.scala 46:19:@12240.4]
  wire [7:0] _T_16429; // @[Mux.scala 46:16:@12241.4]
  wire  _T_16430; // @[Mux.scala 46:19:@12242.4]
  wire [7:0] _T_16431; // @[Mux.scala 46:16:@12243.4]
  wire  _T_16432; // @[Mux.scala 46:19:@12244.4]
  wire [7:0] _T_16433; // @[Mux.scala 46:16:@12245.4]
  wire  _T_16434; // @[Mux.scala 46:19:@12246.4]
  wire [7:0] _T_16435; // @[Mux.scala 46:16:@12247.4]
  wire  _T_16436; // @[Mux.scala 46:19:@12248.4]
  wire [7:0] _T_16437; // @[Mux.scala 46:16:@12249.4]
  wire  _T_16438; // @[Mux.scala 46:19:@12250.4]
  wire [7:0] _T_16439; // @[Mux.scala 46:16:@12251.4]
  wire  _T_16440; // @[Mux.scala 46:19:@12252.4]
  wire [7:0] _T_16441; // @[Mux.scala 46:16:@12253.4]
  wire  _T_16442; // @[Mux.scala 46:19:@12254.4]
  wire [7:0] _T_16443; // @[Mux.scala 46:16:@12255.4]
  wire  _T_16444; // @[Mux.scala 46:19:@12256.4]
  wire [7:0] _T_16445; // @[Mux.scala 46:16:@12257.4]
  wire  _T_16446; // @[Mux.scala 46:19:@12258.4]
  wire [7:0] _T_16447; // @[Mux.scala 46:16:@12259.4]
  wire  _T_16448; // @[Mux.scala 46:19:@12260.4]
  wire [7:0] _T_16449; // @[Mux.scala 46:16:@12261.4]
  wire  _T_16450; // @[Mux.scala 46:19:@12262.4]
  wire [7:0] _T_16451; // @[Mux.scala 46:16:@12263.4]
  wire  _T_16452; // @[Mux.scala 46:19:@12264.4]
  wire [7:0] _T_16453; // @[Mux.scala 46:16:@12265.4]
  wire  _T_16454; // @[Mux.scala 46:19:@12266.4]
  wire [7:0] _T_16455; // @[Mux.scala 46:16:@12267.4]
  wire  _T_16456; // @[Mux.scala 46:19:@12268.4]
  wire [7:0] _T_16457; // @[Mux.scala 46:16:@12269.4]
  wire  _T_16458; // @[Mux.scala 46:19:@12270.4]
  wire [7:0] _T_16459; // @[Mux.scala 46:16:@12271.4]
  wire  _T_16460; // @[Mux.scala 46:19:@12272.4]
  wire [7:0] _T_16461; // @[Mux.scala 46:16:@12273.4]
  wire  _T_16462; // @[Mux.scala 46:19:@12274.4]
  wire [7:0] _T_16463; // @[Mux.scala 46:16:@12275.4]
  wire  _T_16464; // @[Mux.scala 46:19:@12276.4]
  wire [7:0] _T_16465; // @[Mux.scala 46:16:@12277.4]
  wire  _T_16466; // @[Mux.scala 46:19:@12278.4]
  wire [7:0] _T_16467; // @[Mux.scala 46:16:@12279.4]
  wire  _T_16468; // @[Mux.scala 46:19:@12280.4]
  wire [7:0] _T_16469; // @[Mux.scala 46:16:@12281.4]
  wire  _T_16470; // @[Mux.scala 46:19:@12282.4]
  wire [7:0] _T_16471; // @[Mux.scala 46:16:@12283.4]
  wire  _T_16472; // @[Mux.scala 46:19:@12284.4]
  wire [7:0] _T_16473; // @[Mux.scala 46:16:@12285.4]
  wire  _T_16474; // @[Mux.scala 46:19:@12286.4]
  wire [7:0] _T_16475; // @[Mux.scala 46:16:@12287.4]
  wire  _T_16476; // @[Mux.scala 46:19:@12288.4]
  wire [7:0] _T_16477; // @[Mux.scala 46:16:@12289.4]
  wire  _T_16478; // @[Mux.scala 46:19:@12290.4]
  wire [7:0] _T_16479; // @[Mux.scala 46:16:@12291.4]
  wire  _T_16480; // @[Mux.scala 46:19:@12292.4]
  wire [7:0] _T_16481; // @[Mux.scala 46:16:@12293.4]
  wire  _T_16482; // @[Mux.scala 46:19:@12294.4]
  wire [7:0] _T_16483; // @[Mux.scala 46:16:@12295.4]
  wire  _T_16484; // @[Mux.scala 46:19:@12296.4]
  wire [7:0] _T_16485; // @[Mux.scala 46:16:@12297.4]
  wire  _T_16486; // @[Mux.scala 46:19:@12298.4]
  wire [7:0] _T_16487; // @[Mux.scala 46:16:@12299.4]
  wire  _T_16488; // @[Mux.scala 46:19:@12300.4]
  wire [7:0] _T_16489; // @[Mux.scala 46:16:@12301.4]
  wire  _T_16490; // @[Mux.scala 46:19:@12302.4]
  wire [7:0] _T_16491; // @[Mux.scala 46:16:@12303.4]
  wire  _T_16492; // @[Mux.scala 46:19:@12304.4]
  wire [7:0] _T_16493; // @[Mux.scala 46:16:@12305.4]
  wire  _T_16494; // @[Mux.scala 46:19:@12306.4]
  wire [7:0] _T_16495; // @[Mux.scala 46:16:@12307.4]
  wire  _T_16496; // @[Mux.scala 46:19:@12308.4]
  wire [7:0] _T_16497; // @[Mux.scala 46:16:@12309.4]
  wire  _T_16498; // @[Mux.scala 46:19:@12310.4]
  wire [7:0] _T_16499; // @[Mux.scala 46:16:@12311.4]
  wire  _T_16500; // @[Mux.scala 46:19:@12312.4]
  wire [7:0] _T_16501; // @[Mux.scala 46:16:@12313.4]
  wire  _T_16502; // @[Mux.scala 46:19:@12314.4]
  wire [7:0] _T_16503; // @[Mux.scala 46:16:@12315.4]
  wire  _T_16504; // @[Mux.scala 46:19:@12316.4]
  wire [7:0] _T_16505; // @[Mux.scala 46:16:@12317.4]
  wire  _T_16506; // @[Mux.scala 46:19:@12318.4]
  wire [7:0] _T_16507; // @[Mux.scala 46:16:@12319.4]
  wire  _T_16508; // @[Mux.scala 46:19:@12320.4]
  wire [7:0] _T_16509; // @[Mux.scala 46:16:@12321.4]
  wire  _T_16510; // @[Mux.scala 46:19:@12322.4]
  wire [7:0] _T_16511; // @[Mux.scala 46:16:@12323.4]
  wire  _T_16512; // @[Mux.scala 46:19:@12324.4]
  wire [7:0] _T_16513; // @[Mux.scala 46:16:@12325.4]
  wire  _T_16514; // @[Mux.scala 46:19:@12326.4]
  wire [7:0] _T_16515; // @[Mux.scala 46:16:@12327.4]
  wire  _T_16516; // @[Mux.scala 46:19:@12328.4]
  wire [7:0] _T_16517; // @[Mux.scala 46:16:@12329.4]
  wire  _T_16518; // @[Mux.scala 46:19:@12330.4]
  wire [7:0] _T_16519; // @[Mux.scala 46:16:@12331.4]
  wire  _T_16520; // @[Mux.scala 46:19:@12332.4]
  wire [7:0] _T_16521; // @[Mux.scala 46:16:@12333.4]
  wire  _T_16522; // @[Mux.scala 46:19:@12334.4]
  wire [7:0] _T_16523; // @[Mux.scala 46:16:@12335.4]
  wire  _T_16524; // @[Mux.scala 46:19:@12336.4]
  wire [7:0] _T_16525; // @[Mux.scala 46:16:@12337.4]
  wire  _T_16526; // @[Mux.scala 46:19:@12338.4]
  wire [7:0] _T_16527; // @[Mux.scala 46:16:@12339.4]
  wire  _T_16528; // @[Mux.scala 46:19:@12340.4]
  wire [7:0] _T_16529; // @[Mux.scala 46:16:@12341.4]
  wire  _T_16530; // @[Mux.scala 46:19:@12342.4]
  wire [7:0] _T_16531; // @[Mux.scala 46:16:@12343.4]
  wire  _T_16591; // @[Mux.scala 46:19:@12345.4]
  wire [7:0] _T_16592; // @[Mux.scala 46:16:@12346.4]
  wire  _T_16593; // @[Mux.scala 46:19:@12347.4]
  wire [7:0] _T_16594; // @[Mux.scala 46:16:@12348.4]
  wire  _T_16595; // @[Mux.scala 46:19:@12349.4]
  wire [7:0] _T_16596; // @[Mux.scala 46:16:@12350.4]
  wire  _T_16597; // @[Mux.scala 46:19:@12351.4]
  wire [7:0] _T_16598; // @[Mux.scala 46:16:@12352.4]
  wire  _T_16599; // @[Mux.scala 46:19:@12353.4]
  wire [7:0] _T_16600; // @[Mux.scala 46:16:@12354.4]
  wire  _T_16601; // @[Mux.scala 46:19:@12355.4]
  wire [7:0] _T_16602; // @[Mux.scala 46:16:@12356.4]
  wire  _T_16603; // @[Mux.scala 46:19:@12357.4]
  wire [7:0] _T_16604; // @[Mux.scala 46:16:@12358.4]
  wire  _T_16605; // @[Mux.scala 46:19:@12359.4]
  wire [7:0] _T_16606; // @[Mux.scala 46:16:@12360.4]
  wire  _T_16607; // @[Mux.scala 46:19:@12361.4]
  wire [7:0] _T_16608; // @[Mux.scala 46:16:@12362.4]
  wire  _T_16609; // @[Mux.scala 46:19:@12363.4]
  wire [7:0] _T_16610; // @[Mux.scala 46:16:@12364.4]
  wire  _T_16611; // @[Mux.scala 46:19:@12365.4]
  wire [7:0] _T_16612; // @[Mux.scala 46:16:@12366.4]
  wire  _T_16613; // @[Mux.scala 46:19:@12367.4]
  wire [7:0] _T_16614; // @[Mux.scala 46:16:@12368.4]
  wire  _T_16615; // @[Mux.scala 46:19:@12369.4]
  wire [7:0] _T_16616; // @[Mux.scala 46:16:@12370.4]
  wire  _T_16617; // @[Mux.scala 46:19:@12371.4]
  wire [7:0] _T_16618; // @[Mux.scala 46:16:@12372.4]
  wire  _T_16619; // @[Mux.scala 46:19:@12373.4]
  wire [7:0] _T_16620; // @[Mux.scala 46:16:@12374.4]
  wire  _T_16621; // @[Mux.scala 46:19:@12375.4]
  wire [7:0] _T_16622; // @[Mux.scala 46:16:@12376.4]
  wire  _T_16623; // @[Mux.scala 46:19:@12377.4]
  wire [7:0] _T_16624; // @[Mux.scala 46:16:@12378.4]
  wire  _T_16625; // @[Mux.scala 46:19:@12379.4]
  wire [7:0] _T_16626; // @[Mux.scala 46:16:@12380.4]
  wire  _T_16627; // @[Mux.scala 46:19:@12381.4]
  wire [7:0] _T_16628; // @[Mux.scala 46:16:@12382.4]
  wire  _T_16629; // @[Mux.scala 46:19:@12383.4]
  wire [7:0] _T_16630; // @[Mux.scala 46:16:@12384.4]
  wire  _T_16631; // @[Mux.scala 46:19:@12385.4]
  wire [7:0] _T_16632; // @[Mux.scala 46:16:@12386.4]
  wire  _T_16633; // @[Mux.scala 46:19:@12387.4]
  wire [7:0] _T_16634; // @[Mux.scala 46:16:@12388.4]
  wire  _T_16635; // @[Mux.scala 46:19:@12389.4]
  wire [7:0] _T_16636; // @[Mux.scala 46:16:@12390.4]
  wire  _T_16637; // @[Mux.scala 46:19:@12391.4]
  wire [7:0] _T_16638; // @[Mux.scala 46:16:@12392.4]
  wire  _T_16639; // @[Mux.scala 46:19:@12393.4]
  wire [7:0] _T_16640; // @[Mux.scala 46:16:@12394.4]
  wire  _T_16641; // @[Mux.scala 46:19:@12395.4]
  wire [7:0] _T_16642; // @[Mux.scala 46:16:@12396.4]
  wire  _T_16643; // @[Mux.scala 46:19:@12397.4]
  wire [7:0] _T_16644; // @[Mux.scala 46:16:@12398.4]
  wire  _T_16645; // @[Mux.scala 46:19:@12399.4]
  wire [7:0] _T_16646; // @[Mux.scala 46:16:@12400.4]
  wire  _T_16647; // @[Mux.scala 46:19:@12401.4]
  wire [7:0] _T_16648; // @[Mux.scala 46:16:@12402.4]
  wire  _T_16649; // @[Mux.scala 46:19:@12403.4]
  wire [7:0] _T_16650; // @[Mux.scala 46:16:@12404.4]
  wire  _T_16651; // @[Mux.scala 46:19:@12405.4]
  wire [7:0] _T_16652; // @[Mux.scala 46:16:@12406.4]
  wire  _T_16653; // @[Mux.scala 46:19:@12407.4]
  wire [7:0] _T_16654; // @[Mux.scala 46:16:@12408.4]
  wire  _T_16655; // @[Mux.scala 46:19:@12409.4]
  wire [7:0] _T_16656; // @[Mux.scala 46:16:@12410.4]
  wire  _T_16657; // @[Mux.scala 46:19:@12411.4]
  wire [7:0] _T_16658; // @[Mux.scala 46:16:@12412.4]
  wire  _T_16659; // @[Mux.scala 46:19:@12413.4]
  wire [7:0] _T_16660; // @[Mux.scala 46:16:@12414.4]
  wire  _T_16661; // @[Mux.scala 46:19:@12415.4]
  wire [7:0] _T_16662; // @[Mux.scala 46:16:@12416.4]
  wire  _T_16663; // @[Mux.scala 46:19:@12417.4]
  wire [7:0] _T_16664; // @[Mux.scala 46:16:@12418.4]
  wire  _T_16665; // @[Mux.scala 46:19:@12419.4]
  wire [7:0] _T_16666; // @[Mux.scala 46:16:@12420.4]
  wire  _T_16667; // @[Mux.scala 46:19:@12421.4]
  wire [7:0] _T_16668; // @[Mux.scala 46:16:@12422.4]
  wire  _T_16669; // @[Mux.scala 46:19:@12423.4]
  wire [7:0] _T_16670; // @[Mux.scala 46:16:@12424.4]
  wire  _T_16671; // @[Mux.scala 46:19:@12425.4]
  wire [7:0] _T_16672; // @[Mux.scala 46:16:@12426.4]
  wire  _T_16673; // @[Mux.scala 46:19:@12427.4]
  wire [7:0] _T_16674; // @[Mux.scala 46:16:@12428.4]
  wire  _T_16675; // @[Mux.scala 46:19:@12429.4]
  wire [7:0] _T_16676; // @[Mux.scala 46:16:@12430.4]
  wire  _T_16677; // @[Mux.scala 46:19:@12431.4]
  wire [7:0] _T_16678; // @[Mux.scala 46:16:@12432.4]
  wire  _T_16679; // @[Mux.scala 46:19:@12433.4]
  wire [7:0] _T_16680; // @[Mux.scala 46:16:@12434.4]
  wire  _T_16681; // @[Mux.scala 46:19:@12435.4]
  wire [7:0] _T_16682; // @[Mux.scala 46:16:@12436.4]
  wire  _T_16683; // @[Mux.scala 46:19:@12437.4]
  wire [7:0] _T_16684; // @[Mux.scala 46:16:@12438.4]
  wire  _T_16685; // @[Mux.scala 46:19:@12439.4]
  wire [7:0] _T_16686; // @[Mux.scala 46:16:@12440.4]
  wire  _T_16687; // @[Mux.scala 46:19:@12441.4]
  wire [7:0] _T_16688; // @[Mux.scala 46:16:@12442.4]
  wire  _T_16689; // @[Mux.scala 46:19:@12443.4]
  wire [7:0] _T_16690; // @[Mux.scala 46:16:@12444.4]
  wire  _T_16691; // @[Mux.scala 46:19:@12445.4]
  wire [7:0] _T_16692; // @[Mux.scala 46:16:@12446.4]
  wire  _T_16693; // @[Mux.scala 46:19:@12447.4]
  wire [7:0] _T_16694; // @[Mux.scala 46:16:@12448.4]
  wire  _T_16695; // @[Mux.scala 46:19:@12449.4]
  wire [7:0] _T_16696; // @[Mux.scala 46:16:@12450.4]
  wire  _T_16697; // @[Mux.scala 46:19:@12451.4]
  wire [7:0] _T_16698; // @[Mux.scala 46:16:@12452.4]
  wire  _T_16699; // @[Mux.scala 46:19:@12453.4]
  wire [7:0] _T_16700; // @[Mux.scala 46:16:@12454.4]
  wire  _T_16701; // @[Mux.scala 46:19:@12455.4]
  wire [7:0] _T_16702; // @[Mux.scala 46:16:@12456.4]
  wire  _T_16703; // @[Mux.scala 46:19:@12457.4]
  wire [7:0] _T_16704; // @[Mux.scala 46:16:@12458.4]
  wire  _T_16705; // @[Mux.scala 46:19:@12459.4]
  wire [7:0] _T_16706; // @[Mux.scala 46:16:@12460.4]
  wire  _T_16767; // @[Mux.scala 46:19:@12462.4]
  wire [7:0] _T_16768; // @[Mux.scala 46:16:@12463.4]
  wire  _T_16769; // @[Mux.scala 46:19:@12464.4]
  wire [7:0] _T_16770; // @[Mux.scala 46:16:@12465.4]
  wire  _T_16771; // @[Mux.scala 46:19:@12466.4]
  wire [7:0] _T_16772; // @[Mux.scala 46:16:@12467.4]
  wire  _T_16773; // @[Mux.scala 46:19:@12468.4]
  wire [7:0] _T_16774; // @[Mux.scala 46:16:@12469.4]
  wire  _T_16775; // @[Mux.scala 46:19:@12470.4]
  wire [7:0] _T_16776; // @[Mux.scala 46:16:@12471.4]
  wire  _T_16777; // @[Mux.scala 46:19:@12472.4]
  wire [7:0] _T_16778; // @[Mux.scala 46:16:@12473.4]
  wire  _T_16779; // @[Mux.scala 46:19:@12474.4]
  wire [7:0] _T_16780; // @[Mux.scala 46:16:@12475.4]
  wire  _T_16781; // @[Mux.scala 46:19:@12476.4]
  wire [7:0] _T_16782; // @[Mux.scala 46:16:@12477.4]
  wire  _T_16783; // @[Mux.scala 46:19:@12478.4]
  wire [7:0] _T_16784; // @[Mux.scala 46:16:@12479.4]
  wire  _T_16785; // @[Mux.scala 46:19:@12480.4]
  wire [7:0] _T_16786; // @[Mux.scala 46:16:@12481.4]
  wire  _T_16787; // @[Mux.scala 46:19:@12482.4]
  wire [7:0] _T_16788; // @[Mux.scala 46:16:@12483.4]
  wire  _T_16789; // @[Mux.scala 46:19:@12484.4]
  wire [7:0] _T_16790; // @[Mux.scala 46:16:@12485.4]
  wire  _T_16791; // @[Mux.scala 46:19:@12486.4]
  wire [7:0] _T_16792; // @[Mux.scala 46:16:@12487.4]
  wire  _T_16793; // @[Mux.scala 46:19:@12488.4]
  wire [7:0] _T_16794; // @[Mux.scala 46:16:@12489.4]
  wire  _T_16795; // @[Mux.scala 46:19:@12490.4]
  wire [7:0] _T_16796; // @[Mux.scala 46:16:@12491.4]
  wire  _T_16797; // @[Mux.scala 46:19:@12492.4]
  wire [7:0] _T_16798; // @[Mux.scala 46:16:@12493.4]
  wire  _T_16799; // @[Mux.scala 46:19:@12494.4]
  wire [7:0] _T_16800; // @[Mux.scala 46:16:@12495.4]
  wire  _T_16801; // @[Mux.scala 46:19:@12496.4]
  wire [7:0] _T_16802; // @[Mux.scala 46:16:@12497.4]
  wire  _T_16803; // @[Mux.scala 46:19:@12498.4]
  wire [7:0] _T_16804; // @[Mux.scala 46:16:@12499.4]
  wire  _T_16805; // @[Mux.scala 46:19:@12500.4]
  wire [7:0] _T_16806; // @[Mux.scala 46:16:@12501.4]
  wire  _T_16807; // @[Mux.scala 46:19:@12502.4]
  wire [7:0] _T_16808; // @[Mux.scala 46:16:@12503.4]
  wire  _T_16809; // @[Mux.scala 46:19:@12504.4]
  wire [7:0] _T_16810; // @[Mux.scala 46:16:@12505.4]
  wire  _T_16811; // @[Mux.scala 46:19:@12506.4]
  wire [7:0] _T_16812; // @[Mux.scala 46:16:@12507.4]
  wire  _T_16813; // @[Mux.scala 46:19:@12508.4]
  wire [7:0] _T_16814; // @[Mux.scala 46:16:@12509.4]
  wire  _T_16815; // @[Mux.scala 46:19:@12510.4]
  wire [7:0] _T_16816; // @[Mux.scala 46:16:@12511.4]
  wire  _T_16817; // @[Mux.scala 46:19:@12512.4]
  wire [7:0] _T_16818; // @[Mux.scala 46:16:@12513.4]
  wire  _T_16819; // @[Mux.scala 46:19:@12514.4]
  wire [7:0] _T_16820; // @[Mux.scala 46:16:@12515.4]
  wire  _T_16821; // @[Mux.scala 46:19:@12516.4]
  wire [7:0] _T_16822; // @[Mux.scala 46:16:@12517.4]
  wire  _T_16823; // @[Mux.scala 46:19:@12518.4]
  wire [7:0] _T_16824; // @[Mux.scala 46:16:@12519.4]
  wire  _T_16825; // @[Mux.scala 46:19:@12520.4]
  wire [7:0] _T_16826; // @[Mux.scala 46:16:@12521.4]
  wire  _T_16827; // @[Mux.scala 46:19:@12522.4]
  wire [7:0] _T_16828; // @[Mux.scala 46:16:@12523.4]
  wire  _T_16829; // @[Mux.scala 46:19:@12524.4]
  wire [7:0] _T_16830; // @[Mux.scala 46:16:@12525.4]
  wire  _T_16831; // @[Mux.scala 46:19:@12526.4]
  wire [7:0] _T_16832; // @[Mux.scala 46:16:@12527.4]
  wire  _T_16833; // @[Mux.scala 46:19:@12528.4]
  wire [7:0] _T_16834; // @[Mux.scala 46:16:@12529.4]
  wire  _T_16835; // @[Mux.scala 46:19:@12530.4]
  wire [7:0] _T_16836; // @[Mux.scala 46:16:@12531.4]
  wire  _T_16837; // @[Mux.scala 46:19:@12532.4]
  wire [7:0] _T_16838; // @[Mux.scala 46:16:@12533.4]
  wire  _T_16839; // @[Mux.scala 46:19:@12534.4]
  wire [7:0] _T_16840; // @[Mux.scala 46:16:@12535.4]
  wire  _T_16841; // @[Mux.scala 46:19:@12536.4]
  wire [7:0] _T_16842; // @[Mux.scala 46:16:@12537.4]
  wire  _T_16843; // @[Mux.scala 46:19:@12538.4]
  wire [7:0] _T_16844; // @[Mux.scala 46:16:@12539.4]
  wire  _T_16845; // @[Mux.scala 46:19:@12540.4]
  wire [7:0] _T_16846; // @[Mux.scala 46:16:@12541.4]
  wire  _T_16847; // @[Mux.scala 46:19:@12542.4]
  wire [7:0] _T_16848; // @[Mux.scala 46:16:@12543.4]
  wire  _T_16849; // @[Mux.scala 46:19:@12544.4]
  wire [7:0] _T_16850; // @[Mux.scala 46:16:@12545.4]
  wire  _T_16851; // @[Mux.scala 46:19:@12546.4]
  wire [7:0] _T_16852; // @[Mux.scala 46:16:@12547.4]
  wire  _T_16853; // @[Mux.scala 46:19:@12548.4]
  wire [7:0] _T_16854; // @[Mux.scala 46:16:@12549.4]
  wire  _T_16855; // @[Mux.scala 46:19:@12550.4]
  wire [7:0] _T_16856; // @[Mux.scala 46:16:@12551.4]
  wire  _T_16857; // @[Mux.scala 46:19:@12552.4]
  wire [7:0] _T_16858; // @[Mux.scala 46:16:@12553.4]
  wire  _T_16859; // @[Mux.scala 46:19:@12554.4]
  wire [7:0] _T_16860; // @[Mux.scala 46:16:@12555.4]
  wire  _T_16861; // @[Mux.scala 46:19:@12556.4]
  wire [7:0] _T_16862; // @[Mux.scala 46:16:@12557.4]
  wire  _T_16863; // @[Mux.scala 46:19:@12558.4]
  wire [7:0] _T_16864; // @[Mux.scala 46:16:@12559.4]
  wire  _T_16865; // @[Mux.scala 46:19:@12560.4]
  wire [7:0] _T_16866; // @[Mux.scala 46:16:@12561.4]
  wire  _T_16867; // @[Mux.scala 46:19:@12562.4]
  wire [7:0] _T_16868; // @[Mux.scala 46:16:@12563.4]
  wire  _T_16869; // @[Mux.scala 46:19:@12564.4]
  wire [7:0] _T_16870; // @[Mux.scala 46:16:@12565.4]
  wire  _T_16871; // @[Mux.scala 46:19:@12566.4]
  wire [7:0] _T_16872; // @[Mux.scala 46:16:@12567.4]
  wire  _T_16873; // @[Mux.scala 46:19:@12568.4]
  wire [7:0] _T_16874; // @[Mux.scala 46:16:@12569.4]
  wire  _T_16875; // @[Mux.scala 46:19:@12570.4]
  wire [7:0] _T_16876; // @[Mux.scala 46:16:@12571.4]
  wire  _T_16877; // @[Mux.scala 46:19:@12572.4]
  wire [7:0] _T_16878; // @[Mux.scala 46:16:@12573.4]
  wire  _T_16879; // @[Mux.scala 46:19:@12574.4]
  wire [7:0] _T_16880; // @[Mux.scala 46:16:@12575.4]
  wire  _T_16881; // @[Mux.scala 46:19:@12576.4]
  wire [7:0] _T_16882; // @[Mux.scala 46:16:@12577.4]
  wire  _T_16883; // @[Mux.scala 46:19:@12578.4]
  wire [7:0] _T_16884; // @[Mux.scala 46:16:@12579.4]
  wire  _T_16946; // @[Mux.scala 46:19:@12581.4]
  wire [7:0] _T_16947; // @[Mux.scala 46:16:@12582.4]
  wire  _T_16948; // @[Mux.scala 46:19:@12583.4]
  wire [7:0] _T_16949; // @[Mux.scala 46:16:@12584.4]
  wire  _T_16950; // @[Mux.scala 46:19:@12585.4]
  wire [7:0] _T_16951; // @[Mux.scala 46:16:@12586.4]
  wire  _T_16952; // @[Mux.scala 46:19:@12587.4]
  wire [7:0] _T_16953; // @[Mux.scala 46:16:@12588.4]
  wire  _T_16954; // @[Mux.scala 46:19:@12589.4]
  wire [7:0] _T_16955; // @[Mux.scala 46:16:@12590.4]
  wire  _T_16956; // @[Mux.scala 46:19:@12591.4]
  wire [7:0] _T_16957; // @[Mux.scala 46:16:@12592.4]
  wire  _T_16958; // @[Mux.scala 46:19:@12593.4]
  wire [7:0] _T_16959; // @[Mux.scala 46:16:@12594.4]
  wire  _T_16960; // @[Mux.scala 46:19:@12595.4]
  wire [7:0] _T_16961; // @[Mux.scala 46:16:@12596.4]
  wire  _T_16962; // @[Mux.scala 46:19:@12597.4]
  wire [7:0] _T_16963; // @[Mux.scala 46:16:@12598.4]
  wire  _T_16964; // @[Mux.scala 46:19:@12599.4]
  wire [7:0] _T_16965; // @[Mux.scala 46:16:@12600.4]
  wire  _T_16966; // @[Mux.scala 46:19:@12601.4]
  wire [7:0] _T_16967; // @[Mux.scala 46:16:@12602.4]
  wire  _T_16968; // @[Mux.scala 46:19:@12603.4]
  wire [7:0] _T_16969; // @[Mux.scala 46:16:@12604.4]
  wire  _T_16970; // @[Mux.scala 46:19:@12605.4]
  wire [7:0] _T_16971; // @[Mux.scala 46:16:@12606.4]
  wire  _T_16972; // @[Mux.scala 46:19:@12607.4]
  wire [7:0] _T_16973; // @[Mux.scala 46:16:@12608.4]
  wire  _T_16974; // @[Mux.scala 46:19:@12609.4]
  wire [7:0] _T_16975; // @[Mux.scala 46:16:@12610.4]
  wire  _T_16976; // @[Mux.scala 46:19:@12611.4]
  wire [7:0] _T_16977; // @[Mux.scala 46:16:@12612.4]
  wire  _T_16978; // @[Mux.scala 46:19:@12613.4]
  wire [7:0] _T_16979; // @[Mux.scala 46:16:@12614.4]
  wire  _T_16980; // @[Mux.scala 46:19:@12615.4]
  wire [7:0] _T_16981; // @[Mux.scala 46:16:@12616.4]
  wire  _T_16982; // @[Mux.scala 46:19:@12617.4]
  wire [7:0] _T_16983; // @[Mux.scala 46:16:@12618.4]
  wire  _T_16984; // @[Mux.scala 46:19:@12619.4]
  wire [7:0] _T_16985; // @[Mux.scala 46:16:@12620.4]
  wire  _T_16986; // @[Mux.scala 46:19:@12621.4]
  wire [7:0] _T_16987; // @[Mux.scala 46:16:@12622.4]
  wire  _T_16988; // @[Mux.scala 46:19:@12623.4]
  wire [7:0] _T_16989; // @[Mux.scala 46:16:@12624.4]
  wire  _T_16990; // @[Mux.scala 46:19:@12625.4]
  wire [7:0] _T_16991; // @[Mux.scala 46:16:@12626.4]
  wire  _T_16992; // @[Mux.scala 46:19:@12627.4]
  wire [7:0] _T_16993; // @[Mux.scala 46:16:@12628.4]
  wire  _T_16994; // @[Mux.scala 46:19:@12629.4]
  wire [7:0] _T_16995; // @[Mux.scala 46:16:@12630.4]
  wire  _T_16996; // @[Mux.scala 46:19:@12631.4]
  wire [7:0] _T_16997; // @[Mux.scala 46:16:@12632.4]
  wire  _T_16998; // @[Mux.scala 46:19:@12633.4]
  wire [7:0] _T_16999; // @[Mux.scala 46:16:@12634.4]
  wire  _T_17000; // @[Mux.scala 46:19:@12635.4]
  wire [7:0] _T_17001; // @[Mux.scala 46:16:@12636.4]
  wire  _T_17002; // @[Mux.scala 46:19:@12637.4]
  wire [7:0] _T_17003; // @[Mux.scala 46:16:@12638.4]
  wire  _T_17004; // @[Mux.scala 46:19:@12639.4]
  wire [7:0] _T_17005; // @[Mux.scala 46:16:@12640.4]
  wire  _T_17006; // @[Mux.scala 46:19:@12641.4]
  wire [7:0] _T_17007; // @[Mux.scala 46:16:@12642.4]
  wire  _T_17008; // @[Mux.scala 46:19:@12643.4]
  wire [7:0] _T_17009; // @[Mux.scala 46:16:@12644.4]
  wire  _T_17010; // @[Mux.scala 46:19:@12645.4]
  wire [7:0] _T_17011; // @[Mux.scala 46:16:@12646.4]
  wire  _T_17012; // @[Mux.scala 46:19:@12647.4]
  wire [7:0] _T_17013; // @[Mux.scala 46:16:@12648.4]
  wire  _T_17014; // @[Mux.scala 46:19:@12649.4]
  wire [7:0] _T_17015; // @[Mux.scala 46:16:@12650.4]
  wire  _T_17016; // @[Mux.scala 46:19:@12651.4]
  wire [7:0] _T_17017; // @[Mux.scala 46:16:@12652.4]
  wire  _T_17018; // @[Mux.scala 46:19:@12653.4]
  wire [7:0] _T_17019; // @[Mux.scala 46:16:@12654.4]
  wire  _T_17020; // @[Mux.scala 46:19:@12655.4]
  wire [7:0] _T_17021; // @[Mux.scala 46:16:@12656.4]
  wire  _T_17022; // @[Mux.scala 46:19:@12657.4]
  wire [7:0] _T_17023; // @[Mux.scala 46:16:@12658.4]
  wire  _T_17024; // @[Mux.scala 46:19:@12659.4]
  wire [7:0] _T_17025; // @[Mux.scala 46:16:@12660.4]
  wire  _T_17026; // @[Mux.scala 46:19:@12661.4]
  wire [7:0] _T_17027; // @[Mux.scala 46:16:@12662.4]
  wire  _T_17028; // @[Mux.scala 46:19:@12663.4]
  wire [7:0] _T_17029; // @[Mux.scala 46:16:@12664.4]
  wire  _T_17030; // @[Mux.scala 46:19:@12665.4]
  wire [7:0] _T_17031; // @[Mux.scala 46:16:@12666.4]
  wire  _T_17032; // @[Mux.scala 46:19:@12667.4]
  wire [7:0] _T_17033; // @[Mux.scala 46:16:@12668.4]
  wire  _T_17034; // @[Mux.scala 46:19:@12669.4]
  wire [7:0] _T_17035; // @[Mux.scala 46:16:@12670.4]
  wire  _T_17036; // @[Mux.scala 46:19:@12671.4]
  wire [7:0] _T_17037; // @[Mux.scala 46:16:@12672.4]
  wire  _T_17038; // @[Mux.scala 46:19:@12673.4]
  wire [7:0] _T_17039; // @[Mux.scala 46:16:@12674.4]
  wire  _T_17040; // @[Mux.scala 46:19:@12675.4]
  wire [7:0] _T_17041; // @[Mux.scala 46:16:@12676.4]
  wire  _T_17042; // @[Mux.scala 46:19:@12677.4]
  wire [7:0] _T_17043; // @[Mux.scala 46:16:@12678.4]
  wire  _T_17044; // @[Mux.scala 46:19:@12679.4]
  wire [7:0] _T_17045; // @[Mux.scala 46:16:@12680.4]
  wire  _T_17046; // @[Mux.scala 46:19:@12681.4]
  wire [7:0] _T_17047; // @[Mux.scala 46:16:@12682.4]
  wire  _T_17048; // @[Mux.scala 46:19:@12683.4]
  wire [7:0] _T_17049; // @[Mux.scala 46:16:@12684.4]
  wire  _T_17050; // @[Mux.scala 46:19:@12685.4]
  wire [7:0] _T_17051; // @[Mux.scala 46:16:@12686.4]
  wire  _T_17052; // @[Mux.scala 46:19:@12687.4]
  wire [7:0] _T_17053; // @[Mux.scala 46:16:@12688.4]
  wire  _T_17054; // @[Mux.scala 46:19:@12689.4]
  wire [7:0] _T_17055; // @[Mux.scala 46:16:@12690.4]
  wire  _T_17056; // @[Mux.scala 46:19:@12691.4]
  wire [7:0] _T_17057; // @[Mux.scala 46:16:@12692.4]
  wire  _T_17058; // @[Mux.scala 46:19:@12693.4]
  wire [7:0] _T_17059; // @[Mux.scala 46:16:@12694.4]
  wire  _T_17060; // @[Mux.scala 46:19:@12695.4]
  wire [7:0] _T_17061; // @[Mux.scala 46:16:@12696.4]
  wire  _T_17062; // @[Mux.scala 46:19:@12697.4]
  wire [7:0] _T_17063; // @[Mux.scala 46:16:@12698.4]
  wire  _T_17064; // @[Mux.scala 46:19:@12699.4]
  wire [7:0] _T_17065; // @[Mux.scala 46:16:@12700.4]
  wire  _T_17128; // @[Mux.scala 46:19:@12702.4]
  wire [7:0] _T_17129; // @[Mux.scala 46:16:@12703.4]
  wire  _T_17130; // @[Mux.scala 46:19:@12704.4]
  wire [7:0] _T_17131; // @[Mux.scala 46:16:@12705.4]
  wire  _T_17132; // @[Mux.scala 46:19:@12706.4]
  wire [7:0] _T_17133; // @[Mux.scala 46:16:@12707.4]
  wire  _T_17134; // @[Mux.scala 46:19:@12708.4]
  wire [7:0] _T_17135; // @[Mux.scala 46:16:@12709.4]
  wire  _T_17136; // @[Mux.scala 46:19:@12710.4]
  wire [7:0] _T_17137; // @[Mux.scala 46:16:@12711.4]
  wire  _T_17138; // @[Mux.scala 46:19:@12712.4]
  wire [7:0] _T_17139; // @[Mux.scala 46:16:@12713.4]
  wire  _T_17140; // @[Mux.scala 46:19:@12714.4]
  wire [7:0] _T_17141; // @[Mux.scala 46:16:@12715.4]
  wire  _T_17142; // @[Mux.scala 46:19:@12716.4]
  wire [7:0] _T_17143; // @[Mux.scala 46:16:@12717.4]
  wire  _T_17144; // @[Mux.scala 46:19:@12718.4]
  wire [7:0] _T_17145; // @[Mux.scala 46:16:@12719.4]
  wire  _T_17146; // @[Mux.scala 46:19:@12720.4]
  wire [7:0] _T_17147; // @[Mux.scala 46:16:@12721.4]
  wire  _T_17148; // @[Mux.scala 46:19:@12722.4]
  wire [7:0] _T_17149; // @[Mux.scala 46:16:@12723.4]
  wire  _T_17150; // @[Mux.scala 46:19:@12724.4]
  wire [7:0] _T_17151; // @[Mux.scala 46:16:@12725.4]
  wire  _T_17152; // @[Mux.scala 46:19:@12726.4]
  wire [7:0] _T_17153; // @[Mux.scala 46:16:@12727.4]
  wire  _T_17154; // @[Mux.scala 46:19:@12728.4]
  wire [7:0] _T_17155; // @[Mux.scala 46:16:@12729.4]
  wire  _T_17156; // @[Mux.scala 46:19:@12730.4]
  wire [7:0] _T_17157; // @[Mux.scala 46:16:@12731.4]
  wire  _T_17158; // @[Mux.scala 46:19:@12732.4]
  wire [7:0] _T_17159; // @[Mux.scala 46:16:@12733.4]
  wire  _T_17160; // @[Mux.scala 46:19:@12734.4]
  wire [7:0] _T_17161; // @[Mux.scala 46:16:@12735.4]
  wire  _T_17162; // @[Mux.scala 46:19:@12736.4]
  wire [7:0] _T_17163; // @[Mux.scala 46:16:@12737.4]
  wire  _T_17164; // @[Mux.scala 46:19:@12738.4]
  wire [7:0] _T_17165; // @[Mux.scala 46:16:@12739.4]
  wire  _T_17166; // @[Mux.scala 46:19:@12740.4]
  wire [7:0] _T_17167; // @[Mux.scala 46:16:@12741.4]
  wire  _T_17168; // @[Mux.scala 46:19:@12742.4]
  wire [7:0] _T_17169; // @[Mux.scala 46:16:@12743.4]
  wire  _T_17170; // @[Mux.scala 46:19:@12744.4]
  wire [7:0] _T_17171; // @[Mux.scala 46:16:@12745.4]
  wire  _T_17172; // @[Mux.scala 46:19:@12746.4]
  wire [7:0] _T_17173; // @[Mux.scala 46:16:@12747.4]
  wire  _T_17174; // @[Mux.scala 46:19:@12748.4]
  wire [7:0] _T_17175; // @[Mux.scala 46:16:@12749.4]
  wire  _T_17176; // @[Mux.scala 46:19:@12750.4]
  wire [7:0] _T_17177; // @[Mux.scala 46:16:@12751.4]
  wire  _T_17178; // @[Mux.scala 46:19:@12752.4]
  wire [7:0] _T_17179; // @[Mux.scala 46:16:@12753.4]
  wire  _T_17180; // @[Mux.scala 46:19:@12754.4]
  wire [7:0] _T_17181; // @[Mux.scala 46:16:@12755.4]
  wire  _T_17182; // @[Mux.scala 46:19:@12756.4]
  wire [7:0] _T_17183; // @[Mux.scala 46:16:@12757.4]
  wire  _T_17184; // @[Mux.scala 46:19:@12758.4]
  wire [7:0] _T_17185; // @[Mux.scala 46:16:@12759.4]
  wire  _T_17186; // @[Mux.scala 46:19:@12760.4]
  wire [7:0] _T_17187; // @[Mux.scala 46:16:@12761.4]
  wire  _T_17188; // @[Mux.scala 46:19:@12762.4]
  wire [7:0] _T_17189; // @[Mux.scala 46:16:@12763.4]
  wire  _T_17190; // @[Mux.scala 46:19:@12764.4]
  wire [7:0] _T_17191; // @[Mux.scala 46:16:@12765.4]
  wire  _T_17192; // @[Mux.scala 46:19:@12766.4]
  wire [7:0] _T_17193; // @[Mux.scala 46:16:@12767.4]
  wire  _T_17194; // @[Mux.scala 46:19:@12768.4]
  wire [7:0] _T_17195; // @[Mux.scala 46:16:@12769.4]
  wire  _T_17196; // @[Mux.scala 46:19:@12770.4]
  wire [7:0] _T_17197; // @[Mux.scala 46:16:@12771.4]
  wire  _T_17198; // @[Mux.scala 46:19:@12772.4]
  wire [7:0] _T_17199; // @[Mux.scala 46:16:@12773.4]
  wire  _T_17200; // @[Mux.scala 46:19:@12774.4]
  wire [7:0] _T_17201; // @[Mux.scala 46:16:@12775.4]
  wire  _T_17202; // @[Mux.scala 46:19:@12776.4]
  wire [7:0] _T_17203; // @[Mux.scala 46:16:@12777.4]
  wire  _T_17204; // @[Mux.scala 46:19:@12778.4]
  wire [7:0] _T_17205; // @[Mux.scala 46:16:@12779.4]
  wire  _T_17206; // @[Mux.scala 46:19:@12780.4]
  wire [7:0] _T_17207; // @[Mux.scala 46:16:@12781.4]
  wire  _T_17208; // @[Mux.scala 46:19:@12782.4]
  wire [7:0] _T_17209; // @[Mux.scala 46:16:@12783.4]
  wire  _T_17210; // @[Mux.scala 46:19:@12784.4]
  wire [7:0] _T_17211; // @[Mux.scala 46:16:@12785.4]
  wire  _T_17212; // @[Mux.scala 46:19:@12786.4]
  wire [7:0] _T_17213; // @[Mux.scala 46:16:@12787.4]
  wire  _T_17214; // @[Mux.scala 46:19:@12788.4]
  wire [7:0] _T_17215; // @[Mux.scala 46:16:@12789.4]
  wire  _T_17216; // @[Mux.scala 46:19:@12790.4]
  wire [7:0] _T_17217; // @[Mux.scala 46:16:@12791.4]
  wire  _T_17218; // @[Mux.scala 46:19:@12792.4]
  wire [7:0] _T_17219; // @[Mux.scala 46:16:@12793.4]
  wire  _T_17220; // @[Mux.scala 46:19:@12794.4]
  wire [7:0] _T_17221; // @[Mux.scala 46:16:@12795.4]
  wire  _T_17222; // @[Mux.scala 46:19:@12796.4]
  wire [7:0] _T_17223; // @[Mux.scala 46:16:@12797.4]
  wire  _T_17224; // @[Mux.scala 46:19:@12798.4]
  wire [7:0] _T_17225; // @[Mux.scala 46:16:@12799.4]
  wire  _T_17226; // @[Mux.scala 46:19:@12800.4]
  wire [7:0] _T_17227; // @[Mux.scala 46:16:@12801.4]
  wire  _T_17228; // @[Mux.scala 46:19:@12802.4]
  wire [7:0] _T_17229; // @[Mux.scala 46:16:@12803.4]
  wire  _T_17230; // @[Mux.scala 46:19:@12804.4]
  wire [7:0] _T_17231; // @[Mux.scala 46:16:@12805.4]
  wire  _T_17232; // @[Mux.scala 46:19:@12806.4]
  wire [7:0] _T_17233; // @[Mux.scala 46:16:@12807.4]
  wire  _T_17234; // @[Mux.scala 46:19:@12808.4]
  wire [7:0] _T_17235; // @[Mux.scala 46:16:@12809.4]
  wire  _T_17236; // @[Mux.scala 46:19:@12810.4]
  wire [7:0] _T_17237; // @[Mux.scala 46:16:@12811.4]
  wire  _T_17238; // @[Mux.scala 46:19:@12812.4]
  wire [7:0] _T_17239; // @[Mux.scala 46:16:@12813.4]
  wire  _T_17240; // @[Mux.scala 46:19:@12814.4]
  wire [7:0] _T_17241; // @[Mux.scala 46:16:@12815.4]
  wire  _T_17242; // @[Mux.scala 46:19:@12816.4]
  wire [7:0] _T_17243; // @[Mux.scala 46:16:@12817.4]
  wire  _T_17244; // @[Mux.scala 46:19:@12818.4]
  wire [7:0] _T_17245; // @[Mux.scala 46:16:@12819.4]
  wire  _T_17246; // @[Mux.scala 46:19:@12820.4]
  wire [7:0] _T_17247; // @[Mux.scala 46:16:@12821.4]
  wire  _T_17248; // @[Mux.scala 46:19:@12822.4]
  wire [7:0] _T_17249; // @[Mux.scala 46:16:@12823.4]
  wire  _T_17313; // @[Mux.scala 46:19:@12825.4]
  wire [7:0] _T_17314; // @[Mux.scala 46:16:@12826.4]
  wire  _T_17315; // @[Mux.scala 46:19:@12827.4]
  wire [7:0] _T_17316; // @[Mux.scala 46:16:@12828.4]
  wire  _T_17317; // @[Mux.scala 46:19:@12829.4]
  wire [7:0] _T_17318; // @[Mux.scala 46:16:@12830.4]
  wire  _T_17319; // @[Mux.scala 46:19:@12831.4]
  wire [7:0] _T_17320; // @[Mux.scala 46:16:@12832.4]
  wire  _T_17321; // @[Mux.scala 46:19:@12833.4]
  wire [7:0] _T_17322; // @[Mux.scala 46:16:@12834.4]
  wire  _T_17323; // @[Mux.scala 46:19:@12835.4]
  wire [7:0] _T_17324; // @[Mux.scala 46:16:@12836.4]
  wire  _T_17325; // @[Mux.scala 46:19:@12837.4]
  wire [7:0] _T_17326; // @[Mux.scala 46:16:@12838.4]
  wire  _T_17327; // @[Mux.scala 46:19:@12839.4]
  wire [7:0] _T_17328; // @[Mux.scala 46:16:@12840.4]
  wire  _T_17329; // @[Mux.scala 46:19:@12841.4]
  wire [7:0] _T_17330; // @[Mux.scala 46:16:@12842.4]
  wire  _T_17331; // @[Mux.scala 46:19:@12843.4]
  wire [7:0] _T_17332; // @[Mux.scala 46:16:@12844.4]
  wire  _T_17333; // @[Mux.scala 46:19:@12845.4]
  wire [7:0] _T_17334; // @[Mux.scala 46:16:@12846.4]
  wire  _T_17335; // @[Mux.scala 46:19:@12847.4]
  wire [7:0] _T_17336; // @[Mux.scala 46:16:@12848.4]
  wire  _T_17337; // @[Mux.scala 46:19:@12849.4]
  wire [7:0] _T_17338; // @[Mux.scala 46:16:@12850.4]
  wire  _T_17339; // @[Mux.scala 46:19:@12851.4]
  wire [7:0] _T_17340; // @[Mux.scala 46:16:@12852.4]
  wire  _T_17341; // @[Mux.scala 46:19:@12853.4]
  wire [7:0] _T_17342; // @[Mux.scala 46:16:@12854.4]
  wire  _T_17343; // @[Mux.scala 46:19:@12855.4]
  wire [7:0] _T_17344; // @[Mux.scala 46:16:@12856.4]
  wire  _T_17345; // @[Mux.scala 46:19:@12857.4]
  wire [7:0] _T_17346; // @[Mux.scala 46:16:@12858.4]
  wire  _T_17347; // @[Mux.scala 46:19:@12859.4]
  wire [7:0] _T_17348; // @[Mux.scala 46:16:@12860.4]
  wire  _T_17349; // @[Mux.scala 46:19:@12861.4]
  wire [7:0] _T_17350; // @[Mux.scala 46:16:@12862.4]
  wire  _T_17351; // @[Mux.scala 46:19:@12863.4]
  wire [7:0] _T_17352; // @[Mux.scala 46:16:@12864.4]
  wire  _T_17353; // @[Mux.scala 46:19:@12865.4]
  wire [7:0] _T_17354; // @[Mux.scala 46:16:@12866.4]
  wire  _T_17355; // @[Mux.scala 46:19:@12867.4]
  wire [7:0] _T_17356; // @[Mux.scala 46:16:@12868.4]
  wire  _T_17357; // @[Mux.scala 46:19:@12869.4]
  wire [7:0] _T_17358; // @[Mux.scala 46:16:@12870.4]
  wire  _T_17359; // @[Mux.scala 46:19:@12871.4]
  wire [7:0] _T_17360; // @[Mux.scala 46:16:@12872.4]
  wire  _T_17361; // @[Mux.scala 46:19:@12873.4]
  wire [7:0] _T_17362; // @[Mux.scala 46:16:@12874.4]
  wire  _T_17363; // @[Mux.scala 46:19:@12875.4]
  wire [7:0] _T_17364; // @[Mux.scala 46:16:@12876.4]
  wire  _T_17365; // @[Mux.scala 46:19:@12877.4]
  wire [7:0] _T_17366; // @[Mux.scala 46:16:@12878.4]
  wire  _T_17367; // @[Mux.scala 46:19:@12879.4]
  wire [7:0] _T_17368; // @[Mux.scala 46:16:@12880.4]
  wire  _T_17369; // @[Mux.scala 46:19:@12881.4]
  wire [7:0] _T_17370; // @[Mux.scala 46:16:@12882.4]
  wire  _T_17371; // @[Mux.scala 46:19:@12883.4]
  wire [7:0] _T_17372; // @[Mux.scala 46:16:@12884.4]
  wire  _T_17373; // @[Mux.scala 46:19:@12885.4]
  wire [7:0] _T_17374; // @[Mux.scala 46:16:@12886.4]
  wire  _T_17375; // @[Mux.scala 46:19:@12887.4]
  wire [7:0] _T_17376; // @[Mux.scala 46:16:@12888.4]
  wire  _T_17377; // @[Mux.scala 46:19:@12889.4]
  wire [7:0] _T_17378; // @[Mux.scala 46:16:@12890.4]
  wire  _T_17379; // @[Mux.scala 46:19:@12891.4]
  wire [7:0] _T_17380; // @[Mux.scala 46:16:@12892.4]
  wire  _T_17381; // @[Mux.scala 46:19:@12893.4]
  wire [7:0] _T_17382; // @[Mux.scala 46:16:@12894.4]
  wire  _T_17383; // @[Mux.scala 46:19:@12895.4]
  wire [7:0] _T_17384; // @[Mux.scala 46:16:@12896.4]
  wire  _T_17385; // @[Mux.scala 46:19:@12897.4]
  wire [7:0] _T_17386; // @[Mux.scala 46:16:@12898.4]
  wire  _T_17387; // @[Mux.scala 46:19:@12899.4]
  wire [7:0] _T_17388; // @[Mux.scala 46:16:@12900.4]
  wire  _T_17389; // @[Mux.scala 46:19:@12901.4]
  wire [7:0] _T_17390; // @[Mux.scala 46:16:@12902.4]
  wire  _T_17391; // @[Mux.scala 46:19:@12903.4]
  wire [7:0] _T_17392; // @[Mux.scala 46:16:@12904.4]
  wire  _T_17393; // @[Mux.scala 46:19:@12905.4]
  wire [7:0] _T_17394; // @[Mux.scala 46:16:@12906.4]
  wire  _T_17395; // @[Mux.scala 46:19:@12907.4]
  wire [7:0] _T_17396; // @[Mux.scala 46:16:@12908.4]
  wire  _T_17397; // @[Mux.scala 46:19:@12909.4]
  wire [7:0] _T_17398; // @[Mux.scala 46:16:@12910.4]
  wire  _T_17399; // @[Mux.scala 46:19:@12911.4]
  wire [7:0] _T_17400; // @[Mux.scala 46:16:@12912.4]
  wire  _T_17401; // @[Mux.scala 46:19:@12913.4]
  wire [7:0] _T_17402; // @[Mux.scala 46:16:@12914.4]
  wire  _T_17403; // @[Mux.scala 46:19:@12915.4]
  wire [7:0] _T_17404; // @[Mux.scala 46:16:@12916.4]
  wire  _T_17405; // @[Mux.scala 46:19:@12917.4]
  wire [7:0] _T_17406; // @[Mux.scala 46:16:@12918.4]
  wire  _T_17407; // @[Mux.scala 46:19:@12919.4]
  wire [7:0] _T_17408; // @[Mux.scala 46:16:@12920.4]
  wire  _T_17409; // @[Mux.scala 46:19:@12921.4]
  wire [7:0] _T_17410; // @[Mux.scala 46:16:@12922.4]
  wire  _T_17411; // @[Mux.scala 46:19:@12923.4]
  wire [7:0] _T_17412; // @[Mux.scala 46:16:@12924.4]
  wire  _T_17413; // @[Mux.scala 46:19:@12925.4]
  wire [7:0] _T_17414; // @[Mux.scala 46:16:@12926.4]
  wire  _T_17415; // @[Mux.scala 46:19:@12927.4]
  wire [7:0] _T_17416; // @[Mux.scala 46:16:@12928.4]
  wire  _T_17417; // @[Mux.scala 46:19:@12929.4]
  wire [7:0] _T_17418; // @[Mux.scala 46:16:@12930.4]
  wire  _T_17419; // @[Mux.scala 46:19:@12931.4]
  wire [7:0] _T_17420; // @[Mux.scala 46:16:@12932.4]
  wire  _T_17421; // @[Mux.scala 46:19:@12933.4]
  wire [7:0] _T_17422; // @[Mux.scala 46:16:@12934.4]
  wire  _T_17423; // @[Mux.scala 46:19:@12935.4]
  wire [7:0] _T_17424; // @[Mux.scala 46:16:@12936.4]
  wire  _T_17425; // @[Mux.scala 46:19:@12937.4]
  wire [7:0] _T_17426; // @[Mux.scala 46:16:@12938.4]
  wire  _T_17427; // @[Mux.scala 46:19:@12939.4]
  wire [7:0] _T_17428; // @[Mux.scala 46:16:@12940.4]
  wire  _T_17429; // @[Mux.scala 46:19:@12941.4]
  wire [7:0] _T_17430; // @[Mux.scala 46:16:@12942.4]
  wire  _T_17431; // @[Mux.scala 46:19:@12943.4]
  wire [7:0] _T_17432; // @[Mux.scala 46:16:@12944.4]
  wire  _T_17433; // @[Mux.scala 46:19:@12945.4]
  wire [7:0] _T_17434; // @[Mux.scala 46:16:@12946.4]
  wire  _T_17435; // @[Mux.scala 46:19:@12947.4]
  wire [7:0] _T_17436; // @[Mux.scala 46:16:@12948.4]
  wire  _T_17501; // @[Mux.scala 46:19:@12950.4]
  wire [7:0] _T_17502; // @[Mux.scala 46:16:@12951.4]
  wire  _T_17503; // @[Mux.scala 46:19:@12952.4]
  wire [7:0] _T_17504; // @[Mux.scala 46:16:@12953.4]
  wire  _T_17505; // @[Mux.scala 46:19:@12954.4]
  wire [7:0] _T_17506; // @[Mux.scala 46:16:@12955.4]
  wire  _T_17507; // @[Mux.scala 46:19:@12956.4]
  wire [7:0] _T_17508; // @[Mux.scala 46:16:@12957.4]
  wire  _T_17509; // @[Mux.scala 46:19:@12958.4]
  wire [7:0] _T_17510; // @[Mux.scala 46:16:@12959.4]
  wire  _T_17511; // @[Mux.scala 46:19:@12960.4]
  wire [7:0] _T_17512; // @[Mux.scala 46:16:@12961.4]
  wire  _T_17513; // @[Mux.scala 46:19:@12962.4]
  wire [7:0] _T_17514; // @[Mux.scala 46:16:@12963.4]
  wire  _T_17515; // @[Mux.scala 46:19:@12964.4]
  wire [7:0] _T_17516; // @[Mux.scala 46:16:@12965.4]
  wire  _T_17517; // @[Mux.scala 46:19:@12966.4]
  wire [7:0] _T_17518; // @[Mux.scala 46:16:@12967.4]
  wire  _T_17519; // @[Mux.scala 46:19:@12968.4]
  wire [7:0] _T_17520; // @[Mux.scala 46:16:@12969.4]
  wire  _T_17521; // @[Mux.scala 46:19:@12970.4]
  wire [7:0] _T_17522; // @[Mux.scala 46:16:@12971.4]
  wire  _T_17523; // @[Mux.scala 46:19:@12972.4]
  wire [7:0] _T_17524; // @[Mux.scala 46:16:@12973.4]
  wire  _T_17525; // @[Mux.scala 46:19:@12974.4]
  wire [7:0] _T_17526; // @[Mux.scala 46:16:@12975.4]
  wire  _T_17527; // @[Mux.scala 46:19:@12976.4]
  wire [7:0] _T_17528; // @[Mux.scala 46:16:@12977.4]
  wire  _T_17529; // @[Mux.scala 46:19:@12978.4]
  wire [7:0] _T_17530; // @[Mux.scala 46:16:@12979.4]
  wire  _T_17531; // @[Mux.scala 46:19:@12980.4]
  wire [7:0] _T_17532; // @[Mux.scala 46:16:@12981.4]
  wire  _T_17533; // @[Mux.scala 46:19:@12982.4]
  wire [7:0] _T_17534; // @[Mux.scala 46:16:@12983.4]
  wire  _T_17535; // @[Mux.scala 46:19:@12984.4]
  wire [7:0] _T_17536; // @[Mux.scala 46:16:@12985.4]
  wire  _T_17537; // @[Mux.scala 46:19:@12986.4]
  wire [7:0] _T_17538; // @[Mux.scala 46:16:@12987.4]
  wire  _T_17539; // @[Mux.scala 46:19:@12988.4]
  wire [7:0] _T_17540; // @[Mux.scala 46:16:@12989.4]
  wire  _T_17541; // @[Mux.scala 46:19:@12990.4]
  wire [7:0] _T_17542; // @[Mux.scala 46:16:@12991.4]
  wire  _T_17543; // @[Mux.scala 46:19:@12992.4]
  wire [7:0] _T_17544; // @[Mux.scala 46:16:@12993.4]
  wire  _T_17545; // @[Mux.scala 46:19:@12994.4]
  wire [7:0] _T_17546; // @[Mux.scala 46:16:@12995.4]
  wire  _T_17547; // @[Mux.scala 46:19:@12996.4]
  wire [7:0] _T_17548; // @[Mux.scala 46:16:@12997.4]
  wire  _T_17549; // @[Mux.scala 46:19:@12998.4]
  wire [7:0] _T_17550; // @[Mux.scala 46:16:@12999.4]
  wire  _T_17551; // @[Mux.scala 46:19:@13000.4]
  wire [7:0] _T_17552; // @[Mux.scala 46:16:@13001.4]
  wire  _T_17553; // @[Mux.scala 46:19:@13002.4]
  wire [7:0] _T_17554; // @[Mux.scala 46:16:@13003.4]
  wire  _T_17555; // @[Mux.scala 46:19:@13004.4]
  wire [7:0] _T_17556; // @[Mux.scala 46:16:@13005.4]
  wire  _T_17557; // @[Mux.scala 46:19:@13006.4]
  wire [7:0] _T_17558; // @[Mux.scala 46:16:@13007.4]
  wire  _T_17559; // @[Mux.scala 46:19:@13008.4]
  wire [7:0] _T_17560; // @[Mux.scala 46:16:@13009.4]
  wire  _T_17561; // @[Mux.scala 46:19:@13010.4]
  wire [7:0] _T_17562; // @[Mux.scala 46:16:@13011.4]
  wire  _T_17563; // @[Mux.scala 46:19:@13012.4]
  wire [7:0] _T_17564; // @[Mux.scala 46:16:@13013.4]
  wire  _T_17565; // @[Mux.scala 46:19:@13014.4]
  wire [7:0] _T_17566; // @[Mux.scala 46:16:@13015.4]
  wire  _T_17567; // @[Mux.scala 46:19:@13016.4]
  wire [7:0] _T_17568; // @[Mux.scala 46:16:@13017.4]
  wire  _T_17569; // @[Mux.scala 46:19:@13018.4]
  wire [7:0] _T_17570; // @[Mux.scala 46:16:@13019.4]
  wire  _T_17571; // @[Mux.scala 46:19:@13020.4]
  wire [7:0] _T_17572; // @[Mux.scala 46:16:@13021.4]
  wire  _T_17573; // @[Mux.scala 46:19:@13022.4]
  wire [7:0] _T_17574; // @[Mux.scala 46:16:@13023.4]
  wire  _T_17575; // @[Mux.scala 46:19:@13024.4]
  wire [7:0] _T_17576; // @[Mux.scala 46:16:@13025.4]
  wire  _T_17577; // @[Mux.scala 46:19:@13026.4]
  wire [7:0] _T_17578; // @[Mux.scala 46:16:@13027.4]
  wire  _T_17579; // @[Mux.scala 46:19:@13028.4]
  wire [7:0] _T_17580; // @[Mux.scala 46:16:@13029.4]
  wire  _T_17581; // @[Mux.scala 46:19:@13030.4]
  wire [7:0] _T_17582; // @[Mux.scala 46:16:@13031.4]
  wire  _T_17583; // @[Mux.scala 46:19:@13032.4]
  wire [7:0] _T_17584; // @[Mux.scala 46:16:@13033.4]
  wire  _T_17585; // @[Mux.scala 46:19:@13034.4]
  wire [7:0] _T_17586; // @[Mux.scala 46:16:@13035.4]
  wire  _T_17587; // @[Mux.scala 46:19:@13036.4]
  wire [7:0] _T_17588; // @[Mux.scala 46:16:@13037.4]
  wire  _T_17589; // @[Mux.scala 46:19:@13038.4]
  wire [7:0] _T_17590; // @[Mux.scala 46:16:@13039.4]
  wire  _T_17591; // @[Mux.scala 46:19:@13040.4]
  wire [7:0] _T_17592; // @[Mux.scala 46:16:@13041.4]
  wire  _T_17593; // @[Mux.scala 46:19:@13042.4]
  wire [7:0] _T_17594; // @[Mux.scala 46:16:@13043.4]
  wire  _T_17595; // @[Mux.scala 46:19:@13044.4]
  wire [7:0] _T_17596; // @[Mux.scala 46:16:@13045.4]
  wire  _T_17597; // @[Mux.scala 46:19:@13046.4]
  wire [7:0] _T_17598; // @[Mux.scala 46:16:@13047.4]
  wire  _T_17599; // @[Mux.scala 46:19:@13048.4]
  wire [7:0] _T_17600; // @[Mux.scala 46:16:@13049.4]
  wire  _T_17601; // @[Mux.scala 46:19:@13050.4]
  wire [7:0] _T_17602; // @[Mux.scala 46:16:@13051.4]
  wire  _T_17603; // @[Mux.scala 46:19:@13052.4]
  wire [7:0] _T_17604; // @[Mux.scala 46:16:@13053.4]
  wire  _T_17605; // @[Mux.scala 46:19:@13054.4]
  wire [7:0] _T_17606; // @[Mux.scala 46:16:@13055.4]
  wire  _T_17607; // @[Mux.scala 46:19:@13056.4]
  wire [7:0] _T_17608; // @[Mux.scala 46:16:@13057.4]
  wire  _T_17609; // @[Mux.scala 46:19:@13058.4]
  wire [7:0] _T_17610; // @[Mux.scala 46:16:@13059.4]
  wire  _T_17611; // @[Mux.scala 46:19:@13060.4]
  wire [7:0] _T_17612; // @[Mux.scala 46:16:@13061.4]
  wire  _T_17613; // @[Mux.scala 46:19:@13062.4]
  wire [7:0] _T_17614; // @[Mux.scala 46:16:@13063.4]
  wire  _T_17615; // @[Mux.scala 46:19:@13064.4]
  wire [7:0] _T_17616; // @[Mux.scala 46:16:@13065.4]
  wire  _T_17617; // @[Mux.scala 46:19:@13066.4]
  wire [7:0] _T_17618; // @[Mux.scala 46:16:@13067.4]
  wire  _T_17619; // @[Mux.scala 46:19:@13068.4]
  wire [7:0] _T_17620; // @[Mux.scala 46:16:@13069.4]
  wire  _T_17621; // @[Mux.scala 46:19:@13070.4]
  wire [7:0] _T_17622; // @[Mux.scala 46:16:@13071.4]
  wire  _T_17623; // @[Mux.scala 46:19:@13072.4]
  wire [7:0] _T_17624; // @[Mux.scala 46:16:@13073.4]
  wire  _T_17625; // @[Mux.scala 46:19:@13074.4]
  wire [7:0] _T_17626; // @[Mux.scala 46:16:@13075.4]
  wire  _T_17692; // @[Mux.scala 46:19:@13077.4]
  wire [7:0] _T_17693; // @[Mux.scala 46:16:@13078.4]
  wire  _T_17694; // @[Mux.scala 46:19:@13079.4]
  wire [7:0] _T_17695; // @[Mux.scala 46:16:@13080.4]
  wire  _T_17696; // @[Mux.scala 46:19:@13081.4]
  wire [7:0] _T_17697; // @[Mux.scala 46:16:@13082.4]
  wire  _T_17698; // @[Mux.scala 46:19:@13083.4]
  wire [7:0] _T_17699; // @[Mux.scala 46:16:@13084.4]
  wire  _T_17700; // @[Mux.scala 46:19:@13085.4]
  wire [7:0] _T_17701; // @[Mux.scala 46:16:@13086.4]
  wire  _T_17702; // @[Mux.scala 46:19:@13087.4]
  wire [7:0] _T_17703; // @[Mux.scala 46:16:@13088.4]
  wire  _T_17704; // @[Mux.scala 46:19:@13089.4]
  wire [7:0] _T_17705; // @[Mux.scala 46:16:@13090.4]
  wire  _T_17706; // @[Mux.scala 46:19:@13091.4]
  wire [7:0] _T_17707; // @[Mux.scala 46:16:@13092.4]
  wire  _T_17708; // @[Mux.scala 46:19:@13093.4]
  wire [7:0] _T_17709; // @[Mux.scala 46:16:@13094.4]
  wire  _T_17710; // @[Mux.scala 46:19:@13095.4]
  wire [7:0] _T_17711; // @[Mux.scala 46:16:@13096.4]
  wire  _T_17712; // @[Mux.scala 46:19:@13097.4]
  wire [7:0] _T_17713; // @[Mux.scala 46:16:@13098.4]
  wire  _T_17714; // @[Mux.scala 46:19:@13099.4]
  wire [7:0] _T_17715; // @[Mux.scala 46:16:@13100.4]
  wire  _T_17716; // @[Mux.scala 46:19:@13101.4]
  wire [7:0] _T_17717; // @[Mux.scala 46:16:@13102.4]
  wire  _T_17718; // @[Mux.scala 46:19:@13103.4]
  wire [7:0] _T_17719; // @[Mux.scala 46:16:@13104.4]
  wire  _T_17720; // @[Mux.scala 46:19:@13105.4]
  wire [7:0] _T_17721; // @[Mux.scala 46:16:@13106.4]
  wire  _T_17722; // @[Mux.scala 46:19:@13107.4]
  wire [7:0] _T_17723; // @[Mux.scala 46:16:@13108.4]
  wire  _T_17724; // @[Mux.scala 46:19:@13109.4]
  wire [7:0] _T_17725; // @[Mux.scala 46:16:@13110.4]
  wire  _T_17726; // @[Mux.scala 46:19:@13111.4]
  wire [7:0] _T_17727; // @[Mux.scala 46:16:@13112.4]
  wire  _T_17728; // @[Mux.scala 46:19:@13113.4]
  wire [7:0] _T_17729; // @[Mux.scala 46:16:@13114.4]
  wire  _T_17730; // @[Mux.scala 46:19:@13115.4]
  wire [7:0] _T_17731; // @[Mux.scala 46:16:@13116.4]
  wire  _T_17732; // @[Mux.scala 46:19:@13117.4]
  wire [7:0] _T_17733; // @[Mux.scala 46:16:@13118.4]
  wire  _T_17734; // @[Mux.scala 46:19:@13119.4]
  wire [7:0] _T_17735; // @[Mux.scala 46:16:@13120.4]
  wire  _T_17736; // @[Mux.scala 46:19:@13121.4]
  wire [7:0] _T_17737; // @[Mux.scala 46:16:@13122.4]
  wire  _T_17738; // @[Mux.scala 46:19:@13123.4]
  wire [7:0] _T_17739; // @[Mux.scala 46:16:@13124.4]
  wire  _T_17740; // @[Mux.scala 46:19:@13125.4]
  wire [7:0] _T_17741; // @[Mux.scala 46:16:@13126.4]
  wire  _T_17742; // @[Mux.scala 46:19:@13127.4]
  wire [7:0] _T_17743; // @[Mux.scala 46:16:@13128.4]
  wire  _T_17744; // @[Mux.scala 46:19:@13129.4]
  wire [7:0] _T_17745; // @[Mux.scala 46:16:@13130.4]
  wire  _T_17746; // @[Mux.scala 46:19:@13131.4]
  wire [7:0] _T_17747; // @[Mux.scala 46:16:@13132.4]
  wire  _T_17748; // @[Mux.scala 46:19:@13133.4]
  wire [7:0] _T_17749; // @[Mux.scala 46:16:@13134.4]
  wire  _T_17750; // @[Mux.scala 46:19:@13135.4]
  wire [7:0] _T_17751; // @[Mux.scala 46:16:@13136.4]
  wire  _T_17752; // @[Mux.scala 46:19:@13137.4]
  wire [7:0] _T_17753; // @[Mux.scala 46:16:@13138.4]
  wire  _T_17754; // @[Mux.scala 46:19:@13139.4]
  wire [7:0] _T_17755; // @[Mux.scala 46:16:@13140.4]
  wire  _T_17756; // @[Mux.scala 46:19:@13141.4]
  wire [7:0] _T_17757; // @[Mux.scala 46:16:@13142.4]
  wire  _T_17758; // @[Mux.scala 46:19:@13143.4]
  wire [7:0] _T_17759; // @[Mux.scala 46:16:@13144.4]
  wire  _T_17760; // @[Mux.scala 46:19:@13145.4]
  wire [7:0] _T_17761; // @[Mux.scala 46:16:@13146.4]
  wire  _T_17762; // @[Mux.scala 46:19:@13147.4]
  wire [7:0] _T_17763; // @[Mux.scala 46:16:@13148.4]
  wire  _T_17764; // @[Mux.scala 46:19:@13149.4]
  wire [7:0] _T_17765; // @[Mux.scala 46:16:@13150.4]
  wire  _T_17766; // @[Mux.scala 46:19:@13151.4]
  wire [7:0] _T_17767; // @[Mux.scala 46:16:@13152.4]
  wire  _T_17768; // @[Mux.scala 46:19:@13153.4]
  wire [7:0] _T_17769; // @[Mux.scala 46:16:@13154.4]
  wire  _T_17770; // @[Mux.scala 46:19:@13155.4]
  wire [7:0] _T_17771; // @[Mux.scala 46:16:@13156.4]
  wire  _T_17772; // @[Mux.scala 46:19:@13157.4]
  wire [7:0] _T_17773; // @[Mux.scala 46:16:@13158.4]
  wire  _T_17774; // @[Mux.scala 46:19:@13159.4]
  wire [7:0] _T_17775; // @[Mux.scala 46:16:@13160.4]
  wire  _T_17776; // @[Mux.scala 46:19:@13161.4]
  wire [7:0] _T_17777; // @[Mux.scala 46:16:@13162.4]
  wire  _T_17778; // @[Mux.scala 46:19:@13163.4]
  wire [7:0] _T_17779; // @[Mux.scala 46:16:@13164.4]
  wire  _T_17780; // @[Mux.scala 46:19:@13165.4]
  wire [7:0] _T_17781; // @[Mux.scala 46:16:@13166.4]
  wire  _T_17782; // @[Mux.scala 46:19:@13167.4]
  wire [7:0] _T_17783; // @[Mux.scala 46:16:@13168.4]
  wire  _T_17784; // @[Mux.scala 46:19:@13169.4]
  wire [7:0] _T_17785; // @[Mux.scala 46:16:@13170.4]
  wire  _T_17786; // @[Mux.scala 46:19:@13171.4]
  wire [7:0] _T_17787; // @[Mux.scala 46:16:@13172.4]
  wire  _T_17788; // @[Mux.scala 46:19:@13173.4]
  wire [7:0] _T_17789; // @[Mux.scala 46:16:@13174.4]
  wire  _T_17790; // @[Mux.scala 46:19:@13175.4]
  wire [7:0] _T_17791; // @[Mux.scala 46:16:@13176.4]
  wire  _T_17792; // @[Mux.scala 46:19:@13177.4]
  wire [7:0] _T_17793; // @[Mux.scala 46:16:@13178.4]
  wire  _T_17794; // @[Mux.scala 46:19:@13179.4]
  wire [7:0] _T_17795; // @[Mux.scala 46:16:@13180.4]
  wire  _T_17796; // @[Mux.scala 46:19:@13181.4]
  wire [7:0] _T_17797; // @[Mux.scala 46:16:@13182.4]
  wire  _T_17798; // @[Mux.scala 46:19:@13183.4]
  wire [7:0] _T_17799; // @[Mux.scala 46:16:@13184.4]
  wire  _T_17800; // @[Mux.scala 46:19:@13185.4]
  wire [7:0] _T_17801; // @[Mux.scala 46:16:@13186.4]
  wire  _T_17802; // @[Mux.scala 46:19:@13187.4]
  wire [7:0] _T_17803; // @[Mux.scala 46:16:@13188.4]
  wire  _T_17804; // @[Mux.scala 46:19:@13189.4]
  wire [7:0] _T_17805; // @[Mux.scala 46:16:@13190.4]
  wire  _T_17806; // @[Mux.scala 46:19:@13191.4]
  wire [7:0] _T_17807; // @[Mux.scala 46:16:@13192.4]
  wire  _T_17808; // @[Mux.scala 46:19:@13193.4]
  wire [7:0] _T_17809; // @[Mux.scala 46:16:@13194.4]
  wire  _T_17810; // @[Mux.scala 46:19:@13195.4]
  wire [7:0] _T_17811; // @[Mux.scala 46:16:@13196.4]
  wire  _T_17812; // @[Mux.scala 46:19:@13197.4]
  wire [7:0] _T_17813; // @[Mux.scala 46:16:@13198.4]
  wire  _T_17814; // @[Mux.scala 46:19:@13199.4]
  wire [7:0] _T_17815; // @[Mux.scala 46:16:@13200.4]
  wire  _T_17816; // @[Mux.scala 46:19:@13201.4]
  wire [7:0] _T_17817; // @[Mux.scala 46:16:@13202.4]
  wire  _T_17818; // @[Mux.scala 46:19:@13203.4]
  wire [7:0] _T_17819; // @[Mux.scala 46:16:@13204.4]
  reg  _T_17822; // @[NV_NVDLA_CSC_WL_dec.scala 94:27:@13206.4]
  reg [31:0] _RAND_225;
  reg  _T_17961_0; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_226;
  reg  _T_17961_1; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_227;
  reg  _T_17961_2; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_228;
  reg  _T_17961_3; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_229;
  reg  _T_17961_4; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_230;
  reg  _T_17961_5; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_231;
  reg  _T_17961_6; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_232;
  reg  _T_17961_7; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_233;
  reg  _T_17961_8; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_234;
  reg  _T_17961_9; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_235;
  reg  _T_17961_10; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_236;
  reg  _T_17961_11; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_237;
  reg  _T_17961_12; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_238;
  reg  _T_17961_13; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_239;
  reg  _T_17961_14; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_240;
  reg  _T_17961_15; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_241;
  reg  _T_17961_16; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_242;
  reg  _T_17961_17; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_243;
  reg  _T_17961_18; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_244;
  reg  _T_17961_19; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_245;
  reg  _T_17961_20; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_246;
  reg  _T_17961_21; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_247;
  reg  _T_17961_22; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_248;
  reg  _T_17961_23; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_249;
  reg  _T_17961_24; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_250;
  reg  _T_17961_25; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_251;
  reg  _T_17961_26; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_252;
  reg  _T_17961_27; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_253;
  reg  _T_17961_28; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_254;
  reg  _T_17961_29; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_255;
  reg  _T_17961_30; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_256;
  reg  _T_17961_31; // @[NV_NVDLA_CSC_WL_dec.scala 95:25:@13240.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_18065_0; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_18065_1; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_18065_2; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_18065_3; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_18065_4; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_18065_5; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_18065_6; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_18065_7; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_18065_8; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_18065_9; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_18065_10; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_18065_11; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_18065_12; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_18065_13; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_18065_14; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_18065_15; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_18065_16; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_18065_17; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_18065_18; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_18065_19; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_18065_20; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_18065_21; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_18065_22; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_18065_23; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_281;
  reg [7:0] _T_18065_24; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_282;
  reg [7:0] _T_18065_25; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_283;
  reg [7:0] _T_18065_26; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_284;
  reg [7:0] _T_18065_27; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_285;
  reg [7:0] _T_18065_28; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_286;
  reg [7:0] _T_18065_29; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_287;
  reg [7:0] _T_18065_30; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_288;
  reg [7:0] _T_18065_31; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_289;
  reg [7:0] _T_18065_32; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_290;
  reg [7:0] _T_18065_33; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_291;
  reg [7:0] _T_18065_34; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_292;
  reg [7:0] _T_18065_35; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_293;
  reg [7:0] _T_18065_36; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_294;
  reg [7:0] _T_18065_37; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_295;
  reg [7:0] _T_18065_38; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_296;
  reg [7:0] _T_18065_39; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_297;
  reg [7:0] _T_18065_40; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_298;
  reg [7:0] _T_18065_41; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_299;
  reg [7:0] _T_18065_42; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_300;
  reg [7:0] _T_18065_43; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_301;
  reg [7:0] _T_18065_44; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_302;
  reg [7:0] _T_18065_45; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_303;
  reg [7:0] _T_18065_46; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_304;
  reg [7:0] _T_18065_47; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_305;
  reg [7:0] _T_18065_48; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_306;
  reg [7:0] _T_18065_49; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_307;
  reg [7:0] _T_18065_50; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_308;
  reg [7:0] _T_18065_51; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_309;
  reg [7:0] _T_18065_52; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_310;
  reg [7:0] _T_18065_53; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_311;
  reg [7:0] _T_18065_54; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_312;
  reg [7:0] _T_18065_55; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_313;
  reg [7:0] _T_18065_56; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_314;
  reg [7:0] _T_18065_57; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_315;
  reg [7:0] _T_18065_58; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_316;
  reg [7:0] _T_18065_59; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_317;
  reg [7:0] _T_18065_60; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_318;
  reg [7:0] _T_18065_61; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_319;
  reg [7:0] _T_18065_62; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_320;
  reg [7:0] _T_18065_63; // @[NV_NVDLA_CSC_WL_dec.scala 96:26:@13241.4]
  reg [31:0] _RAND_321;
  wire  _GEN_224; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_230; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_231; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_232; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_233; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_234; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_235; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_236; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_237; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_238; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_239; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_240; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_241; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_242; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_243; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_244; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_245; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_246; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_247; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_248; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_249; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_250; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_251; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_252; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_253; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_254; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire  _GEN_255; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  wire [7:0] _GEN_256; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13278.6]
  wire [7:0] _GEN_258; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13286.6]
  wire [7:0] _GEN_260; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13294.6]
  wire [7:0] _GEN_262; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13302.6]
  wire [7:0] _GEN_264; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13310.6]
  wire [7:0] _GEN_266; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13318.6]
  wire [7:0] _GEN_268; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13326.6]
  wire [7:0] _GEN_270; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13334.6]
  wire [7:0] _GEN_272; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13342.6]
  wire [7:0] _GEN_274; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13350.6]
  wire [7:0] _GEN_276; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13358.6]
  wire [7:0] _GEN_278; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13366.6]
  wire [7:0] _GEN_280; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13374.6]
  wire [7:0] _GEN_282; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13382.6]
  wire [7:0] _GEN_284; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13390.6]
  wire [7:0] _GEN_286; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13398.6]
  wire [7:0] _GEN_288; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13406.6]
  wire [7:0] _GEN_290; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13414.6]
  wire [7:0] _GEN_292; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13422.6]
  wire [7:0] _GEN_294; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13430.6]
  wire [7:0] _GEN_296; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13438.6]
  wire [7:0] _GEN_298; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13446.6]
  wire [7:0] _GEN_300; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13454.6]
  wire [7:0] _GEN_302; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13462.6]
  wire [7:0] _GEN_304; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13470.6]
  wire [7:0] _GEN_306; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13478.6]
  wire [7:0] _GEN_308; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13486.6]
  wire [7:0] _GEN_310; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13494.6]
  wire [7:0] _GEN_312; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13502.6]
  wire [7:0] _GEN_314; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13510.6]
  wire [7:0] _GEN_316; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13518.6]
  wire [7:0] _GEN_318; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13526.6]
  wire [7:0] _GEN_320; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13534.6]
  wire [7:0] _GEN_322; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13542.6]
  wire [7:0] _GEN_324; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13550.6]
  wire [7:0] _GEN_326; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13558.6]
  wire [7:0] _GEN_328; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13566.6]
  wire [7:0] _GEN_330; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13574.6]
  wire [7:0] _GEN_332; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13582.6]
  wire [7:0] _GEN_334; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13590.6]
  wire [7:0] _GEN_336; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13598.6]
  wire [7:0] _GEN_338; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13606.6]
  wire [7:0] _GEN_340; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13614.6]
  wire [7:0] _GEN_342; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13622.6]
  wire [7:0] _GEN_344; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13630.6]
  wire [7:0] _GEN_346; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13638.6]
  wire [7:0] _GEN_348; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13646.6]
  wire [7:0] _GEN_350; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13654.6]
  wire [7:0] _GEN_352; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13662.6]
  wire [7:0] _GEN_354; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13670.6]
  wire [7:0] _GEN_356; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13678.6]
  wire [7:0] _GEN_358; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13686.6]
  wire [7:0] _GEN_360; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13694.6]
  wire [7:0] _GEN_362; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13702.6]
  wire [7:0] _GEN_364; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13710.6]
  wire [7:0] _GEN_366; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13718.6]
  wire [7:0] _GEN_368; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13726.6]
  wire [7:0] _GEN_370; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13734.6]
  wire [7:0] _GEN_372; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13742.6]
  wire [7:0] _GEN_374; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13750.6]
  wire [7:0] _GEN_376; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13758.6]
  wire [7:0] _GEN_378; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13766.6]
  wire [7:0] _GEN_380; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13774.6]
  wire [7:0] _GEN_382; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13782.6]
  wire  _T_18267; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13790.4]
  wire  _T_18269; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13792.4]
  wire  _T_18271; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13794.4]
  wire  _T_18273; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13796.4]
  wire  _T_18275; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13798.4]
  wire  _T_18277; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13800.4]
  wire  _T_18279; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13802.4]
  wire  _T_18281; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13804.4]
  wire  _T_18283; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13806.4]
  wire  _T_18285; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13808.4]
  wire  _T_18287; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13810.4]
  wire  _T_18289; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13812.4]
  wire  _T_18291; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13814.4]
  wire  _T_18293; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13816.4]
  wire  _T_18295; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13818.4]
  wire  _T_18297; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13820.4]
  wire  _T_18299; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13822.4]
  wire  _T_18301; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13824.4]
  wire  _T_18303; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13826.4]
  wire  _T_18305; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13828.4]
  wire  _T_18307; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13830.4]
  wire  _T_18309; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13832.4]
  wire  _T_18311; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13834.4]
  wire  _T_18313; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13836.4]
  wire  _T_18315; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13838.4]
  wire  _T_18317; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13840.4]
  wire  _T_18319; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13842.4]
  wire  _T_18321; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13844.4]
  wire  _T_18323; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13846.4]
  wire  _T_18325; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13848.4]
  wire  _T_18327; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13850.4]
  wire  _T_18329; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13852.4]
  wire  _T_18331; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13854.4]
  wire  _T_18333; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13856.4]
  wire  _T_18335; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13858.4]
  wire  _T_18337; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13860.4]
  wire  _T_18339; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13862.4]
  wire  _T_18341; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13864.4]
  wire  _T_18343; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13866.4]
  wire  _T_18345; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13868.4]
  wire  _T_18347; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13870.4]
  wire  _T_18349; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13872.4]
  wire  _T_18351; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13874.4]
  wire  _T_18353; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13876.4]
  wire  _T_18355; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13878.4]
  wire  _T_18357; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13880.4]
  wire  _T_18359; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13882.4]
  wire  _T_18361; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13884.4]
  wire  _T_18363; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13886.4]
  wire  _T_18365; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13888.4]
  wire  _T_18367; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13890.4]
  wire  _T_18369; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13892.4]
  wire  _T_18371; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13894.4]
  wire  _T_18373; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13896.4]
  wire  _T_18375; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13898.4]
  wire  _T_18377; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13900.4]
  wire  _T_18379; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13902.4]
  wire  _T_18381; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13904.4]
  wire  _T_18383; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13906.4]
  wire  _T_18385; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13908.4]
  wire  _T_18387; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13910.4]
  wire  _T_18389; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13912.4]
  wire  _T_18391; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13914.4]
  wire  _T_18393; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13916.4]
  reg  _T_18396; // @[NV_NVDLA_CSC_WL_dec.scala 122:27:@13918.4]
  reg [31:0] _RAND_322;
  reg  _T_18400_0; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_323;
  reg  _T_18400_1; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_324;
  reg  _T_18400_2; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_325;
  reg  _T_18400_3; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_326;
  reg  _T_18400_4; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_327;
  reg  _T_18400_5; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_328;
  reg  _T_18400_6; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_329;
  reg  _T_18400_7; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_330;
  reg  _T_18400_8; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_331;
  reg  _T_18400_9; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_332;
  reg  _T_18400_10; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_333;
  reg  _T_18400_11; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_334;
  reg  _T_18400_12; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_335;
  reg  _T_18400_13; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_336;
  reg  _T_18400_14; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_337;
  reg  _T_18400_15; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_338;
  reg  _T_18400_16; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_339;
  reg  _T_18400_17; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_340;
  reg  _T_18400_18; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_341;
  reg  _T_18400_19; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_342;
  reg  _T_18400_20; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_343;
  reg  _T_18400_21; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_344;
  reg  _T_18400_22; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_345;
  reg  _T_18400_23; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_346;
  reg  _T_18400_24; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_347;
  reg  _T_18400_25; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_348;
  reg  _T_18400_26; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_349;
  reg  _T_18400_27; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_350;
  reg  _T_18400_28; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_351;
  reg  _T_18400_29; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_352;
  reg  _T_18400_30; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_353;
  reg  _T_18400_31; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_354;
  reg  _T_18400_32; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_355;
  reg  _T_18400_33; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_356;
  reg  _T_18400_34; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_357;
  reg  _T_18400_35; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_358;
  reg  _T_18400_36; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_359;
  reg  _T_18400_37; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_360;
  reg  _T_18400_38; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_361;
  reg  _T_18400_39; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_362;
  reg  _T_18400_40; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_363;
  reg  _T_18400_41; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_364;
  reg  _T_18400_42; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_365;
  reg  _T_18400_43; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_366;
  reg  _T_18400_44; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_367;
  reg  _T_18400_45; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_368;
  reg  _T_18400_46; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_369;
  reg  _T_18400_47; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_370;
  reg  _T_18400_48; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_371;
  reg  _T_18400_49; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_372;
  reg  _T_18400_50; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_373;
  reg  _T_18400_51; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_374;
  reg  _T_18400_52; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_375;
  reg  _T_18400_53; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_376;
  reg  _T_18400_54; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_377;
  reg  _T_18400_55; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_378;
  reg  _T_18400_56; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_379;
  reg  _T_18400_57; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_380;
  reg  _T_18400_58; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_381;
  reg  _T_18400_59; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_382;
  reg  _T_18400_60; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_383;
  reg  _T_18400_61; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_384;
  reg  _T_18400_62; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_385;
  reg  _T_18400_63; // @[NV_NVDLA_CSC_WL_dec.scala 123:22:@13919.4]
  reg [31:0] _RAND_386;
  reg  _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_387;
  reg  _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_388;
  reg  _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_389;
  reg  _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_390;
  reg  _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_391;
  reg  _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_392;
  reg  _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_393;
  reg  _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_394;
  reg  _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_395;
  reg  _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_396;
  reg  _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_397;
  reg  _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_398;
  reg  _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_399;
  reg  _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_400;
  reg  _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_401;
  reg  _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_402;
  reg  _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_403;
  reg  _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_404;
  reg  _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_405;
  reg  _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_406;
  reg  _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_407;
  reg  _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_408;
  reg  _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_409;
  reg  _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_410;
  reg  _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_411;
  reg  _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_412;
  reg  _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_413;
  reg  _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_414;
  reg  _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_415;
  reg  _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_416;
  reg  _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_417;
  reg  _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 124:25:@13953.4]
  reg [31:0] _RAND_418;
  reg [7:0] _T_18709_0; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_419;
  reg [7:0] _T_18709_1; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_420;
  reg [7:0] _T_18709_2; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_421;
  reg [7:0] _T_18709_3; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_422;
  reg [7:0] _T_18709_4; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_423;
  reg [7:0] _T_18709_5; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_424;
  reg [7:0] _T_18709_6; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_425;
  reg [7:0] _T_18709_7; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_426;
  reg [7:0] _T_18709_8; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_427;
  reg [7:0] _T_18709_9; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_428;
  reg [7:0] _T_18709_10; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_429;
  reg [7:0] _T_18709_11; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_430;
  reg [7:0] _T_18709_12; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_431;
  reg [7:0] _T_18709_13; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_432;
  reg [7:0] _T_18709_14; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_433;
  reg [7:0] _T_18709_15; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_434;
  reg [7:0] _T_18709_16; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_435;
  reg [7:0] _T_18709_17; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_436;
  reg [7:0] _T_18709_18; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_437;
  reg [7:0] _T_18709_19; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_438;
  reg [7:0] _T_18709_20; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_439;
  reg [7:0] _T_18709_21; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_440;
  reg [7:0] _T_18709_22; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_441;
  reg [7:0] _T_18709_23; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_442;
  reg [7:0] _T_18709_24; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_443;
  reg [7:0] _T_18709_25; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_444;
  reg [7:0] _T_18709_26; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_445;
  reg [7:0] _T_18709_27; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_446;
  reg [7:0] _T_18709_28; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_447;
  reg [7:0] _T_18709_29; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_448;
  reg [7:0] _T_18709_30; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_449;
  reg [7:0] _T_18709_31; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_450;
  reg [7:0] _T_18709_32; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_451;
  reg [7:0] _T_18709_33; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_452;
  reg [7:0] _T_18709_34; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_453;
  reg [7:0] _T_18709_35; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_454;
  reg [7:0] _T_18709_36; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_455;
  reg [7:0] _T_18709_37; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_456;
  reg [7:0] _T_18709_38; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_457;
  reg [7:0] _T_18709_39; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_458;
  reg [7:0] _T_18709_40; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_459;
  reg [7:0] _T_18709_41; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_460;
  reg [7:0] _T_18709_42; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_461;
  reg [7:0] _T_18709_43; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_462;
  reg [7:0] _T_18709_44; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_463;
  reg [7:0] _T_18709_45; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_464;
  reg [7:0] _T_18709_46; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_465;
  reg [7:0] _T_18709_47; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_466;
  reg [7:0] _T_18709_48; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_467;
  reg [7:0] _T_18709_49; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_468;
  reg [7:0] _T_18709_50; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_469;
  reg [7:0] _T_18709_51; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_470;
  reg [7:0] _T_18709_52; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_471;
  reg [7:0] _T_18709_53; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_472;
  reg [7:0] _T_18709_54; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_473;
  reg [7:0] _T_18709_55; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_474;
  reg [7:0] _T_18709_56; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_475;
  reg [7:0] _T_18709_57; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_476;
  reg [7:0] _T_18709_58; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_477;
  reg [7:0] _T_18709_59; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_478;
  reg [7:0] _T_18709_60; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_479;
  reg [7:0] _T_18709_61; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_480;
  reg [7:0] _T_18709_62; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_481;
  reg [7:0] _T_18709_63; // @[NV_NVDLA_CSC_WL_dec.scala 125:26:@13954.4]
  reg [31:0] _RAND_482;
  wire  _GEN_448; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_449; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_450; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_451; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_452; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_453; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_454; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_455; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_456; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_457; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_458; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_459; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_460; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_461; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_462; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_463; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_464; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_465; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_466; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_467; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_468; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_469; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_470; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_471; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_472; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_473; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_474; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_475; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_476; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_477; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_478; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  wire  _GEN_479; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _T_1771 = io_input_mask_en[8]; // @[NV_NVDLA_CSC_WL_dec.scala 56:48:@8.4]
  assign _T_1906_0 = _T_1771 ? io_input_bits_mask_0 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_1 = _T_1771 ? io_input_bits_mask_1 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_2 = _T_1771 ? io_input_bits_mask_2 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_3 = _T_1771 ? io_input_bits_mask_3 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_4 = _T_1771 ? io_input_bits_mask_4 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_5 = _T_1771 ? io_input_bits_mask_5 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_6 = _T_1771 ? io_input_bits_mask_6 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_7 = _T_1771 ? io_input_bits_mask_7 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_8 = _T_1771 ? io_input_bits_mask_8 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_9 = _T_1771 ? io_input_bits_mask_9 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_10 = _T_1771 ? io_input_bits_mask_10 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_11 = _T_1771 ? io_input_bits_mask_11 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_12 = _T_1771 ? io_input_bits_mask_12 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_13 = _T_1771 ? io_input_bits_mask_13 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_14 = _T_1771 ? io_input_bits_mask_14 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_15 = _T_1771 ? io_input_bits_mask_15 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_16 = _T_1771 ? io_input_bits_mask_16 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_17 = _T_1771 ? io_input_bits_mask_17 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_18 = _T_1771 ? io_input_bits_mask_18 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_19 = _T_1771 ? io_input_bits_mask_19 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_20 = _T_1771 ? io_input_bits_mask_20 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_21 = _T_1771 ? io_input_bits_mask_21 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_22 = _T_1771 ? io_input_bits_mask_22 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_23 = _T_1771 ? io_input_bits_mask_23 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_24 = _T_1771 ? io_input_bits_mask_24 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_25 = _T_1771 ? io_input_bits_mask_25 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_26 = _T_1771 ? io_input_bits_mask_26 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_27 = _T_1771 ? io_input_bits_mask_27 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_28 = _T_1771 ? io_input_bits_mask_28 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_29 = _T_1771 ? io_input_bits_mask_29 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_30 = _T_1771 ? io_input_bits_mask_30 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_31 = _T_1771 ? io_input_bits_mask_31 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_32 = _T_1771 ? io_input_bits_mask_32 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_33 = _T_1771 ? io_input_bits_mask_33 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_34 = _T_1771 ? io_input_bits_mask_34 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_35 = _T_1771 ? io_input_bits_mask_35 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_36 = _T_1771 ? io_input_bits_mask_36 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_37 = _T_1771 ? io_input_bits_mask_37 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_38 = _T_1771 ? io_input_bits_mask_38 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_39 = _T_1771 ? io_input_bits_mask_39 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_40 = _T_1771 ? io_input_bits_mask_40 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_41 = _T_1771 ? io_input_bits_mask_41 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_42 = _T_1771 ? io_input_bits_mask_42 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_43 = _T_1771 ? io_input_bits_mask_43 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_44 = _T_1771 ? io_input_bits_mask_44 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_45 = _T_1771 ? io_input_bits_mask_45 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_46 = _T_1771 ? io_input_bits_mask_46 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_47 = _T_1771 ? io_input_bits_mask_47 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_48 = _T_1771 ? io_input_bits_mask_48 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_49 = _T_1771 ? io_input_bits_mask_49 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_50 = _T_1771 ? io_input_bits_mask_50 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_51 = _T_1771 ? io_input_bits_mask_51 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_52 = _T_1771 ? io_input_bits_mask_52 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_53 = _T_1771 ? io_input_bits_mask_53 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_54 = _T_1771 ? io_input_bits_mask_54 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_55 = _T_1771 ? io_input_bits_mask_55 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_56 = _T_1771 ? io_input_bits_mask_56 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_57 = _T_1771 ? io_input_bits_mask_57 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_58 = _T_1771 ? io_input_bits_mask_58 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_59 = _T_1771 ? io_input_bits_mask_59 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_60 = _T_1771 ? io_input_bits_mask_60 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_61 = _T_1771 ? io_input_bits_mask_61 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_62 = _T_1771 ? io_input_bits_mask_62 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_1906_63 = _T_1771 ? io_input_bits_mask_63 : 1'h0; // @[NV_NVDLA_CSC_WL_dec.scala 56:31:@74.4]
  assign _T_2174 = {_T_1906_7,_T_1906_6,_T_1906_5,_T_1906_4,_T_1906_3,_T_1906_2,_T_1906_1,_T_1906_0}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@82.4]
  assign _T_2182 = {_T_1906_15,_T_1906_14,_T_1906_13,_T_1906_12,_T_1906_11,_T_1906_10,_T_1906_9,_T_1906_8,_T_2174}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@90.4]
  assign _T_2189 = {_T_1906_23,_T_1906_22,_T_1906_21,_T_1906_20,_T_1906_19,_T_1906_18,_T_1906_17,_T_1906_16}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@97.4]
  assign _T_2198 = {_T_1906_31,_T_1906_30,_T_1906_29,_T_1906_28,_T_1906_27,_T_1906_26,_T_1906_25,_T_1906_24,_T_2189,_T_2182}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@106.4]
  assign _T_2205 = {_T_1906_39,_T_1906_38,_T_1906_37,_T_1906_36,_T_1906_35,_T_1906_34,_T_1906_33,_T_1906_32}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@113.4]
  assign _T_2213 = {_T_1906_47,_T_1906_46,_T_1906_45,_T_1906_44,_T_1906_43,_T_1906_42,_T_1906_41,_T_1906_40,_T_2205}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@121.4]
  assign _T_2220 = {_T_1906_55,_T_1906_54,_T_1906_53,_T_1906_52,_T_1906_51,_T_1906_50,_T_1906_49,_T_1906_48}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@128.4]
  assign _T_2229 = {_T_1906_63,_T_1906_62,_T_1906_61,_T_1906_60,_T_1906_59,_T_1906_58,_T_1906_57,_T_1906_56,_T_2220,_T_2213}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@137.4]
  assign _T_2230 = {_T_2229,_T_2198}; // @[NV_NVDLA_CSC_WL_dec.scala 60:53:@138.4]
  assign _T_2231 = _T_2230[0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@139.4]
  assign _T_2296 = _T_2230[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@205.4]
  assign _T_2297 = _T_2296[0]; // @[Bitwise.scala 50:65:@206.4]
  assign _T_2298 = _T_2296[1]; // @[Bitwise.scala 50:65:@207.4]
  assign _T_2299 = _T_2297 + _T_2298; // @[Bitwise.scala 48:55:@208.4]
  assign _T_2363 = _T_2230[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@273.4]
  assign _T_2364 = _T_2363[0]; // @[Bitwise.scala 50:65:@274.4]
  assign _T_2365 = _T_2363[1]; // @[Bitwise.scala 50:65:@275.4]
  assign _T_2366 = _T_2363[2]; // @[Bitwise.scala 50:65:@276.4]
  assign _T_2367 = _T_2365 + _T_2366; // @[Bitwise.scala 48:55:@277.4]
  assign _GEN_544 = {{1'd0}, _T_2364}; // @[Bitwise.scala 48:55:@278.4]
  assign _T_2368 = _GEN_544 + _T_2367; // @[Bitwise.scala 48:55:@278.4]
  assign _T_2432 = _T_2230[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@343.4]
  assign _T_2433 = _T_2432[0]; // @[Bitwise.scala 50:65:@344.4]
  assign _T_2434 = _T_2432[1]; // @[Bitwise.scala 50:65:@345.4]
  assign _T_2435 = _T_2432[2]; // @[Bitwise.scala 50:65:@346.4]
  assign _T_2436 = _T_2432[3]; // @[Bitwise.scala 50:65:@347.4]
  assign _T_2437 = _T_2433 + _T_2434; // @[Bitwise.scala 48:55:@348.4]
  assign _T_2438 = _T_2435 + _T_2436; // @[Bitwise.scala 48:55:@349.4]
  assign _T_2439 = _T_2437 + _T_2438; // @[Bitwise.scala 48:55:@350.4]
  assign _T_2503 = _T_2230[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@415.4]
  assign _T_2504 = _T_2503[0]; // @[Bitwise.scala 50:65:@416.4]
  assign _T_2505 = _T_2503[1]; // @[Bitwise.scala 50:65:@417.4]
  assign _T_2506 = _T_2503[2]; // @[Bitwise.scala 50:65:@418.4]
  assign _T_2507 = _T_2503[3]; // @[Bitwise.scala 50:65:@419.4]
  assign _T_2508 = _T_2503[4]; // @[Bitwise.scala 50:65:@420.4]
  assign _T_2509 = _T_2504 + _T_2505; // @[Bitwise.scala 48:55:@421.4]
  assign _T_2510 = _T_2507 + _T_2508; // @[Bitwise.scala 48:55:@422.4]
  assign _GEN_545 = {{1'd0}, _T_2506}; // @[Bitwise.scala 48:55:@423.4]
  assign _T_2511 = _GEN_545 + _T_2510; // @[Bitwise.scala 48:55:@423.4]
  assign _GEN_546 = {{1'd0}, _T_2509}; // @[Bitwise.scala 48:55:@424.4]
  assign _T_2512 = _GEN_546 + _T_2511; // @[Bitwise.scala 48:55:@424.4]
  assign _T_2576 = _T_2230[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@489.4]
  assign _T_2577 = _T_2576[0]; // @[Bitwise.scala 50:65:@490.4]
  assign _T_2578 = _T_2576[1]; // @[Bitwise.scala 50:65:@491.4]
  assign _T_2579 = _T_2576[2]; // @[Bitwise.scala 50:65:@492.4]
  assign _T_2580 = _T_2576[3]; // @[Bitwise.scala 50:65:@493.4]
  assign _T_2581 = _T_2576[4]; // @[Bitwise.scala 50:65:@494.4]
  assign _T_2582 = _T_2576[5]; // @[Bitwise.scala 50:65:@495.4]
  assign _T_2583 = _T_2578 + _T_2579; // @[Bitwise.scala 48:55:@496.4]
  assign _GEN_547 = {{1'd0}, _T_2577}; // @[Bitwise.scala 48:55:@497.4]
  assign _T_2584 = _GEN_547 + _T_2583; // @[Bitwise.scala 48:55:@497.4]
  assign _T_2585 = _T_2581 + _T_2582; // @[Bitwise.scala 48:55:@498.4]
  assign _GEN_548 = {{1'd0}, _T_2580}; // @[Bitwise.scala 48:55:@499.4]
  assign _T_2586 = _GEN_548 + _T_2585; // @[Bitwise.scala 48:55:@499.4]
  assign _T_2587 = _T_2584 + _T_2586; // @[Bitwise.scala 48:55:@500.4]
  assign _T_2651 = _T_2230[6:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@565.4]
  assign _T_2652 = _T_2651[0]; // @[Bitwise.scala 50:65:@566.4]
  assign _T_2653 = _T_2651[1]; // @[Bitwise.scala 50:65:@567.4]
  assign _T_2654 = _T_2651[2]; // @[Bitwise.scala 50:65:@568.4]
  assign _T_2655 = _T_2651[3]; // @[Bitwise.scala 50:65:@569.4]
  assign _T_2656 = _T_2651[4]; // @[Bitwise.scala 50:65:@570.4]
  assign _T_2657 = _T_2651[5]; // @[Bitwise.scala 50:65:@571.4]
  assign _T_2658 = _T_2651[6]; // @[Bitwise.scala 50:65:@572.4]
  assign _T_2659 = _T_2653 + _T_2654; // @[Bitwise.scala 48:55:@573.4]
  assign _GEN_549 = {{1'd0}, _T_2652}; // @[Bitwise.scala 48:55:@574.4]
  assign _T_2660 = _GEN_549 + _T_2659; // @[Bitwise.scala 48:55:@574.4]
  assign _T_2661 = _T_2655 + _T_2656; // @[Bitwise.scala 48:55:@575.4]
  assign _T_2662 = _T_2657 + _T_2658; // @[Bitwise.scala 48:55:@576.4]
  assign _T_2663 = _T_2661 + _T_2662; // @[Bitwise.scala 48:55:@577.4]
  assign _T_2664 = _T_2660 + _T_2663; // @[Bitwise.scala 48:55:@578.4]
  assign _T_2728 = _T_2230[7:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@643.4]
  assign _T_2729 = _T_2728[0]; // @[Bitwise.scala 50:65:@644.4]
  assign _T_2730 = _T_2728[1]; // @[Bitwise.scala 50:65:@645.4]
  assign _T_2731 = _T_2728[2]; // @[Bitwise.scala 50:65:@646.4]
  assign _T_2732 = _T_2728[3]; // @[Bitwise.scala 50:65:@647.4]
  assign _T_2733 = _T_2728[4]; // @[Bitwise.scala 50:65:@648.4]
  assign _T_2734 = _T_2728[5]; // @[Bitwise.scala 50:65:@649.4]
  assign _T_2735 = _T_2728[6]; // @[Bitwise.scala 50:65:@650.4]
  assign _T_2736 = _T_2728[7]; // @[Bitwise.scala 50:65:@651.4]
  assign _T_2737 = _T_2729 + _T_2730; // @[Bitwise.scala 48:55:@652.4]
  assign _T_2738 = _T_2731 + _T_2732; // @[Bitwise.scala 48:55:@653.4]
  assign _T_2739 = _T_2737 + _T_2738; // @[Bitwise.scala 48:55:@654.4]
  assign _T_2740 = _T_2733 + _T_2734; // @[Bitwise.scala 48:55:@655.4]
  assign _T_2741 = _T_2735 + _T_2736; // @[Bitwise.scala 48:55:@656.4]
  assign _T_2742 = _T_2740 + _T_2741; // @[Bitwise.scala 48:55:@657.4]
  assign _T_2743 = _T_2739 + _T_2742; // @[Bitwise.scala 48:55:@658.4]
  assign _T_2807 = _T_2230[8:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@723.4]
  assign _T_2808 = _T_2807[0]; // @[Bitwise.scala 50:65:@724.4]
  assign _T_2809 = _T_2807[1]; // @[Bitwise.scala 50:65:@725.4]
  assign _T_2810 = _T_2807[2]; // @[Bitwise.scala 50:65:@726.4]
  assign _T_2811 = _T_2807[3]; // @[Bitwise.scala 50:65:@727.4]
  assign _T_2812 = _T_2807[4]; // @[Bitwise.scala 50:65:@728.4]
  assign _T_2813 = _T_2807[5]; // @[Bitwise.scala 50:65:@729.4]
  assign _T_2814 = _T_2807[6]; // @[Bitwise.scala 50:65:@730.4]
  assign _T_2815 = _T_2807[7]; // @[Bitwise.scala 50:65:@731.4]
  assign _T_2816 = _T_2807[8]; // @[Bitwise.scala 50:65:@732.4]
  assign _T_2817 = _T_2808 + _T_2809; // @[Bitwise.scala 48:55:@733.4]
  assign _T_2818 = _T_2810 + _T_2811; // @[Bitwise.scala 48:55:@734.4]
  assign _T_2819 = _T_2817 + _T_2818; // @[Bitwise.scala 48:55:@735.4]
  assign _T_2820 = _T_2812 + _T_2813; // @[Bitwise.scala 48:55:@736.4]
  assign _T_2821 = _T_2815 + _T_2816; // @[Bitwise.scala 48:55:@737.4]
  assign _GEN_550 = {{1'd0}, _T_2814}; // @[Bitwise.scala 48:55:@738.4]
  assign _T_2822 = _GEN_550 + _T_2821; // @[Bitwise.scala 48:55:@738.4]
  assign _GEN_551 = {{1'd0}, _T_2820}; // @[Bitwise.scala 48:55:@739.4]
  assign _T_2823 = _GEN_551 + _T_2822; // @[Bitwise.scala 48:55:@739.4]
  assign _GEN_552 = {{1'd0}, _T_2819}; // @[Bitwise.scala 48:55:@740.4]
  assign _T_2824 = _GEN_552 + _T_2823; // @[Bitwise.scala 48:55:@740.4]
  assign _T_2888 = _T_2230[9:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@805.4]
  assign _T_2889 = _T_2888[0]; // @[Bitwise.scala 50:65:@806.4]
  assign _T_2890 = _T_2888[1]; // @[Bitwise.scala 50:65:@807.4]
  assign _T_2891 = _T_2888[2]; // @[Bitwise.scala 50:65:@808.4]
  assign _T_2892 = _T_2888[3]; // @[Bitwise.scala 50:65:@809.4]
  assign _T_2893 = _T_2888[4]; // @[Bitwise.scala 50:65:@810.4]
  assign _T_2894 = _T_2888[5]; // @[Bitwise.scala 50:65:@811.4]
  assign _T_2895 = _T_2888[6]; // @[Bitwise.scala 50:65:@812.4]
  assign _T_2896 = _T_2888[7]; // @[Bitwise.scala 50:65:@813.4]
  assign _T_2897 = _T_2888[8]; // @[Bitwise.scala 50:65:@814.4]
  assign _T_2898 = _T_2888[9]; // @[Bitwise.scala 50:65:@815.4]
  assign _T_2899 = _T_2889 + _T_2890; // @[Bitwise.scala 48:55:@816.4]
  assign _T_2900 = _T_2892 + _T_2893; // @[Bitwise.scala 48:55:@817.4]
  assign _GEN_553 = {{1'd0}, _T_2891}; // @[Bitwise.scala 48:55:@818.4]
  assign _T_2901 = _GEN_553 + _T_2900; // @[Bitwise.scala 48:55:@818.4]
  assign _GEN_554 = {{1'd0}, _T_2899}; // @[Bitwise.scala 48:55:@819.4]
  assign _T_2902 = _GEN_554 + _T_2901; // @[Bitwise.scala 48:55:@819.4]
  assign _T_2903 = _T_2894 + _T_2895; // @[Bitwise.scala 48:55:@820.4]
  assign _T_2904 = _T_2897 + _T_2898; // @[Bitwise.scala 48:55:@821.4]
  assign _GEN_555 = {{1'd0}, _T_2896}; // @[Bitwise.scala 48:55:@822.4]
  assign _T_2905 = _GEN_555 + _T_2904; // @[Bitwise.scala 48:55:@822.4]
  assign _GEN_556 = {{1'd0}, _T_2903}; // @[Bitwise.scala 48:55:@823.4]
  assign _T_2906 = _GEN_556 + _T_2905; // @[Bitwise.scala 48:55:@823.4]
  assign _T_2907 = _T_2902 + _T_2906; // @[Bitwise.scala 48:55:@824.4]
  assign _T_2971 = _T_2230[10:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@889.4]
  assign _T_2972 = _T_2971[0]; // @[Bitwise.scala 50:65:@890.4]
  assign _T_2973 = _T_2971[1]; // @[Bitwise.scala 50:65:@891.4]
  assign _T_2974 = _T_2971[2]; // @[Bitwise.scala 50:65:@892.4]
  assign _T_2975 = _T_2971[3]; // @[Bitwise.scala 50:65:@893.4]
  assign _T_2976 = _T_2971[4]; // @[Bitwise.scala 50:65:@894.4]
  assign _T_2977 = _T_2971[5]; // @[Bitwise.scala 50:65:@895.4]
  assign _T_2978 = _T_2971[6]; // @[Bitwise.scala 50:65:@896.4]
  assign _T_2979 = _T_2971[7]; // @[Bitwise.scala 50:65:@897.4]
  assign _T_2980 = _T_2971[8]; // @[Bitwise.scala 50:65:@898.4]
  assign _T_2981 = _T_2971[9]; // @[Bitwise.scala 50:65:@899.4]
  assign _T_2982 = _T_2971[10]; // @[Bitwise.scala 50:65:@900.4]
  assign _T_2983 = _T_2972 + _T_2973; // @[Bitwise.scala 48:55:@901.4]
  assign _T_2984 = _T_2975 + _T_2976; // @[Bitwise.scala 48:55:@902.4]
  assign _GEN_557 = {{1'd0}, _T_2974}; // @[Bitwise.scala 48:55:@903.4]
  assign _T_2985 = _GEN_557 + _T_2984; // @[Bitwise.scala 48:55:@903.4]
  assign _GEN_558 = {{1'd0}, _T_2983}; // @[Bitwise.scala 48:55:@904.4]
  assign _T_2986 = _GEN_558 + _T_2985; // @[Bitwise.scala 48:55:@904.4]
  assign _T_2987 = _T_2978 + _T_2979; // @[Bitwise.scala 48:55:@905.4]
  assign _GEN_559 = {{1'd0}, _T_2977}; // @[Bitwise.scala 48:55:@906.4]
  assign _T_2988 = _GEN_559 + _T_2987; // @[Bitwise.scala 48:55:@906.4]
  assign _T_2989 = _T_2981 + _T_2982; // @[Bitwise.scala 48:55:@907.4]
  assign _GEN_560 = {{1'd0}, _T_2980}; // @[Bitwise.scala 48:55:@908.4]
  assign _T_2990 = _GEN_560 + _T_2989; // @[Bitwise.scala 48:55:@908.4]
  assign _T_2991 = _T_2988 + _T_2990; // @[Bitwise.scala 48:55:@909.4]
  assign _T_2992 = _T_2986 + _T_2991; // @[Bitwise.scala 48:55:@910.4]
  assign _T_3056 = _T_2230[11:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@975.4]
  assign _T_3057 = _T_3056[0]; // @[Bitwise.scala 50:65:@976.4]
  assign _T_3058 = _T_3056[1]; // @[Bitwise.scala 50:65:@977.4]
  assign _T_3059 = _T_3056[2]; // @[Bitwise.scala 50:65:@978.4]
  assign _T_3060 = _T_3056[3]; // @[Bitwise.scala 50:65:@979.4]
  assign _T_3061 = _T_3056[4]; // @[Bitwise.scala 50:65:@980.4]
  assign _T_3062 = _T_3056[5]; // @[Bitwise.scala 50:65:@981.4]
  assign _T_3063 = _T_3056[6]; // @[Bitwise.scala 50:65:@982.4]
  assign _T_3064 = _T_3056[7]; // @[Bitwise.scala 50:65:@983.4]
  assign _T_3065 = _T_3056[8]; // @[Bitwise.scala 50:65:@984.4]
  assign _T_3066 = _T_3056[9]; // @[Bitwise.scala 50:65:@985.4]
  assign _T_3067 = _T_3056[10]; // @[Bitwise.scala 50:65:@986.4]
  assign _T_3068 = _T_3056[11]; // @[Bitwise.scala 50:65:@987.4]
  assign _T_3069 = _T_3058 + _T_3059; // @[Bitwise.scala 48:55:@988.4]
  assign _GEN_561 = {{1'd0}, _T_3057}; // @[Bitwise.scala 48:55:@989.4]
  assign _T_3070 = _GEN_561 + _T_3069; // @[Bitwise.scala 48:55:@989.4]
  assign _T_3071 = _T_3061 + _T_3062; // @[Bitwise.scala 48:55:@990.4]
  assign _GEN_562 = {{1'd0}, _T_3060}; // @[Bitwise.scala 48:55:@991.4]
  assign _T_3072 = _GEN_562 + _T_3071; // @[Bitwise.scala 48:55:@991.4]
  assign _T_3073 = _T_3070 + _T_3072; // @[Bitwise.scala 48:55:@992.4]
  assign _T_3074 = _T_3064 + _T_3065; // @[Bitwise.scala 48:55:@993.4]
  assign _GEN_563 = {{1'd0}, _T_3063}; // @[Bitwise.scala 48:55:@994.4]
  assign _T_3075 = _GEN_563 + _T_3074; // @[Bitwise.scala 48:55:@994.4]
  assign _T_3076 = _T_3067 + _T_3068; // @[Bitwise.scala 48:55:@995.4]
  assign _GEN_564 = {{1'd0}, _T_3066}; // @[Bitwise.scala 48:55:@996.4]
  assign _T_3077 = _GEN_564 + _T_3076; // @[Bitwise.scala 48:55:@996.4]
  assign _T_3078 = _T_3075 + _T_3077; // @[Bitwise.scala 48:55:@997.4]
  assign _T_3079 = _T_3073 + _T_3078; // @[Bitwise.scala 48:55:@998.4]
  assign _T_3143 = _T_2230[12:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1063.4]
  assign _T_3144 = _T_3143[0]; // @[Bitwise.scala 50:65:@1064.4]
  assign _T_3145 = _T_3143[1]; // @[Bitwise.scala 50:65:@1065.4]
  assign _T_3146 = _T_3143[2]; // @[Bitwise.scala 50:65:@1066.4]
  assign _T_3147 = _T_3143[3]; // @[Bitwise.scala 50:65:@1067.4]
  assign _T_3148 = _T_3143[4]; // @[Bitwise.scala 50:65:@1068.4]
  assign _T_3149 = _T_3143[5]; // @[Bitwise.scala 50:65:@1069.4]
  assign _T_3150 = _T_3143[6]; // @[Bitwise.scala 50:65:@1070.4]
  assign _T_3151 = _T_3143[7]; // @[Bitwise.scala 50:65:@1071.4]
  assign _T_3152 = _T_3143[8]; // @[Bitwise.scala 50:65:@1072.4]
  assign _T_3153 = _T_3143[9]; // @[Bitwise.scala 50:65:@1073.4]
  assign _T_3154 = _T_3143[10]; // @[Bitwise.scala 50:65:@1074.4]
  assign _T_3155 = _T_3143[11]; // @[Bitwise.scala 50:65:@1075.4]
  assign _T_3156 = _T_3143[12]; // @[Bitwise.scala 50:65:@1076.4]
  assign _T_3157 = _T_3145 + _T_3146; // @[Bitwise.scala 48:55:@1077.4]
  assign _GEN_565 = {{1'd0}, _T_3144}; // @[Bitwise.scala 48:55:@1078.4]
  assign _T_3158 = _GEN_565 + _T_3157; // @[Bitwise.scala 48:55:@1078.4]
  assign _T_3159 = _T_3148 + _T_3149; // @[Bitwise.scala 48:55:@1079.4]
  assign _GEN_566 = {{1'd0}, _T_3147}; // @[Bitwise.scala 48:55:@1080.4]
  assign _T_3160 = _GEN_566 + _T_3159; // @[Bitwise.scala 48:55:@1080.4]
  assign _T_3161 = _T_3158 + _T_3160; // @[Bitwise.scala 48:55:@1081.4]
  assign _T_3162 = _T_3151 + _T_3152; // @[Bitwise.scala 48:55:@1082.4]
  assign _GEN_567 = {{1'd0}, _T_3150}; // @[Bitwise.scala 48:55:@1083.4]
  assign _T_3163 = _GEN_567 + _T_3162; // @[Bitwise.scala 48:55:@1083.4]
  assign _T_3164 = _T_3153 + _T_3154; // @[Bitwise.scala 48:55:@1084.4]
  assign _T_3165 = _T_3155 + _T_3156; // @[Bitwise.scala 48:55:@1085.4]
  assign _T_3166 = _T_3164 + _T_3165; // @[Bitwise.scala 48:55:@1086.4]
  assign _T_3167 = _T_3163 + _T_3166; // @[Bitwise.scala 48:55:@1087.4]
  assign _T_3168 = _T_3161 + _T_3167; // @[Bitwise.scala 48:55:@1088.4]
  assign _T_3232 = _T_2230[13:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1153.4]
  assign _T_3233 = _T_3232[0]; // @[Bitwise.scala 50:65:@1154.4]
  assign _T_3234 = _T_3232[1]; // @[Bitwise.scala 50:65:@1155.4]
  assign _T_3235 = _T_3232[2]; // @[Bitwise.scala 50:65:@1156.4]
  assign _T_3236 = _T_3232[3]; // @[Bitwise.scala 50:65:@1157.4]
  assign _T_3237 = _T_3232[4]; // @[Bitwise.scala 50:65:@1158.4]
  assign _T_3238 = _T_3232[5]; // @[Bitwise.scala 50:65:@1159.4]
  assign _T_3239 = _T_3232[6]; // @[Bitwise.scala 50:65:@1160.4]
  assign _T_3240 = _T_3232[7]; // @[Bitwise.scala 50:65:@1161.4]
  assign _T_3241 = _T_3232[8]; // @[Bitwise.scala 50:65:@1162.4]
  assign _T_3242 = _T_3232[9]; // @[Bitwise.scala 50:65:@1163.4]
  assign _T_3243 = _T_3232[10]; // @[Bitwise.scala 50:65:@1164.4]
  assign _T_3244 = _T_3232[11]; // @[Bitwise.scala 50:65:@1165.4]
  assign _T_3245 = _T_3232[12]; // @[Bitwise.scala 50:65:@1166.4]
  assign _T_3246 = _T_3232[13]; // @[Bitwise.scala 50:65:@1167.4]
  assign _T_3247 = _T_3234 + _T_3235; // @[Bitwise.scala 48:55:@1168.4]
  assign _GEN_568 = {{1'd0}, _T_3233}; // @[Bitwise.scala 48:55:@1169.4]
  assign _T_3248 = _GEN_568 + _T_3247; // @[Bitwise.scala 48:55:@1169.4]
  assign _T_3249 = _T_3236 + _T_3237; // @[Bitwise.scala 48:55:@1170.4]
  assign _T_3250 = _T_3238 + _T_3239; // @[Bitwise.scala 48:55:@1171.4]
  assign _T_3251 = _T_3249 + _T_3250; // @[Bitwise.scala 48:55:@1172.4]
  assign _T_3252 = _T_3248 + _T_3251; // @[Bitwise.scala 48:55:@1173.4]
  assign _T_3253 = _T_3241 + _T_3242; // @[Bitwise.scala 48:55:@1174.4]
  assign _GEN_569 = {{1'd0}, _T_3240}; // @[Bitwise.scala 48:55:@1175.4]
  assign _T_3254 = _GEN_569 + _T_3253; // @[Bitwise.scala 48:55:@1175.4]
  assign _T_3255 = _T_3243 + _T_3244; // @[Bitwise.scala 48:55:@1176.4]
  assign _T_3256 = _T_3245 + _T_3246; // @[Bitwise.scala 48:55:@1177.4]
  assign _T_3257 = _T_3255 + _T_3256; // @[Bitwise.scala 48:55:@1178.4]
  assign _T_3258 = _T_3254 + _T_3257; // @[Bitwise.scala 48:55:@1179.4]
  assign _T_3259 = _T_3252 + _T_3258; // @[Bitwise.scala 48:55:@1180.4]
  assign _T_3323 = _T_2230[14:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1245.4]
  assign _T_3324 = _T_3323[0]; // @[Bitwise.scala 50:65:@1246.4]
  assign _T_3325 = _T_3323[1]; // @[Bitwise.scala 50:65:@1247.4]
  assign _T_3326 = _T_3323[2]; // @[Bitwise.scala 50:65:@1248.4]
  assign _T_3327 = _T_3323[3]; // @[Bitwise.scala 50:65:@1249.4]
  assign _T_3328 = _T_3323[4]; // @[Bitwise.scala 50:65:@1250.4]
  assign _T_3329 = _T_3323[5]; // @[Bitwise.scala 50:65:@1251.4]
  assign _T_3330 = _T_3323[6]; // @[Bitwise.scala 50:65:@1252.4]
  assign _T_3331 = _T_3323[7]; // @[Bitwise.scala 50:65:@1253.4]
  assign _T_3332 = _T_3323[8]; // @[Bitwise.scala 50:65:@1254.4]
  assign _T_3333 = _T_3323[9]; // @[Bitwise.scala 50:65:@1255.4]
  assign _T_3334 = _T_3323[10]; // @[Bitwise.scala 50:65:@1256.4]
  assign _T_3335 = _T_3323[11]; // @[Bitwise.scala 50:65:@1257.4]
  assign _T_3336 = _T_3323[12]; // @[Bitwise.scala 50:65:@1258.4]
  assign _T_3337 = _T_3323[13]; // @[Bitwise.scala 50:65:@1259.4]
  assign _T_3338 = _T_3323[14]; // @[Bitwise.scala 50:65:@1260.4]
  assign _T_3339 = _T_3325 + _T_3326; // @[Bitwise.scala 48:55:@1261.4]
  assign _GEN_570 = {{1'd0}, _T_3324}; // @[Bitwise.scala 48:55:@1262.4]
  assign _T_3340 = _GEN_570 + _T_3339; // @[Bitwise.scala 48:55:@1262.4]
  assign _T_3341 = _T_3327 + _T_3328; // @[Bitwise.scala 48:55:@1263.4]
  assign _T_3342 = _T_3329 + _T_3330; // @[Bitwise.scala 48:55:@1264.4]
  assign _T_3343 = _T_3341 + _T_3342; // @[Bitwise.scala 48:55:@1265.4]
  assign _T_3344 = _T_3340 + _T_3343; // @[Bitwise.scala 48:55:@1266.4]
  assign _T_3345 = _T_3331 + _T_3332; // @[Bitwise.scala 48:55:@1267.4]
  assign _T_3346 = _T_3333 + _T_3334; // @[Bitwise.scala 48:55:@1268.4]
  assign _T_3347 = _T_3345 + _T_3346; // @[Bitwise.scala 48:55:@1269.4]
  assign _T_3348 = _T_3335 + _T_3336; // @[Bitwise.scala 48:55:@1270.4]
  assign _T_3349 = _T_3337 + _T_3338; // @[Bitwise.scala 48:55:@1271.4]
  assign _T_3350 = _T_3348 + _T_3349; // @[Bitwise.scala 48:55:@1272.4]
  assign _T_3351 = _T_3347 + _T_3350; // @[Bitwise.scala 48:55:@1273.4]
  assign _T_3352 = _T_3344 + _T_3351; // @[Bitwise.scala 48:55:@1274.4]
  assign _T_3416 = _T_2230[15:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1339.4]
  assign _T_3417 = _T_3416[0]; // @[Bitwise.scala 50:65:@1340.4]
  assign _T_3418 = _T_3416[1]; // @[Bitwise.scala 50:65:@1341.4]
  assign _T_3419 = _T_3416[2]; // @[Bitwise.scala 50:65:@1342.4]
  assign _T_3420 = _T_3416[3]; // @[Bitwise.scala 50:65:@1343.4]
  assign _T_3421 = _T_3416[4]; // @[Bitwise.scala 50:65:@1344.4]
  assign _T_3422 = _T_3416[5]; // @[Bitwise.scala 50:65:@1345.4]
  assign _T_3423 = _T_3416[6]; // @[Bitwise.scala 50:65:@1346.4]
  assign _T_3424 = _T_3416[7]; // @[Bitwise.scala 50:65:@1347.4]
  assign _T_3425 = _T_3416[8]; // @[Bitwise.scala 50:65:@1348.4]
  assign _T_3426 = _T_3416[9]; // @[Bitwise.scala 50:65:@1349.4]
  assign _T_3427 = _T_3416[10]; // @[Bitwise.scala 50:65:@1350.4]
  assign _T_3428 = _T_3416[11]; // @[Bitwise.scala 50:65:@1351.4]
  assign _T_3429 = _T_3416[12]; // @[Bitwise.scala 50:65:@1352.4]
  assign _T_3430 = _T_3416[13]; // @[Bitwise.scala 50:65:@1353.4]
  assign _T_3431 = _T_3416[14]; // @[Bitwise.scala 50:65:@1354.4]
  assign _T_3432 = _T_3416[15]; // @[Bitwise.scala 50:65:@1355.4]
  assign _T_3433 = _T_3417 + _T_3418; // @[Bitwise.scala 48:55:@1356.4]
  assign _T_3434 = _T_3419 + _T_3420; // @[Bitwise.scala 48:55:@1357.4]
  assign _T_3435 = _T_3433 + _T_3434; // @[Bitwise.scala 48:55:@1358.4]
  assign _T_3436 = _T_3421 + _T_3422; // @[Bitwise.scala 48:55:@1359.4]
  assign _T_3437 = _T_3423 + _T_3424; // @[Bitwise.scala 48:55:@1360.4]
  assign _T_3438 = _T_3436 + _T_3437; // @[Bitwise.scala 48:55:@1361.4]
  assign _T_3439 = _T_3435 + _T_3438; // @[Bitwise.scala 48:55:@1362.4]
  assign _T_3440 = _T_3425 + _T_3426; // @[Bitwise.scala 48:55:@1363.4]
  assign _T_3441 = _T_3427 + _T_3428; // @[Bitwise.scala 48:55:@1364.4]
  assign _T_3442 = _T_3440 + _T_3441; // @[Bitwise.scala 48:55:@1365.4]
  assign _T_3443 = _T_3429 + _T_3430; // @[Bitwise.scala 48:55:@1366.4]
  assign _T_3444 = _T_3431 + _T_3432; // @[Bitwise.scala 48:55:@1367.4]
  assign _T_3445 = _T_3443 + _T_3444; // @[Bitwise.scala 48:55:@1368.4]
  assign _T_3446 = _T_3442 + _T_3445; // @[Bitwise.scala 48:55:@1369.4]
  assign _T_3447 = _T_3439 + _T_3446; // @[Bitwise.scala 48:55:@1370.4]
  assign _T_3511 = _T_2230[16:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1435.4]
  assign _T_3512 = _T_3511[0]; // @[Bitwise.scala 50:65:@1436.4]
  assign _T_3513 = _T_3511[1]; // @[Bitwise.scala 50:65:@1437.4]
  assign _T_3514 = _T_3511[2]; // @[Bitwise.scala 50:65:@1438.4]
  assign _T_3515 = _T_3511[3]; // @[Bitwise.scala 50:65:@1439.4]
  assign _T_3516 = _T_3511[4]; // @[Bitwise.scala 50:65:@1440.4]
  assign _T_3517 = _T_3511[5]; // @[Bitwise.scala 50:65:@1441.4]
  assign _T_3518 = _T_3511[6]; // @[Bitwise.scala 50:65:@1442.4]
  assign _T_3519 = _T_3511[7]; // @[Bitwise.scala 50:65:@1443.4]
  assign _T_3520 = _T_3511[8]; // @[Bitwise.scala 50:65:@1444.4]
  assign _T_3521 = _T_3511[9]; // @[Bitwise.scala 50:65:@1445.4]
  assign _T_3522 = _T_3511[10]; // @[Bitwise.scala 50:65:@1446.4]
  assign _T_3523 = _T_3511[11]; // @[Bitwise.scala 50:65:@1447.4]
  assign _T_3524 = _T_3511[12]; // @[Bitwise.scala 50:65:@1448.4]
  assign _T_3525 = _T_3511[13]; // @[Bitwise.scala 50:65:@1449.4]
  assign _T_3526 = _T_3511[14]; // @[Bitwise.scala 50:65:@1450.4]
  assign _T_3527 = _T_3511[15]; // @[Bitwise.scala 50:65:@1451.4]
  assign _T_3528 = _T_3511[16]; // @[Bitwise.scala 50:65:@1452.4]
  assign _T_3529 = _T_3512 + _T_3513; // @[Bitwise.scala 48:55:@1453.4]
  assign _T_3530 = _T_3514 + _T_3515; // @[Bitwise.scala 48:55:@1454.4]
  assign _T_3531 = _T_3529 + _T_3530; // @[Bitwise.scala 48:55:@1455.4]
  assign _T_3532 = _T_3516 + _T_3517; // @[Bitwise.scala 48:55:@1456.4]
  assign _T_3533 = _T_3518 + _T_3519; // @[Bitwise.scala 48:55:@1457.4]
  assign _T_3534 = _T_3532 + _T_3533; // @[Bitwise.scala 48:55:@1458.4]
  assign _T_3535 = _T_3531 + _T_3534; // @[Bitwise.scala 48:55:@1459.4]
  assign _T_3536 = _T_3520 + _T_3521; // @[Bitwise.scala 48:55:@1460.4]
  assign _T_3537 = _T_3522 + _T_3523; // @[Bitwise.scala 48:55:@1461.4]
  assign _T_3538 = _T_3536 + _T_3537; // @[Bitwise.scala 48:55:@1462.4]
  assign _T_3539 = _T_3524 + _T_3525; // @[Bitwise.scala 48:55:@1463.4]
  assign _T_3540 = _T_3527 + _T_3528; // @[Bitwise.scala 48:55:@1464.4]
  assign _GEN_571 = {{1'd0}, _T_3526}; // @[Bitwise.scala 48:55:@1465.4]
  assign _T_3541 = _GEN_571 + _T_3540; // @[Bitwise.scala 48:55:@1465.4]
  assign _GEN_572 = {{1'd0}, _T_3539}; // @[Bitwise.scala 48:55:@1466.4]
  assign _T_3542 = _GEN_572 + _T_3541; // @[Bitwise.scala 48:55:@1466.4]
  assign _GEN_573 = {{1'd0}, _T_3538}; // @[Bitwise.scala 48:55:@1467.4]
  assign _T_3543 = _GEN_573 + _T_3542; // @[Bitwise.scala 48:55:@1467.4]
  assign _GEN_574 = {{1'd0}, _T_3535}; // @[Bitwise.scala 48:55:@1468.4]
  assign _T_3544 = _GEN_574 + _T_3543; // @[Bitwise.scala 48:55:@1468.4]
  assign _T_3608 = _T_2230[17:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1533.4]
  assign _T_3609 = _T_3608[0]; // @[Bitwise.scala 50:65:@1534.4]
  assign _T_3610 = _T_3608[1]; // @[Bitwise.scala 50:65:@1535.4]
  assign _T_3611 = _T_3608[2]; // @[Bitwise.scala 50:65:@1536.4]
  assign _T_3612 = _T_3608[3]; // @[Bitwise.scala 50:65:@1537.4]
  assign _T_3613 = _T_3608[4]; // @[Bitwise.scala 50:65:@1538.4]
  assign _T_3614 = _T_3608[5]; // @[Bitwise.scala 50:65:@1539.4]
  assign _T_3615 = _T_3608[6]; // @[Bitwise.scala 50:65:@1540.4]
  assign _T_3616 = _T_3608[7]; // @[Bitwise.scala 50:65:@1541.4]
  assign _T_3617 = _T_3608[8]; // @[Bitwise.scala 50:65:@1542.4]
  assign _T_3618 = _T_3608[9]; // @[Bitwise.scala 50:65:@1543.4]
  assign _T_3619 = _T_3608[10]; // @[Bitwise.scala 50:65:@1544.4]
  assign _T_3620 = _T_3608[11]; // @[Bitwise.scala 50:65:@1545.4]
  assign _T_3621 = _T_3608[12]; // @[Bitwise.scala 50:65:@1546.4]
  assign _T_3622 = _T_3608[13]; // @[Bitwise.scala 50:65:@1547.4]
  assign _T_3623 = _T_3608[14]; // @[Bitwise.scala 50:65:@1548.4]
  assign _T_3624 = _T_3608[15]; // @[Bitwise.scala 50:65:@1549.4]
  assign _T_3625 = _T_3608[16]; // @[Bitwise.scala 50:65:@1550.4]
  assign _T_3626 = _T_3608[17]; // @[Bitwise.scala 50:65:@1551.4]
  assign _T_3627 = _T_3609 + _T_3610; // @[Bitwise.scala 48:55:@1552.4]
  assign _T_3628 = _T_3611 + _T_3612; // @[Bitwise.scala 48:55:@1553.4]
  assign _T_3629 = _T_3627 + _T_3628; // @[Bitwise.scala 48:55:@1554.4]
  assign _T_3630 = _T_3613 + _T_3614; // @[Bitwise.scala 48:55:@1555.4]
  assign _T_3631 = _T_3616 + _T_3617; // @[Bitwise.scala 48:55:@1556.4]
  assign _GEN_575 = {{1'd0}, _T_3615}; // @[Bitwise.scala 48:55:@1557.4]
  assign _T_3632 = _GEN_575 + _T_3631; // @[Bitwise.scala 48:55:@1557.4]
  assign _GEN_576 = {{1'd0}, _T_3630}; // @[Bitwise.scala 48:55:@1558.4]
  assign _T_3633 = _GEN_576 + _T_3632; // @[Bitwise.scala 48:55:@1558.4]
  assign _GEN_577 = {{1'd0}, _T_3629}; // @[Bitwise.scala 48:55:@1559.4]
  assign _T_3634 = _GEN_577 + _T_3633; // @[Bitwise.scala 48:55:@1559.4]
  assign _T_3635 = _T_3618 + _T_3619; // @[Bitwise.scala 48:55:@1560.4]
  assign _T_3636 = _T_3620 + _T_3621; // @[Bitwise.scala 48:55:@1561.4]
  assign _T_3637 = _T_3635 + _T_3636; // @[Bitwise.scala 48:55:@1562.4]
  assign _T_3638 = _T_3622 + _T_3623; // @[Bitwise.scala 48:55:@1563.4]
  assign _T_3639 = _T_3625 + _T_3626; // @[Bitwise.scala 48:55:@1564.4]
  assign _GEN_578 = {{1'd0}, _T_3624}; // @[Bitwise.scala 48:55:@1565.4]
  assign _T_3640 = _GEN_578 + _T_3639; // @[Bitwise.scala 48:55:@1565.4]
  assign _GEN_579 = {{1'd0}, _T_3638}; // @[Bitwise.scala 48:55:@1566.4]
  assign _T_3641 = _GEN_579 + _T_3640; // @[Bitwise.scala 48:55:@1566.4]
  assign _GEN_580 = {{1'd0}, _T_3637}; // @[Bitwise.scala 48:55:@1567.4]
  assign _T_3642 = _GEN_580 + _T_3641; // @[Bitwise.scala 48:55:@1567.4]
  assign _T_3643 = _T_3634 + _T_3642; // @[Bitwise.scala 48:55:@1568.4]
  assign _T_3707 = _T_2230[18:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1633.4]
  assign _T_3708 = _T_3707[0]; // @[Bitwise.scala 50:65:@1634.4]
  assign _T_3709 = _T_3707[1]; // @[Bitwise.scala 50:65:@1635.4]
  assign _T_3710 = _T_3707[2]; // @[Bitwise.scala 50:65:@1636.4]
  assign _T_3711 = _T_3707[3]; // @[Bitwise.scala 50:65:@1637.4]
  assign _T_3712 = _T_3707[4]; // @[Bitwise.scala 50:65:@1638.4]
  assign _T_3713 = _T_3707[5]; // @[Bitwise.scala 50:65:@1639.4]
  assign _T_3714 = _T_3707[6]; // @[Bitwise.scala 50:65:@1640.4]
  assign _T_3715 = _T_3707[7]; // @[Bitwise.scala 50:65:@1641.4]
  assign _T_3716 = _T_3707[8]; // @[Bitwise.scala 50:65:@1642.4]
  assign _T_3717 = _T_3707[9]; // @[Bitwise.scala 50:65:@1643.4]
  assign _T_3718 = _T_3707[10]; // @[Bitwise.scala 50:65:@1644.4]
  assign _T_3719 = _T_3707[11]; // @[Bitwise.scala 50:65:@1645.4]
  assign _T_3720 = _T_3707[12]; // @[Bitwise.scala 50:65:@1646.4]
  assign _T_3721 = _T_3707[13]; // @[Bitwise.scala 50:65:@1647.4]
  assign _T_3722 = _T_3707[14]; // @[Bitwise.scala 50:65:@1648.4]
  assign _T_3723 = _T_3707[15]; // @[Bitwise.scala 50:65:@1649.4]
  assign _T_3724 = _T_3707[16]; // @[Bitwise.scala 50:65:@1650.4]
  assign _T_3725 = _T_3707[17]; // @[Bitwise.scala 50:65:@1651.4]
  assign _T_3726 = _T_3707[18]; // @[Bitwise.scala 50:65:@1652.4]
  assign _T_3727 = _T_3708 + _T_3709; // @[Bitwise.scala 48:55:@1653.4]
  assign _T_3728 = _T_3710 + _T_3711; // @[Bitwise.scala 48:55:@1654.4]
  assign _T_3729 = _T_3727 + _T_3728; // @[Bitwise.scala 48:55:@1655.4]
  assign _T_3730 = _T_3712 + _T_3713; // @[Bitwise.scala 48:55:@1656.4]
  assign _T_3731 = _T_3715 + _T_3716; // @[Bitwise.scala 48:55:@1657.4]
  assign _GEN_581 = {{1'd0}, _T_3714}; // @[Bitwise.scala 48:55:@1658.4]
  assign _T_3732 = _GEN_581 + _T_3731; // @[Bitwise.scala 48:55:@1658.4]
  assign _GEN_582 = {{1'd0}, _T_3730}; // @[Bitwise.scala 48:55:@1659.4]
  assign _T_3733 = _GEN_582 + _T_3732; // @[Bitwise.scala 48:55:@1659.4]
  assign _GEN_583 = {{1'd0}, _T_3729}; // @[Bitwise.scala 48:55:@1660.4]
  assign _T_3734 = _GEN_583 + _T_3733; // @[Bitwise.scala 48:55:@1660.4]
  assign _T_3735 = _T_3717 + _T_3718; // @[Bitwise.scala 48:55:@1661.4]
  assign _T_3736 = _T_3720 + _T_3721; // @[Bitwise.scala 48:55:@1662.4]
  assign _GEN_584 = {{1'd0}, _T_3719}; // @[Bitwise.scala 48:55:@1663.4]
  assign _T_3737 = _GEN_584 + _T_3736; // @[Bitwise.scala 48:55:@1663.4]
  assign _GEN_585 = {{1'd0}, _T_3735}; // @[Bitwise.scala 48:55:@1664.4]
  assign _T_3738 = _GEN_585 + _T_3737; // @[Bitwise.scala 48:55:@1664.4]
  assign _T_3739 = _T_3722 + _T_3723; // @[Bitwise.scala 48:55:@1665.4]
  assign _T_3740 = _T_3725 + _T_3726; // @[Bitwise.scala 48:55:@1666.4]
  assign _GEN_586 = {{1'd0}, _T_3724}; // @[Bitwise.scala 48:55:@1667.4]
  assign _T_3741 = _GEN_586 + _T_3740; // @[Bitwise.scala 48:55:@1667.4]
  assign _GEN_587 = {{1'd0}, _T_3739}; // @[Bitwise.scala 48:55:@1668.4]
  assign _T_3742 = _GEN_587 + _T_3741; // @[Bitwise.scala 48:55:@1668.4]
  assign _T_3743 = _T_3738 + _T_3742; // @[Bitwise.scala 48:55:@1669.4]
  assign _T_3744 = _T_3734 + _T_3743; // @[Bitwise.scala 48:55:@1670.4]
  assign _T_3808 = _T_2230[19:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1735.4]
  assign _T_3809 = _T_3808[0]; // @[Bitwise.scala 50:65:@1736.4]
  assign _T_3810 = _T_3808[1]; // @[Bitwise.scala 50:65:@1737.4]
  assign _T_3811 = _T_3808[2]; // @[Bitwise.scala 50:65:@1738.4]
  assign _T_3812 = _T_3808[3]; // @[Bitwise.scala 50:65:@1739.4]
  assign _T_3813 = _T_3808[4]; // @[Bitwise.scala 50:65:@1740.4]
  assign _T_3814 = _T_3808[5]; // @[Bitwise.scala 50:65:@1741.4]
  assign _T_3815 = _T_3808[6]; // @[Bitwise.scala 50:65:@1742.4]
  assign _T_3816 = _T_3808[7]; // @[Bitwise.scala 50:65:@1743.4]
  assign _T_3817 = _T_3808[8]; // @[Bitwise.scala 50:65:@1744.4]
  assign _T_3818 = _T_3808[9]; // @[Bitwise.scala 50:65:@1745.4]
  assign _T_3819 = _T_3808[10]; // @[Bitwise.scala 50:65:@1746.4]
  assign _T_3820 = _T_3808[11]; // @[Bitwise.scala 50:65:@1747.4]
  assign _T_3821 = _T_3808[12]; // @[Bitwise.scala 50:65:@1748.4]
  assign _T_3822 = _T_3808[13]; // @[Bitwise.scala 50:65:@1749.4]
  assign _T_3823 = _T_3808[14]; // @[Bitwise.scala 50:65:@1750.4]
  assign _T_3824 = _T_3808[15]; // @[Bitwise.scala 50:65:@1751.4]
  assign _T_3825 = _T_3808[16]; // @[Bitwise.scala 50:65:@1752.4]
  assign _T_3826 = _T_3808[17]; // @[Bitwise.scala 50:65:@1753.4]
  assign _T_3827 = _T_3808[18]; // @[Bitwise.scala 50:65:@1754.4]
  assign _T_3828 = _T_3808[19]; // @[Bitwise.scala 50:65:@1755.4]
  assign _T_3829 = _T_3809 + _T_3810; // @[Bitwise.scala 48:55:@1756.4]
  assign _T_3830 = _T_3812 + _T_3813; // @[Bitwise.scala 48:55:@1757.4]
  assign _GEN_588 = {{1'd0}, _T_3811}; // @[Bitwise.scala 48:55:@1758.4]
  assign _T_3831 = _GEN_588 + _T_3830; // @[Bitwise.scala 48:55:@1758.4]
  assign _GEN_589 = {{1'd0}, _T_3829}; // @[Bitwise.scala 48:55:@1759.4]
  assign _T_3832 = _GEN_589 + _T_3831; // @[Bitwise.scala 48:55:@1759.4]
  assign _T_3833 = _T_3814 + _T_3815; // @[Bitwise.scala 48:55:@1760.4]
  assign _T_3834 = _T_3817 + _T_3818; // @[Bitwise.scala 48:55:@1761.4]
  assign _GEN_590 = {{1'd0}, _T_3816}; // @[Bitwise.scala 48:55:@1762.4]
  assign _T_3835 = _GEN_590 + _T_3834; // @[Bitwise.scala 48:55:@1762.4]
  assign _GEN_591 = {{1'd0}, _T_3833}; // @[Bitwise.scala 48:55:@1763.4]
  assign _T_3836 = _GEN_591 + _T_3835; // @[Bitwise.scala 48:55:@1763.4]
  assign _T_3837 = _T_3832 + _T_3836; // @[Bitwise.scala 48:55:@1764.4]
  assign _T_3838 = _T_3819 + _T_3820; // @[Bitwise.scala 48:55:@1765.4]
  assign _T_3839 = _T_3822 + _T_3823; // @[Bitwise.scala 48:55:@1766.4]
  assign _GEN_592 = {{1'd0}, _T_3821}; // @[Bitwise.scala 48:55:@1767.4]
  assign _T_3840 = _GEN_592 + _T_3839; // @[Bitwise.scala 48:55:@1767.4]
  assign _GEN_593 = {{1'd0}, _T_3838}; // @[Bitwise.scala 48:55:@1768.4]
  assign _T_3841 = _GEN_593 + _T_3840; // @[Bitwise.scala 48:55:@1768.4]
  assign _T_3842 = _T_3824 + _T_3825; // @[Bitwise.scala 48:55:@1769.4]
  assign _T_3843 = _T_3827 + _T_3828; // @[Bitwise.scala 48:55:@1770.4]
  assign _GEN_594 = {{1'd0}, _T_3826}; // @[Bitwise.scala 48:55:@1771.4]
  assign _T_3844 = _GEN_594 + _T_3843; // @[Bitwise.scala 48:55:@1771.4]
  assign _GEN_595 = {{1'd0}, _T_3842}; // @[Bitwise.scala 48:55:@1772.4]
  assign _T_3845 = _GEN_595 + _T_3844; // @[Bitwise.scala 48:55:@1772.4]
  assign _T_3846 = _T_3841 + _T_3845; // @[Bitwise.scala 48:55:@1773.4]
  assign _T_3847 = _T_3837 + _T_3846; // @[Bitwise.scala 48:55:@1774.4]
  assign _T_3911 = _T_2230[20:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1839.4]
  assign _T_3912 = _T_3911[0]; // @[Bitwise.scala 50:65:@1840.4]
  assign _T_3913 = _T_3911[1]; // @[Bitwise.scala 50:65:@1841.4]
  assign _T_3914 = _T_3911[2]; // @[Bitwise.scala 50:65:@1842.4]
  assign _T_3915 = _T_3911[3]; // @[Bitwise.scala 50:65:@1843.4]
  assign _T_3916 = _T_3911[4]; // @[Bitwise.scala 50:65:@1844.4]
  assign _T_3917 = _T_3911[5]; // @[Bitwise.scala 50:65:@1845.4]
  assign _T_3918 = _T_3911[6]; // @[Bitwise.scala 50:65:@1846.4]
  assign _T_3919 = _T_3911[7]; // @[Bitwise.scala 50:65:@1847.4]
  assign _T_3920 = _T_3911[8]; // @[Bitwise.scala 50:65:@1848.4]
  assign _T_3921 = _T_3911[9]; // @[Bitwise.scala 50:65:@1849.4]
  assign _T_3922 = _T_3911[10]; // @[Bitwise.scala 50:65:@1850.4]
  assign _T_3923 = _T_3911[11]; // @[Bitwise.scala 50:65:@1851.4]
  assign _T_3924 = _T_3911[12]; // @[Bitwise.scala 50:65:@1852.4]
  assign _T_3925 = _T_3911[13]; // @[Bitwise.scala 50:65:@1853.4]
  assign _T_3926 = _T_3911[14]; // @[Bitwise.scala 50:65:@1854.4]
  assign _T_3927 = _T_3911[15]; // @[Bitwise.scala 50:65:@1855.4]
  assign _T_3928 = _T_3911[16]; // @[Bitwise.scala 50:65:@1856.4]
  assign _T_3929 = _T_3911[17]; // @[Bitwise.scala 50:65:@1857.4]
  assign _T_3930 = _T_3911[18]; // @[Bitwise.scala 50:65:@1858.4]
  assign _T_3931 = _T_3911[19]; // @[Bitwise.scala 50:65:@1859.4]
  assign _T_3932 = _T_3911[20]; // @[Bitwise.scala 50:65:@1860.4]
  assign _T_3933 = _T_3912 + _T_3913; // @[Bitwise.scala 48:55:@1861.4]
  assign _T_3934 = _T_3915 + _T_3916; // @[Bitwise.scala 48:55:@1862.4]
  assign _GEN_596 = {{1'd0}, _T_3914}; // @[Bitwise.scala 48:55:@1863.4]
  assign _T_3935 = _GEN_596 + _T_3934; // @[Bitwise.scala 48:55:@1863.4]
  assign _GEN_597 = {{1'd0}, _T_3933}; // @[Bitwise.scala 48:55:@1864.4]
  assign _T_3936 = _GEN_597 + _T_3935; // @[Bitwise.scala 48:55:@1864.4]
  assign _T_3937 = _T_3917 + _T_3918; // @[Bitwise.scala 48:55:@1865.4]
  assign _T_3938 = _T_3920 + _T_3921; // @[Bitwise.scala 48:55:@1866.4]
  assign _GEN_598 = {{1'd0}, _T_3919}; // @[Bitwise.scala 48:55:@1867.4]
  assign _T_3939 = _GEN_598 + _T_3938; // @[Bitwise.scala 48:55:@1867.4]
  assign _GEN_599 = {{1'd0}, _T_3937}; // @[Bitwise.scala 48:55:@1868.4]
  assign _T_3940 = _GEN_599 + _T_3939; // @[Bitwise.scala 48:55:@1868.4]
  assign _T_3941 = _T_3936 + _T_3940; // @[Bitwise.scala 48:55:@1869.4]
  assign _T_3942 = _T_3922 + _T_3923; // @[Bitwise.scala 48:55:@1870.4]
  assign _T_3943 = _T_3925 + _T_3926; // @[Bitwise.scala 48:55:@1871.4]
  assign _GEN_600 = {{1'd0}, _T_3924}; // @[Bitwise.scala 48:55:@1872.4]
  assign _T_3944 = _GEN_600 + _T_3943; // @[Bitwise.scala 48:55:@1872.4]
  assign _GEN_601 = {{1'd0}, _T_3942}; // @[Bitwise.scala 48:55:@1873.4]
  assign _T_3945 = _GEN_601 + _T_3944; // @[Bitwise.scala 48:55:@1873.4]
  assign _T_3946 = _T_3928 + _T_3929; // @[Bitwise.scala 48:55:@1874.4]
  assign _GEN_602 = {{1'd0}, _T_3927}; // @[Bitwise.scala 48:55:@1875.4]
  assign _T_3947 = _GEN_602 + _T_3946; // @[Bitwise.scala 48:55:@1875.4]
  assign _T_3948 = _T_3931 + _T_3932; // @[Bitwise.scala 48:55:@1876.4]
  assign _GEN_603 = {{1'd0}, _T_3930}; // @[Bitwise.scala 48:55:@1877.4]
  assign _T_3949 = _GEN_603 + _T_3948; // @[Bitwise.scala 48:55:@1877.4]
  assign _T_3950 = _T_3947 + _T_3949; // @[Bitwise.scala 48:55:@1878.4]
  assign _T_3951 = _T_3945 + _T_3950; // @[Bitwise.scala 48:55:@1879.4]
  assign _T_3952 = _T_3941 + _T_3951; // @[Bitwise.scala 48:55:@1880.4]
  assign _T_4016 = _T_2230[21:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@1945.4]
  assign _T_4017 = _T_4016[0]; // @[Bitwise.scala 50:65:@1946.4]
  assign _T_4018 = _T_4016[1]; // @[Bitwise.scala 50:65:@1947.4]
  assign _T_4019 = _T_4016[2]; // @[Bitwise.scala 50:65:@1948.4]
  assign _T_4020 = _T_4016[3]; // @[Bitwise.scala 50:65:@1949.4]
  assign _T_4021 = _T_4016[4]; // @[Bitwise.scala 50:65:@1950.4]
  assign _T_4022 = _T_4016[5]; // @[Bitwise.scala 50:65:@1951.4]
  assign _T_4023 = _T_4016[6]; // @[Bitwise.scala 50:65:@1952.4]
  assign _T_4024 = _T_4016[7]; // @[Bitwise.scala 50:65:@1953.4]
  assign _T_4025 = _T_4016[8]; // @[Bitwise.scala 50:65:@1954.4]
  assign _T_4026 = _T_4016[9]; // @[Bitwise.scala 50:65:@1955.4]
  assign _T_4027 = _T_4016[10]; // @[Bitwise.scala 50:65:@1956.4]
  assign _T_4028 = _T_4016[11]; // @[Bitwise.scala 50:65:@1957.4]
  assign _T_4029 = _T_4016[12]; // @[Bitwise.scala 50:65:@1958.4]
  assign _T_4030 = _T_4016[13]; // @[Bitwise.scala 50:65:@1959.4]
  assign _T_4031 = _T_4016[14]; // @[Bitwise.scala 50:65:@1960.4]
  assign _T_4032 = _T_4016[15]; // @[Bitwise.scala 50:65:@1961.4]
  assign _T_4033 = _T_4016[16]; // @[Bitwise.scala 50:65:@1962.4]
  assign _T_4034 = _T_4016[17]; // @[Bitwise.scala 50:65:@1963.4]
  assign _T_4035 = _T_4016[18]; // @[Bitwise.scala 50:65:@1964.4]
  assign _T_4036 = _T_4016[19]; // @[Bitwise.scala 50:65:@1965.4]
  assign _T_4037 = _T_4016[20]; // @[Bitwise.scala 50:65:@1966.4]
  assign _T_4038 = _T_4016[21]; // @[Bitwise.scala 50:65:@1967.4]
  assign _T_4039 = _T_4017 + _T_4018; // @[Bitwise.scala 48:55:@1968.4]
  assign _T_4040 = _T_4020 + _T_4021; // @[Bitwise.scala 48:55:@1969.4]
  assign _GEN_604 = {{1'd0}, _T_4019}; // @[Bitwise.scala 48:55:@1970.4]
  assign _T_4041 = _GEN_604 + _T_4040; // @[Bitwise.scala 48:55:@1970.4]
  assign _GEN_605 = {{1'd0}, _T_4039}; // @[Bitwise.scala 48:55:@1971.4]
  assign _T_4042 = _GEN_605 + _T_4041; // @[Bitwise.scala 48:55:@1971.4]
  assign _T_4043 = _T_4023 + _T_4024; // @[Bitwise.scala 48:55:@1972.4]
  assign _GEN_606 = {{1'd0}, _T_4022}; // @[Bitwise.scala 48:55:@1973.4]
  assign _T_4044 = _GEN_606 + _T_4043; // @[Bitwise.scala 48:55:@1973.4]
  assign _T_4045 = _T_4026 + _T_4027; // @[Bitwise.scala 48:55:@1974.4]
  assign _GEN_607 = {{1'd0}, _T_4025}; // @[Bitwise.scala 48:55:@1975.4]
  assign _T_4046 = _GEN_607 + _T_4045; // @[Bitwise.scala 48:55:@1975.4]
  assign _T_4047 = _T_4044 + _T_4046; // @[Bitwise.scala 48:55:@1976.4]
  assign _T_4048 = _T_4042 + _T_4047; // @[Bitwise.scala 48:55:@1977.4]
  assign _T_4049 = _T_4028 + _T_4029; // @[Bitwise.scala 48:55:@1978.4]
  assign _T_4050 = _T_4031 + _T_4032; // @[Bitwise.scala 48:55:@1979.4]
  assign _GEN_608 = {{1'd0}, _T_4030}; // @[Bitwise.scala 48:55:@1980.4]
  assign _T_4051 = _GEN_608 + _T_4050; // @[Bitwise.scala 48:55:@1980.4]
  assign _GEN_609 = {{1'd0}, _T_4049}; // @[Bitwise.scala 48:55:@1981.4]
  assign _T_4052 = _GEN_609 + _T_4051; // @[Bitwise.scala 48:55:@1981.4]
  assign _T_4053 = _T_4034 + _T_4035; // @[Bitwise.scala 48:55:@1982.4]
  assign _GEN_610 = {{1'd0}, _T_4033}; // @[Bitwise.scala 48:55:@1983.4]
  assign _T_4054 = _GEN_610 + _T_4053; // @[Bitwise.scala 48:55:@1983.4]
  assign _T_4055 = _T_4037 + _T_4038; // @[Bitwise.scala 48:55:@1984.4]
  assign _GEN_611 = {{1'd0}, _T_4036}; // @[Bitwise.scala 48:55:@1985.4]
  assign _T_4056 = _GEN_611 + _T_4055; // @[Bitwise.scala 48:55:@1985.4]
  assign _T_4057 = _T_4054 + _T_4056; // @[Bitwise.scala 48:55:@1986.4]
  assign _T_4058 = _T_4052 + _T_4057; // @[Bitwise.scala 48:55:@1987.4]
  assign _T_4059 = _T_4048 + _T_4058; // @[Bitwise.scala 48:55:@1988.4]
  assign _T_4123 = _T_2230[22:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2053.4]
  assign _T_4124 = _T_4123[0]; // @[Bitwise.scala 50:65:@2054.4]
  assign _T_4125 = _T_4123[1]; // @[Bitwise.scala 50:65:@2055.4]
  assign _T_4126 = _T_4123[2]; // @[Bitwise.scala 50:65:@2056.4]
  assign _T_4127 = _T_4123[3]; // @[Bitwise.scala 50:65:@2057.4]
  assign _T_4128 = _T_4123[4]; // @[Bitwise.scala 50:65:@2058.4]
  assign _T_4129 = _T_4123[5]; // @[Bitwise.scala 50:65:@2059.4]
  assign _T_4130 = _T_4123[6]; // @[Bitwise.scala 50:65:@2060.4]
  assign _T_4131 = _T_4123[7]; // @[Bitwise.scala 50:65:@2061.4]
  assign _T_4132 = _T_4123[8]; // @[Bitwise.scala 50:65:@2062.4]
  assign _T_4133 = _T_4123[9]; // @[Bitwise.scala 50:65:@2063.4]
  assign _T_4134 = _T_4123[10]; // @[Bitwise.scala 50:65:@2064.4]
  assign _T_4135 = _T_4123[11]; // @[Bitwise.scala 50:65:@2065.4]
  assign _T_4136 = _T_4123[12]; // @[Bitwise.scala 50:65:@2066.4]
  assign _T_4137 = _T_4123[13]; // @[Bitwise.scala 50:65:@2067.4]
  assign _T_4138 = _T_4123[14]; // @[Bitwise.scala 50:65:@2068.4]
  assign _T_4139 = _T_4123[15]; // @[Bitwise.scala 50:65:@2069.4]
  assign _T_4140 = _T_4123[16]; // @[Bitwise.scala 50:65:@2070.4]
  assign _T_4141 = _T_4123[17]; // @[Bitwise.scala 50:65:@2071.4]
  assign _T_4142 = _T_4123[18]; // @[Bitwise.scala 50:65:@2072.4]
  assign _T_4143 = _T_4123[19]; // @[Bitwise.scala 50:65:@2073.4]
  assign _T_4144 = _T_4123[20]; // @[Bitwise.scala 50:65:@2074.4]
  assign _T_4145 = _T_4123[21]; // @[Bitwise.scala 50:65:@2075.4]
  assign _T_4146 = _T_4123[22]; // @[Bitwise.scala 50:65:@2076.4]
  assign _T_4147 = _T_4124 + _T_4125; // @[Bitwise.scala 48:55:@2077.4]
  assign _T_4148 = _T_4127 + _T_4128; // @[Bitwise.scala 48:55:@2078.4]
  assign _GEN_612 = {{1'd0}, _T_4126}; // @[Bitwise.scala 48:55:@2079.4]
  assign _T_4149 = _GEN_612 + _T_4148; // @[Bitwise.scala 48:55:@2079.4]
  assign _GEN_613 = {{1'd0}, _T_4147}; // @[Bitwise.scala 48:55:@2080.4]
  assign _T_4150 = _GEN_613 + _T_4149; // @[Bitwise.scala 48:55:@2080.4]
  assign _T_4151 = _T_4130 + _T_4131; // @[Bitwise.scala 48:55:@2081.4]
  assign _GEN_614 = {{1'd0}, _T_4129}; // @[Bitwise.scala 48:55:@2082.4]
  assign _T_4152 = _GEN_614 + _T_4151; // @[Bitwise.scala 48:55:@2082.4]
  assign _T_4153 = _T_4133 + _T_4134; // @[Bitwise.scala 48:55:@2083.4]
  assign _GEN_615 = {{1'd0}, _T_4132}; // @[Bitwise.scala 48:55:@2084.4]
  assign _T_4154 = _GEN_615 + _T_4153; // @[Bitwise.scala 48:55:@2084.4]
  assign _T_4155 = _T_4152 + _T_4154; // @[Bitwise.scala 48:55:@2085.4]
  assign _T_4156 = _T_4150 + _T_4155; // @[Bitwise.scala 48:55:@2086.4]
  assign _T_4157 = _T_4136 + _T_4137; // @[Bitwise.scala 48:55:@2087.4]
  assign _GEN_616 = {{1'd0}, _T_4135}; // @[Bitwise.scala 48:55:@2088.4]
  assign _T_4158 = _GEN_616 + _T_4157; // @[Bitwise.scala 48:55:@2088.4]
  assign _T_4159 = _T_4139 + _T_4140; // @[Bitwise.scala 48:55:@2089.4]
  assign _GEN_617 = {{1'd0}, _T_4138}; // @[Bitwise.scala 48:55:@2090.4]
  assign _T_4160 = _GEN_617 + _T_4159; // @[Bitwise.scala 48:55:@2090.4]
  assign _T_4161 = _T_4158 + _T_4160; // @[Bitwise.scala 48:55:@2091.4]
  assign _T_4162 = _T_4142 + _T_4143; // @[Bitwise.scala 48:55:@2092.4]
  assign _GEN_618 = {{1'd0}, _T_4141}; // @[Bitwise.scala 48:55:@2093.4]
  assign _T_4163 = _GEN_618 + _T_4162; // @[Bitwise.scala 48:55:@2093.4]
  assign _T_4164 = _T_4145 + _T_4146; // @[Bitwise.scala 48:55:@2094.4]
  assign _GEN_619 = {{1'd0}, _T_4144}; // @[Bitwise.scala 48:55:@2095.4]
  assign _T_4165 = _GEN_619 + _T_4164; // @[Bitwise.scala 48:55:@2095.4]
  assign _T_4166 = _T_4163 + _T_4165; // @[Bitwise.scala 48:55:@2096.4]
  assign _T_4167 = _T_4161 + _T_4166; // @[Bitwise.scala 48:55:@2097.4]
  assign _T_4168 = _T_4156 + _T_4167; // @[Bitwise.scala 48:55:@2098.4]
  assign _T_4232 = _T_2230[23:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2163.4]
  assign _T_4233 = _T_4232[0]; // @[Bitwise.scala 50:65:@2164.4]
  assign _T_4234 = _T_4232[1]; // @[Bitwise.scala 50:65:@2165.4]
  assign _T_4235 = _T_4232[2]; // @[Bitwise.scala 50:65:@2166.4]
  assign _T_4236 = _T_4232[3]; // @[Bitwise.scala 50:65:@2167.4]
  assign _T_4237 = _T_4232[4]; // @[Bitwise.scala 50:65:@2168.4]
  assign _T_4238 = _T_4232[5]; // @[Bitwise.scala 50:65:@2169.4]
  assign _T_4239 = _T_4232[6]; // @[Bitwise.scala 50:65:@2170.4]
  assign _T_4240 = _T_4232[7]; // @[Bitwise.scala 50:65:@2171.4]
  assign _T_4241 = _T_4232[8]; // @[Bitwise.scala 50:65:@2172.4]
  assign _T_4242 = _T_4232[9]; // @[Bitwise.scala 50:65:@2173.4]
  assign _T_4243 = _T_4232[10]; // @[Bitwise.scala 50:65:@2174.4]
  assign _T_4244 = _T_4232[11]; // @[Bitwise.scala 50:65:@2175.4]
  assign _T_4245 = _T_4232[12]; // @[Bitwise.scala 50:65:@2176.4]
  assign _T_4246 = _T_4232[13]; // @[Bitwise.scala 50:65:@2177.4]
  assign _T_4247 = _T_4232[14]; // @[Bitwise.scala 50:65:@2178.4]
  assign _T_4248 = _T_4232[15]; // @[Bitwise.scala 50:65:@2179.4]
  assign _T_4249 = _T_4232[16]; // @[Bitwise.scala 50:65:@2180.4]
  assign _T_4250 = _T_4232[17]; // @[Bitwise.scala 50:65:@2181.4]
  assign _T_4251 = _T_4232[18]; // @[Bitwise.scala 50:65:@2182.4]
  assign _T_4252 = _T_4232[19]; // @[Bitwise.scala 50:65:@2183.4]
  assign _T_4253 = _T_4232[20]; // @[Bitwise.scala 50:65:@2184.4]
  assign _T_4254 = _T_4232[21]; // @[Bitwise.scala 50:65:@2185.4]
  assign _T_4255 = _T_4232[22]; // @[Bitwise.scala 50:65:@2186.4]
  assign _T_4256 = _T_4232[23]; // @[Bitwise.scala 50:65:@2187.4]
  assign _T_4257 = _T_4234 + _T_4235; // @[Bitwise.scala 48:55:@2188.4]
  assign _GEN_620 = {{1'd0}, _T_4233}; // @[Bitwise.scala 48:55:@2189.4]
  assign _T_4258 = _GEN_620 + _T_4257; // @[Bitwise.scala 48:55:@2189.4]
  assign _T_4259 = _T_4237 + _T_4238; // @[Bitwise.scala 48:55:@2190.4]
  assign _GEN_621 = {{1'd0}, _T_4236}; // @[Bitwise.scala 48:55:@2191.4]
  assign _T_4260 = _GEN_621 + _T_4259; // @[Bitwise.scala 48:55:@2191.4]
  assign _T_4261 = _T_4258 + _T_4260; // @[Bitwise.scala 48:55:@2192.4]
  assign _T_4262 = _T_4240 + _T_4241; // @[Bitwise.scala 48:55:@2193.4]
  assign _GEN_622 = {{1'd0}, _T_4239}; // @[Bitwise.scala 48:55:@2194.4]
  assign _T_4263 = _GEN_622 + _T_4262; // @[Bitwise.scala 48:55:@2194.4]
  assign _T_4264 = _T_4243 + _T_4244; // @[Bitwise.scala 48:55:@2195.4]
  assign _GEN_623 = {{1'd0}, _T_4242}; // @[Bitwise.scala 48:55:@2196.4]
  assign _T_4265 = _GEN_623 + _T_4264; // @[Bitwise.scala 48:55:@2196.4]
  assign _T_4266 = _T_4263 + _T_4265; // @[Bitwise.scala 48:55:@2197.4]
  assign _T_4267 = _T_4261 + _T_4266; // @[Bitwise.scala 48:55:@2198.4]
  assign _T_4268 = _T_4246 + _T_4247; // @[Bitwise.scala 48:55:@2199.4]
  assign _GEN_624 = {{1'd0}, _T_4245}; // @[Bitwise.scala 48:55:@2200.4]
  assign _T_4269 = _GEN_624 + _T_4268; // @[Bitwise.scala 48:55:@2200.4]
  assign _T_4270 = _T_4249 + _T_4250; // @[Bitwise.scala 48:55:@2201.4]
  assign _GEN_625 = {{1'd0}, _T_4248}; // @[Bitwise.scala 48:55:@2202.4]
  assign _T_4271 = _GEN_625 + _T_4270; // @[Bitwise.scala 48:55:@2202.4]
  assign _T_4272 = _T_4269 + _T_4271; // @[Bitwise.scala 48:55:@2203.4]
  assign _T_4273 = _T_4252 + _T_4253; // @[Bitwise.scala 48:55:@2204.4]
  assign _GEN_626 = {{1'd0}, _T_4251}; // @[Bitwise.scala 48:55:@2205.4]
  assign _T_4274 = _GEN_626 + _T_4273; // @[Bitwise.scala 48:55:@2205.4]
  assign _T_4275 = _T_4255 + _T_4256; // @[Bitwise.scala 48:55:@2206.4]
  assign _GEN_627 = {{1'd0}, _T_4254}; // @[Bitwise.scala 48:55:@2207.4]
  assign _T_4276 = _GEN_627 + _T_4275; // @[Bitwise.scala 48:55:@2207.4]
  assign _T_4277 = _T_4274 + _T_4276; // @[Bitwise.scala 48:55:@2208.4]
  assign _T_4278 = _T_4272 + _T_4277; // @[Bitwise.scala 48:55:@2209.4]
  assign _T_4279 = _T_4267 + _T_4278; // @[Bitwise.scala 48:55:@2210.4]
  assign _T_4343 = _T_2230[24:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2275.4]
  assign _T_4344 = _T_4343[0]; // @[Bitwise.scala 50:65:@2276.4]
  assign _T_4345 = _T_4343[1]; // @[Bitwise.scala 50:65:@2277.4]
  assign _T_4346 = _T_4343[2]; // @[Bitwise.scala 50:65:@2278.4]
  assign _T_4347 = _T_4343[3]; // @[Bitwise.scala 50:65:@2279.4]
  assign _T_4348 = _T_4343[4]; // @[Bitwise.scala 50:65:@2280.4]
  assign _T_4349 = _T_4343[5]; // @[Bitwise.scala 50:65:@2281.4]
  assign _T_4350 = _T_4343[6]; // @[Bitwise.scala 50:65:@2282.4]
  assign _T_4351 = _T_4343[7]; // @[Bitwise.scala 50:65:@2283.4]
  assign _T_4352 = _T_4343[8]; // @[Bitwise.scala 50:65:@2284.4]
  assign _T_4353 = _T_4343[9]; // @[Bitwise.scala 50:65:@2285.4]
  assign _T_4354 = _T_4343[10]; // @[Bitwise.scala 50:65:@2286.4]
  assign _T_4355 = _T_4343[11]; // @[Bitwise.scala 50:65:@2287.4]
  assign _T_4356 = _T_4343[12]; // @[Bitwise.scala 50:65:@2288.4]
  assign _T_4357 = _T_4343[13]; // @[Bitwise.scala 50:65:@2289.4]
  assign _T_4358 = _T_4343[14]; // @[Bitwise.scala 50:65:@2290.4]
  assign _T_4359 = _T_4343[15]; // @[Bitwise.scala 50:65:@2291.4]
  assign _T_4360 = _T_4343[16]; // @[Bitwise.scala 50:65:@2292.4]
  assign _T_4361 = _T_4343[17]; // @[Bitwise.scala 50:65:@2293.4]
  assign _T_4362 = _T_4343[18]; // @[Bitwise.scala 50:65:@2294.4]
  assign _T_4363 = _T_4343[19]; // @[Bitwise.scala 50:65:@2295.4]
  assign _T_4364 = _T_4343[20]; // @[Bitwise.scala 50:65:@2296.4]
  assign _T_4365 = _T_4343[21]; // @[Bitwise.scala 50:65:@2297.4]
  assign _T_4366 = _T_4343[22]; // @[Bitwise.scala 50:65:@2298.4]
  assign _T_4367 = _T_4343[23]; // @[Bitwise.scala 50:65:@2299.4]
  assign _T_4368 = _T_4343[24]; // @[Bitwise.scala 50:65:@2300.4]
  assign _T_4369 = _T_4345 + _T_4346; // @[Bitwise.scala 48:55:@2301.4]
  assign _GEN_628 = {{1'd0}, _T_4344}; // @[Bitwise.scala 48:55:@2302.4]
  assign _T_4370 = _GEN_628 + _T_4369; // @[Bitwise.scala 48:55:@2302.4]
  assign _T_4371 = _T_4348 + _T_4349; // @[Bitwise.scala 48:55:@2303.4]
  assign _GEN_629 = {{1'd0}, _T_4347}; // @[Bitwise.scala 48:55:@2304.4]
  assign _T_4372 = _GEN_629 + _T_4371; // @[Bitwise.scala 48:55:@2304.4]
  assign _T_4373 = _T_4370 + _T_4372; // @[Bitwise.scala 48:55:@2305.4]
  assign _T_4374 = _T_4351 + _T_4352; // @[Bitwise.scala 48:55:@2306.4]
  assign _GEN_630 = {{1'd0}, _T_4350}; // @[Bitwise.scala 48:55:@2307.4]
  assign _T_4375 = _GEN_630 + _T_4374; // @[Bitwise.scala 48:55:@2307.4]
  assign _T_4376 = _T_4354 + _T_4355; // @[Bitwise.scala 48:55:@2308.4]
  assign _GEN_631 = {{1'd0}, _T_4353}; // @[Bitwise.scala 48:55:@2309.4]
  assign _T_4377 = _GEN_631 + _T_4376; // @[Bitwise.scala 48:55:@2309.4]
  assign _T_4378 = _T_4375 + _T_4377; // @[Bitwise.scala 48:55:@2310.4]
  assign _T_4379 = _T_4373 + _T_4378; // @[Bitwise.scala 48:55:@2311.4]
  assign _T_4380 = _T_4357 + _T_4358; // @[Bitwise.scala 48:55:@2312.4]
  assign _GEN_632 = {{1'd0}, _T_4356}; // @[Bitwise.scala 48:55:@2313.4]
  assign _T_4381 = _GEN_632 + _T_4380; // @[Bitwise.scala 48:55:@2313.4]
  assign _T_4382 = _T_4360 + _T_4361; // @[Bitwise.scala 48:55:@2314.4]
  assign _GEN_633 = {{1'd0}, _T_4359}; // @[Bitwise.scala 48:55:@2315.4]
  assign _T_4383 = _GEN_633 + _T_4382; // @[Bitwise.scala 48:55:@2315.4]
  assign _T_4384 = _T_4381 + _T_4383; // @[Bitwise.scala 48:55:@2316.4]
  assign _T_4385 = _T_4363 + _T_4364; // @[Bitwise.scala 48:55:@2317.4]
  assign _GEN_634 = {{1'd0}, _T_4362}; // @[Bitwise.scala 48:55:@2318.4]
  assign _T_4386 = _GEN_634 + _T_4385; // @[Bitwise.scala 48:55:@2318.4]
  assign _T_4387 = _T_4365 + _T_4366; // @[Bitwise.scala 48:55:@2319.4]
  assign _T_4388 = _T_4367 + _T_4368; // @[Bitwise.scala 48:55:@2320.4]
  assign _T_4389 = _T_4387 + _T_4388; // @[Bitwise.scala 48:55:@2321.4]
  assign _T_4390 = _T_4386 + _T_4389; // @[Bitwise.scala 48:55:@2322.4]
  assign _T_4391 = _T_4384 + _T_4390; // @[Bitwise.scala 48:55:@2323.4]
  assign _T_4392 = _T_4379 + _T_4391; // @[Bitwise.scala 48:55:@2324.4]
  assign _T_4456 = _T_2230[25:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2389.4]
  assign _T_4457 = _T_4456[0]; // @[Bitwise.scala 50:65:@2390.4]
  assign _T_4458 = _T_4456[1]; // @[Bitwise.scala 50:65:@2391.4]
  assign _T_4459 = _T_4456[2]; // @[Bitwise.scala 50:65:@2392.4]
  assign _T_4460 = _T_4456[3]; // @[Bitwise.scala 50:65:@2393.4]
  assign _T_4461 = _T_4456[4]; // @[Bitwise.scala 50:65:@2394.4]
  assign _T_4462 = _T_4456[5]; // @[Bitwise.scala 50:65:@2395.4]
  assign _T_4463 = _T_4456[6]; // @[Bitwise.scala 50:65:@2396.4]
  assign _T_4464 = _T_4456[7]; // @[Bitwise.scala 50:65:@2397.4]
  assign _T_4465 = _T_4456[8]; // @[Bitwise.scala 50:65:@2398.4]
  assign _T_4466 = _T_4456[9]; // @[Bitwise.scala 50:65:@2399.4]
  assign _T_4467 = _T_4456[10]; // @[Bitwise.scala 50:65:@2400.4]
  assign _T_4468 = _T_4456[11]; // @[Bitwise.scala 50:65:@2401.4]
  assign _T_4469 = _T_4456[12]; // @[Bitwise.scala 50:65:@2402.4]
  assign _T_4470 = _T_4456[13]; // @[Bitwise.scala 50:65:@2403.4]
  assign _T_4471 = _T_4456[14]; // @[Bitwise.scala 50:65:@2404.4]
  assign _T_4472 = _T_4456[15]; // @[Bitwise.scala 50:65:@2405.4]
  assign _T_4473 = _T_4456[16]; // @[Bitwise.scala 50:65:@2406.4]
  assign _T_4474 = _T_4456[17]; // @[Bitwise.scala 50:65:@2407.4]
  assign _T_4475 = _T_4456[18]; // @[Bitwise.scala 50:65:@2408.4]
  assign _T_4476 = _T_4456[19]; // @[Bitwise.scala 50:65:@2409.4]
  assign _T_4477 = _T_4456[20]; // @[Bitwise.scala 50:65:@2410.4]
  assign _T_4478 = _T_4456[21]; // @[Bitwise.scala 50:65:@2411.4]
  assign _T_4479 = _T_4456[22]; // @[Bitwise.scala 50:65:@2412.4]
  assign _T_4480 = _T_4456[23]; // @[Bitwise.scala 50:65:@2413.4]
  assign _T_4481 = _T_4456[24]; // @[Bitwise.scala 50:65:@2414.4]
  assign _T_4482 = _T_4456[25]; // @[Bitwise.scala 50:65:@2415.4]
  assign _T_4483 = _T_4458 + _T_4459; // @[Bitwise.scala 48:55:@2416.4]
  assign _GEN_635 = {{1'd0}, _T_4457}; // @[Bitwise.scala 48:55:@2417.4]
  assign _T_4484 = _GEN_635 + _T_4483; // @[Bitwise.scala 48:55:@2417.4]
  assign _T_4485 = _T_4461 + _T_4462; // @[Bitwise.scala 48:55:@2418.4]
  assign _GEN_636 = {{1'd0}, _T_4460}; // @[Bitwise.scala 48:55:@2419.4]
  assign _T_4486 = _GEN_636 + _T_4485; // @[Bitwise.scala 48:55:@2419.4]
  assign _T_4487 = _T_4484 + _T_4486; // @[Bitwise.scala 48:55:@2420.4]
  assign _T_4488 = _T_4464 + _T_4465; // @[Bitwise.scala 48:55:@2421.4]
  assign _GEN_637 = {{1'd0}, _T_4463}; // @[Bitwise.scala 48:55:@2422.4]
  assign _T_4489 = _GEN_637 + _T_4488; // @[Bitwise.scala 48:55:@2422.4]
  assign _T_4490 = _T_4466 + _T_4467; // @[Bitwise.scala 48:55:@2423.4]
  assign _T_4491 = _T_4468 + _T_4469; // @[Bitwise.scala 48:55:@2424.4]
  assign _T_4492 = _T_4490 + _T_4491; // @[Bitwise.scala 48:55:@2425.4]
  assign _T_4493 = _T_4489 + _T_4492; // @[Bitwise.scala 48:55:@2426.4]
  assign _T_4494 = _T_4487 + _T_4493; // @[Bitwise.scala 48:55:@2427.4]
  assign _T_4495 = _T_4471 + _T_4472; // @[Bitwise.scala 48:55:@2428.4]
  assign _GEN_638 = {{1'd0}, _T_4470}; // @[Bitwise.scala 48:55:@2429.4]
  assign _T_4496 = _GEN_638 + _T_4495; // @[Bitwise.scala 48:55:@2429.4]
  assign _T_4497 = _T_4474 + _T_4475; // @[Bitwise.scala 48:55:@2430.4]
  assign _GEN_639 = {{1'd0}, _T_4473}; // @[Bitwise.scala 48:55:@2431.4]
  assign _T_4498 = _GEN_639 + _T_4497; // @[Bitwise.scala 48:55:@2431.4]
  assign _T_4499 = _T_4496 + _T_4498; // @[Bitwise.scala 48:55:@2432.4]
  assign _T_4500 = _T_4477 + _T_4478; // @[Bitwise.scala 48:55:@2433.4]
  assign _GEN_640 = {{1'd0}, _T_4476}; // @[Bitwise.scala 48:55:@2434.4]
  assign _T_4501 = _GEN_640 + _T_4500; // @[Bitwise.scala 48:55:@2434.4]
  assign _T_4502 = _T_4479 + _T_4480; // @[Bitwise.scala 48:55:@2435.4]
  assign _T_4503 = _T_4481 + _T_4482; // @[Bitwise.scala 48:55:@2436.4]
  assign _T_4504 = _T_4502 + _T_4503; // @[Bitwise.scala 48:55:@2437.4]
  assign _T_4505 = _T_4501 + _T_4504; // @[Bitwise.scala 48:55:@2438.4]
  assign _T_4506 = _T_4499 + _T_4505; // @[Bitwise.scala 48:55:@2439.4]
  assign _T_4507 = _T_4494 + _T_4506; // @[Bitwise.scala 48:55:@2440.4]
  assign _T_4571 = _T_2230[26:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2505.4]
  assign _T_4572 = _T_4571[0]; // @[Bitwise.scala 50:65:@2506.4]
  assign _T_4573 = _T_4571[1]; // @[Bitwise.scala 50:65:@2507.4]
  assign _T_4574 = _T_4571[2]; // @[Bitwise.scala 50:65:@2508.4]
  assign _T_4575 = _T_4571[3]; // @[Bitwise.scala 50:65:@2509.4]
  assign _T_4576 = _T_4571[4]; // @[Bitwise.scala 50:65:@2510.4]
  assign _T_4577 = _T_4571[5]; // @[Bitwise.scala 50:65:@2511.4]
  assign _T_4578 = _T_4571[6]; // @[Bitwise.scala 50:65:@2512.4]
  assign _T_4579 = _T_4571[7]; // @[Bitwise.scala 50:65:@2513.4]
  assign _T_4580 = _T_4571[8]; // @[Bitwise.scala 50:65:@2514.4]
  assign _T_4581 = _T_4571[9]; // @[Bitwise.scala 50:65:@2515.4]
  assign _T_4582 = _T_4571[10]; // @[Bitwise.scala 50:65:@2516.4]
  assign _T_4583 = _T_4571[11]; // @[Bitwise.scala 50:65:@2517.4]
  assign _T_4584 = _T_4571[12]; // @[Bitwise.scala 50:65:@2518.4]
  assign _T_4585 = _T_4571[13]; // @[Bitwise.scala 50:65:@2519.4]
  assign _T_4586 = _T_4571[14]; // @[Bitwise.scala 50:65:@2520.4]
  assign _T_4587 = _T_4571[15]; // @[Bitwise.scala 50:65:@2521.4]
  assign _T_4588 = _T_4571[16]; // @[Bitwise.scala 50:65:@2522.4]
  assign _T_4589 = _T_4571[17]; // @[Bitwise.scala 50:65:@2523.4]
  assign _T_4590 = _T_4571[18]; // @[Bitwise.scala 50:65:@2524.4]
  assign _T_4591 = _T_4571[19]; // @[Bitwise.scala 50:65:@2525.4]
  assign _T_4592 = _T_4571[20]; // @[Bitwise.scala 50:65:@2526.4]
  assign _T_4593 = _T_4571[21]; // @[Bitwise.scala 50:65:@2527.4]
  assign _T_4594 = _T_4571[22]; // @[Bitwise.scala 50:65:@2528.4]
  assign _T_4595 = _T_4571[23]; // @[Bitwise.scala 50:65:@2529.4]
  assign _T_4596 = _T_4571[24]; // @[Bitwise.scala 50:65:@2530.4]
  assign _T_4597 = _T_4571[25]; // @[Bitwise.scala 50:65:@2531.4]
  assign _T_4598 = _T_4571[26]; // @[Bitwise.scala 50:65:@2532.4]
  assign _T_4599 = _T_4573 + _T_4574; // @[Bitwise.scala 48:55:@2533.4]
  assign _GEN_641 = {{1'd0}, _T_4572}; // @[Bitwise.scala 48:55:@2534.4]
  assign _T_4600 = _GEN_641 + _T_4599; // @[Bitwise.scala 48:55:@2534.4]
  assign _T_4601 = _T_4576 + _T_4577; // @[Bitwise.scala 48:55:@2535.4]
  assign _GEN_642 = {{1'd0}, _T_4575}; // @[Bitwise.scala 48:55:@2536.4]
  assign _T_4602 = _GEN_642 + _T_4601; // @[Bitwise.scala 48:55:@2536.4]
  assign _T_4603 = _T_4600 + _T_4602; // @[Bitwise.scala 48:55:@2537.4]
  assign _T_4604 = _T_4579 + _T_4580; // @[Bitwise.scala 48:55:@2538.4]
  assign _GEN_643 = {{1'd0}, _T_4578}; // @[Bitwise.scala 48:55:@2539.4]
  assign _T_4605 = _GEN_643 + _T_4604; // @[Bitwise.scala 48:55:@2539.4]
  assign _T_4606 = _T_4581 + _T_4582; // @[Bitwise.scala 48:55:@2540.4]
  assign _T_4607 = _T_4583 + _T_4584; // @[Bitwise.scala 48:55:@2541.4]
  assign _T_4608 = _T_4606 + _T_4607; // @[Bitwise.scala 48:55:@2542.4]
  assign _T_4609 = _T_4605 + _T_4608; // @[Bitwise.scala 48:55:@2543.4]
  assign _T_4610 = _T_4603 + _T_4609; // @[Bitwise.scala 48:55:@2544.4]
  assign _T_4611 = _T_4586 + _T_4587; // @[Bitwise.scala 48:55:@2545.4]
  assign _GEN_644 = {{1'd0}, _T_4585}; // @[Bitwise.scala 48:55:@2546.4]
  assign _T_4612 = _GEN_644 + _T_4611; // @[Bitwise.scala 48:55:@2546.4]
  assign _T_4613 = _T_4588 + _T_4589; // @[Bitwise.scala 48:55:@2547.4]
  assign _T_4614 = _T_4590 + _T_4591; // @[Bitwise.scala 48:55:@2548.4]
  assign _T_4615 = _T_4613 + _T_4614; // @[Bitwise.scala 48:55:@2549.4]
  assign _T_4616 = _T_4612 + _T_4615; // @[Bitwise.scala 48:55:@2550.4]
  assign _T_4617 = _T_4593 + _T_4594; // @[Bitwise.scala 48:55:@2551.4]
  assign _GEN_645 = {{1'd0}, _T_4592}; // @[Bitwise.scala 48:55:@2552.4]
  assign _T_4618 = _GEN_645 + _T_4617; // @[Bitwise.scala 48:55:@2552.4]
  assign _T_4619 = _T_4595 + _T_4596; // @[Bitwise.scala 48:55:@2553.4]
  assign _T_4620 = _T_4597 + _T_4598; // @[Bitwise.scala 48:55:@2554.4]
  assign _T_4621 = _T_4619 + _T_4620; // @[Bitwise.scala 48:55:@2555.4]
  assign _T_4622 = _T_4618 + _T_4621; // @[Bitwise.scala 48:55:@2556.4]
  assign _T_4623 = _T_4616 + _T_4622; // @[Bitwise.scala 48:55:@2557.4]
  assign _T_4624 = _T_4610 + _T_4623; // @[Bitwise.scala 48:55:@2558.4]
  assign _T_4688 = _T_2230[27:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2623.4]
  assign _T_4689 = _T_4688[0]; // @[Bitwise.scala 50:65:@2624.4]
  assign _T_4690 = _T_4688[1]; // @[Bitwise.scala 50:65:@2625.4]
  assign _T_4691 = _T_4688[2]; // @[Bitwise.scala 50:65:@2626.4]
  assign _T_4692 = _T_4688[3]; // @[Bitwise.scala 50:65:@2627.4]
  assign _T_4693 = _T_4688[4]; // @[Bitwise.scala 50:65:@2628.4]
  assign _T_4694 = _T_4688[5]; // @[Bitwise.scala 50:65:@2629.4]
  assign _T_4695 = _T_4688[6]; // @[Bitwise.scala 50:65:@2630.4]
  assign _T_4696 = _T_4688[7]; // @[Bitwise.scala 50:65:@2631.4]
  assign _T_4697 = _T_4688[8]; // @[Bitwise.scala 50:65:@2632.4]
  assign _T_4698 = _T_4688[9]; // @[Bitwise.scala 50:65:@2633.4]
  assign _T_4699 = _T_4688[10]; // @[Bitwise.scala 50:65:@2634.4]
  assign _T_4700 = _T_4688[11]; // @[Bitwise.scala 50:65:@2635.4]
  assign _T_4701 = _T_4688[12]; // @[Bitwise.scala 50:65:@2636.4]
  assign _T_4702 = _T_4688[13]; // @[Bitwise.scala 50:65:@2637.4]
  assign _T_4703 = _T_4688[14]; // @[Bitwise.scala 50:65:@2638.4]
  assign _T_4704 = _T_4688[15]; // @[Bitwise.scala 50:65:@2639.4]
  assign _T_4705 = _T_4688[16]; // @[Bitwise.scala 50:65:@2640.4]
  assign _T_4706 = _T_4688[17]; // @[Bitwise.scala 50:65:@2641.4]
  assign _T_4707 = _T_4688[18]; // @[Bitwise.scala 50:65:@2642.4]
  assign _T_4708 = _T_4688[19]; // @[Bitwise.scala 50:65:@2643.4]
  assign _T_4709 = _T_4688[20]; // @[Bitwise.scala 50:65:@2644.4]
  assign _T_4710 = _T_4688[21]; // @[Bitwise.scala 50:65:@2645.4]
  assign _T_4711 = _T_4688[22]; // @[Bitwise.scala 50:65:@2646.4]
  assign _T_4712 = _T_4688[23]; // @[Bitwise.scala 50:65:@2647.4]
  assign _T_4713 = _T_4688[24]; // @[Bitwise.scala 50:65:@2648.4]
  assign _T_4714 = _T_4688[25]; // @[Bitwise.scala 50:65:@2649.4]
  assign _T_4715 = _T_4688[26]; // @[Bitwise.scala 50:65:@2650.4]
  assign _T_4716 = _T_4688[27]; // @[Bitwise.scala 50:65:@2651.4]
  assign _T_4717 = _T_4690 + _T_4691; // @[Bitwise.scala 48:55:@2652.4]
  assign _GEN_646 = {{1'd0}, _T_4689}; // @[Bitwise.scala 48:55:@2653.4]
  assign _T_4718 = _GEN_646 + _T_4717; // @[Bitwise.scala 48:55:@2653.4]
  assign _T_4719 = _T_4692 + _T_4693; // @[Bitwise.scala 48:55:@2654.4]
  assign _T_4720 = _T_4694 + _T_4695; // @[Bitwise.scala 48:55:@2655.4]
  assign _T_4721 = _T_4719 + _T_4720; // @[Bitwise.scala 48:55:@2656.4]
  assign _T_4722 = _T_4718 + _T_4721; // @[Bitwise.scala 48:55:@2657.4]
  assign _T_4723 = _T_4697 + _T_4698; // @[Bitwise.scala 48:55:@2658.4]
  assign _GEN_647 = {{1'd0}, _T_4696}; // @[Bitwise.scala 48:55:@2659.4]
  assign _T_4724 = _GEN_647 + _T_4723; // @[Bitwise.scala 48:55:@2659.4]
  assign _T_4725 = _T_4699 + _T_4700; // @[Bitwise.scala 48:55:@2660.4]
  assign _T_4726 = _T_4701 + _T_4702; // @[Bitwise.scala 48:55:@2661.4]
  assign _T_4727 = _T_4725 + _T_4726; // @[Bitwise.scala 48:55:@2662.4]
  assign _T_4728 = _T_4724 + _T_4727; // @[Bitwise.scala 48:55:@2663.4]
  assign _T_4729 = _T_4722 + _T_4728; // @[Bitwise.scala 48:55:@2664.4]
  assign _T_4730 = _T_4704 + _T_4705; // @[Bitwise.scala 48:55:@2665.4]
  assign _GEN_648 = {{1'd0}, _T_4703}; // @[Bitwise.scala 48:55:@2666.4]
  assign _T_4731 = _GEN_648 + _T_4730; // @[Bitwise.scala 48:55:@2666.4]
  assign _T_4732 = _T_4706 + _T_4707; // @[Bitwise.scala 48:55:@2667.4]
  assign _T_4733 = _T_4708 + _T_4709; // @[Bitwise.scala 48:55:@2668.4]
  assign _T_4734 = _T_4732 + _T_4733; // @[Bitwise.scala 48:55:@2669.4]
  assign _T_4735 = _T_4731 + _T_4734; // @[Bitwise.scala 48:55:@2670.4]
  assign _T_4736 = _T_4711 + _T_4712; // @[Bitwise.scala 48:55:@2671.4]
  assign _GEN_649 = {{1'd0}, _T_4710}; // @[Bitwise.scala 48:55:@2672.4]
  assign _T_4737 = _GEN_649 + _T_4736; // @[Bitwise.scala 48:55:@2672.4]
  assign _T_4738 = _T_4713 + _T_4714; // @[Bitwise.scala 48:55:@2673.4]
  assign _T_4739 = _T_4715 + _T_4716; // @[Bitwise.scala 48:55:@2674.4]
  assign _T_4740 = _T_4738 + _T_4739; // @[Bitwise.scala 48:55:@2675.4]
  assign _T_4741 = _T_4737 + _T_4740; // @[Bitwise.scala 48:55:@2676.4]
  assign _T_4742 = _T_4735 + _T_4741; // @[Bitwise.scala 48:55:@2677.4]
  assign _T_4743 = _T_4729 + _T_4742; // @[Bitwise.scala 48:55:@2678.4]
  assign _T_4807 = _T_2230[28:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2743.4]
  assign _T_4808 = _T_4807[0]; // @[Bitwise.scala 50:65:@2744.4]
  assign _T_4809 = _T_4807[1]; // @[Bitwise.scala 50:65:@2745.4]
  assign _T_4810 = _T_4807[2]; // @[Bitwise.scala 50:65:@2746.4]
  assign _T_4811 = _T_4807[3]; // @[Bitwise.scala 50:65:@2747.4]
  assign _T_4812 = _T_4807[4]; // @[Bitwise.scala 50:65:@2748.4]
  assign _T_4813 = _T_4807[5]; // @[Bitwise.scala 50:65:@2749.4]
  assign _T_4814 = _T_4807[6]; // @[Bitwise.scala 50:65:@2750.4]
  assign _T_4815 = _T_4807[7]; // @[Bitwise.scala 50:65:@2751.4]
  assign _T_4816 = _T_4807[8]; // @[Bitwise.scala 50:65:@2752.4]
  assign _T_4817 = _T_4807[9]; // @[Bitwise.scala 50:65:@2753.4]
  assign _T_4818 = _T_4807[10]; // @[Bitwise.scala 50:65:@2754.4]
  assign _T_4819 = _T_4807[11]; // @[Bitwise.scala 50:65:@2755.4]
  assign _T_4820 = _T_4807[12]; // @[Bitwise.scala 50:65:@2756.4]
  assign _T_4821 = _T_4807[13]; // @[Bitwise.scala 50:65:@2757.4]
  assign _T_4822 = _T_4807[14]; // @[Bitwise.scala 50:65:@2758.4]
  assign _T_4823 = _T_4807[15]; // @[Bitwise.scala 50:65:@2759.4]
  assign _T_4824 = _T_4807[16]; // @[Bitwise.scala 50:65:@2760.4]
  assign _T_4825 = _T_4807[17]; // @[Bitwise.scala 50:65:@2761.4]
  assign _T_4826 = _T_4807[18]; // @[Bitwise.scala 50:65:@2762.4]
  assign _T_4827 = _T_4807[19]; // @[Bitwise.scala 50:65:@2763.4]
  assign _T_4828 = _T_4807[20]; // @[Bitwise.scala 50:65:@2764.4]
  assign _T_4829 = _T_4807[21]; // @[Bitwise.scala 50:65:@2765.4]
  assign _T_4830 = _T_4807[22]; // @[Bitwise.scala 50:65:@2766.4]
  assign _T_4831 = _T_4807[23]; // @[Bitwise.scala 50:65:@2767.4]
  assign _T_4832 = _T_4807[24]; // @[Bitwise.scala 50:65:@2768.4]
  assign _T_4833 = _T_4807[25]; // @[Bitwise.scala 50:65:@2769.4]
  assign _T_4834 = _T_4807[26]; // @[Bitwise.scala 50:65:@2770.4]
  assign _T_4835 = _T_4807[27]; // @[Bitwise.scala 50:65:@2771.4]
  assign _T_4836 = _T_4807[28]; // @[Bitwise.scala 50:65:@2772.4]
  assign _T_4837 = _T_4809 + _T_4810; // @[Bitwise.scala 48:55:@2773.4]
  assign _GEN_650 = {{1'd0}, _T_4808}; // @[Bitwise.scala 48:55:@2774.4]
  assign _T_4838 = _GEN_650 + _T_4837; // @[Bitwise.scala 48:55:@2774.4]
  assign _T_4839 = _T_4811 + _T_4812; // @[Bitwise.scala 48:55:@2775.4]
  assign _T_4840 = _T_4813 + _T_4814; // @[Bitwise.scala 48:55:@2776.4]
  assign _T_4841 = _T_4839 + _T_4840; // @[Bitwise.scala 48:55:@2777.4]
  assign _T_4842 = _T_4838 + _T_4841; // @[Bitwise.scala 48:55:@2778.4]
  assign _T_4843 = _T_4816 + _T_4817; // @[Bitwise.scala 48:55:@2779.4]
  assign _GEN_651 = {{1'd0}, _T_4815}; // @[Bitwise.scala 48:55:@2780.4]
  assign _T_4844 = _GEN_651 + _T_4843; // @[Bitwise.scala 48:55:@2780.4]
  assign _T_4845 = _T_4818 + _T_4819; // @[Bitwise.scala 48:55:@2781.4]
  assign _T_4846 = _T_4820 + _T_4821; // @[Bitwise.scala 48:55:@2782.4]
  assign _T_4847 = _T_4845 + _T_4846; // @[Bitwise.scala 48:55:@2783.4]
  assign _T_4848 = _T_4844 + _T_4847; // @[Bitwise.scala 48:55:@2784.4]
  assign _T_4849 = _T_4842 + _T_4848; // @[Bitwise.scala 48:55:@2785.4]
  assign _T_4850 = _T_4823 + _T_4824; // @[Bitwise.scala 48:55:@2786.4]
  assign _GEN_652 = {{1'd0}, _T_4822}; // @[Bitwise.scala 48:55:@2787.4]
  assign _T_4851 = _GEN_652 + _T_4850; // @[Bitwise.scala 48:55:@2787.4]
  assign _T_4852 = _T_4825 + _T_4826; // @[Bitwise.scala 48:55:@2788.4]
  assign _T_4853 = _T_4827 + _T_4828; // @[Bitwise.scala 48:55:@2789.4]
  assign _T_4854 = _T_4852 + _T_4853; // @[Bitwise.scala 48:55:@2790.4]
  assign _T_4855 = _T_4851 + _T_4854; // @[Bitwise.scala 48:55:@2791.4]
  assign _T_4856 = _T_4829 + _T_4830; // @[Bitwise.scala 48:55:@2792.4]
  assign _T_4857 = _T_4831 + _T_4832; // @[Bitwise.scala 48:55:@2793.4]
  assign _T_4858 = _T_4856 + _T_4857; // @[Bitwise.scala 48:55:@2794.4]
  assign _T_4859 = _T_4833 + _T_4834; // @[Bitwise.scala 48:55:@2795.4]
  assign _T_4860 = _T_4835 + _T_4836; // @[Bitwise.scala 48:55:@2796.4]
  assign _T_4861 = _T_4859 + _T_4860; // @[Bitwise.scala 48:55:@2797.4]
  assign _T_4862 = _T_4858 + _T_4861; // @[Bitwise.scala 48:55:@2798.4]
  assign _T_4863 = _T_4855 + _T_4862; // @[Bitwise.scala 48:55:@2799.4]
  assign _T_4864 = _T_4849 + _T_4863; // @[Bitwise.scala 48:55:@2800.4]
  assign _T_4928 = _T_2230[29:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2865.4]
  assign _T_4929 = _T_4928[0]; // @[Bitwise.scala 50:65:@2866.4]
  assign _T_4930 = _T_4928[1]; // @[Bitwise.scala 50:65:@2867.4]
  assign _T_4931 = _T_4928[2]; // @[Bitwise.scala 50:65:@2868.4]
  assign _T_4932 = _T_4928[3]; // @[Bitwise.scala 50:65:@2869.4]
  assign _T_4933 = _T_4928[4]; // @[Bitwise.scala 50:65:@2870.4]
  assign _T_4934 = _T_4928[5]; // @[Bitwise.scala 50:65:@2871.4]
  assign _T_4935 = _T_4928[6]; // @[Bitwise.scala 50:65:@2872.4]
  assign _T_4936 = _T_4928[7]; // @[Bitwise.scala 50:65:@2873.4]
  assign _T_4937 = _T_4928[8]; // @[Bitwise.scala 50:65:@2874.4]
  assign _T_4938 = _T_4928[9]; // @[Bitwise.scala 50:65:@2875.4]
  assign _T_4939 = _T_4928[10]; // @[Bitwise.scala 50:65:@2876.4]
  assign _T_4940 = _T_4928[11]; // @[Bitwise.scala 50:65:@2877.4]
  assign _T_4941 = _T_4928[12]; // @[Bitwise.scala 50:65:@2878.4]
  assign _T_4942 = _T_4928[13]; // @[Bitwise.scala 50:65:@2879.4]
  assign _T_4943 = _T_4928[14]; // @[Bitwise.scala 50:65:@2880.4]
  assign _T_4944 = _T_4928[15]; // @[Bitwise.scala 50:65:@2881.4]
  assign _T_4945 = _T_4928[16]; // @[Bitwise.scala 50:65:@2882.4]
  assign _T_4946 = _T_4928[17]; // @[Bitwise.scala 50:65:@2883.4]
  assign _T_4947 = _T_4928[18]; // @[Bitwise.scala 50:65:@2884.4]
  assign _T_4948 = _T_4928[19]; // @[Bitwise.scala 50:65:@2885.4]
  assign _T_4949 = _T_4928[20]; // @[Bitwise.scala 50:65:@2886.4]
  assign _T_4950 = _T_4928[21]; // @[Bitwise.scala 50:65:@2887.4]
  assign _T_4951 = _T_4928[22]; // @[Bitwise.scala 50:65:@2888.4]
  assign _T_4952 = _T_4928[23]; // @[Bitwise.scala 50:65:@2889.4]
  assign _T_4953 = _T_4928[24]; // @[Bitwise.scala 50:65:@2890.4]
  assign _T_4954 = _T_4928[25]; // @[Bitwise.scala 50:65:@2891.4]
  assign _T_4955 = _T_4928[26]; // @[Bitwise.scala 50:65:@2892.4]
  assign _T_4956 = _T_4928[27]; // @[Bitwise.scala 50:65:@2893.4]
  assign _T_4957 = _T_4928[28]; // @[Bitwise.scala 50:65:@2894.4]
  assign _T_4958 = _T_4928[29]; // @[Bitwise.scala 50:65:@2895.4]
  assign _T_4959 = _T_4930 + _T_4931; // @[Bitwise.scala 48:55:@2896.4]
  assign _GEN_653 = {{1'd0}, _T_4929}; // @[Bitwise.scala 48:55:@2897.4]
  assign _T_4960 = _GEN_653 + _T_4959; // @[Bitwise.scala 48:55:@2897.4]
  assign _T_4961 = _T_4932 + _T_4933; // @[Bitwise.scala 48:55:@2898.4]
  assign _T_4962 = _T_4934 + _T_4935; // @[Bitwise.scala 48:55:@2899.4]
  assign _T_4963 = _T_4961 + _T_4962; // @[Bitwise.scala 48:55:@2900.4]
  assign _T_4964 = _T_4960 + _T_4963; // @[Bitwise.scala 48:55:@2901.4]
  assign _T_4965 = _T_4936 + _T_4937; // @[Bitwise.scala 48:55:@2902.4]
  assign _T_4966 = _T_4938 + _T_4939; // @[Bitwise.scala 48:55:@2903.4]
  assign _T_4967 = _T_4965 + _T_4966; // @[Bitwise.scala 48:55:@2904.4]
  assign _T_4968 = _T_4940 + _T_4941; // @[Bitwise.scala 48:55:@2905.4]
  assign _T_4969 = _T_4942 + _T_4943; // @[Bitwise.scala 48:55:@2906.4]
  assign _T_4970 = _T_4968 + _T_4969; // @[Bitwise.scala 48:55:@2907.4]
  assign _T_4971 = _T_4967 + _T_4970; // @[Bitwise.scala 48:55:@2908.4]
  assign _T_4972 = _T_4964 + _T_4971; // @[Bitwise.scala 48:55:@2909.4]
  assign _T_4973 = _T_4945 + _T_4946; // @[Bitwise.scala 48:55:@2910.4]
  assign _GEN_654 = {{1'd0}, _T_4944}; // @[Bitwise.scala 48:55:@2911.4]
  assign _T_4974 = _GEN_654 + _T_4973; // @[Bitwise.scala 48:55:@2911.4]
  assign _T_4975 = _T_4947 + _T_4948; // @[Bitwise.scala 48:55:@2912.4]
  assign _T_4976 = _T_4949 + _T_4950; // @[Bitwise.scala 48:55:@2913.4]
  assign _T_4977 = _T_4975 + _T_4976; // @[Bitwise.scala 48:55:@2914.4]
  assign _T_4978 = _T_4974 + _T_4977; // @[Bitwise.scala 48:55:@2915.4]
  assign _T_4979 = _T_4951 + _T_4952; // @[Bitwise.scala 48:55:@2916.4]
  assign _T_4980 = _T_4953 + _T_4954; // @[Bitwise.scala 48:55:@2917.4]
  assign _T_4981 = _T_4979 + _T_4980; // @[Bitwise.scala 48:55:@2918.4]
  assign _T_4982 = _T_4955 + _T_4956; // @[Bitwise.scala 48:55:@2919.4]
  assign _T_4983 = _T_4957 + _T_4958; // @[Bitwise.scala 48:55:@2920.4]
  assign _T_4984 = _T_4982 + _T_4983; // @[Bitwise.scala 48:55:@2921.4]
  assign _T_4985 = _T_4981 + _T_4984; // @[Bitwise.scala 48:55:@2922.4]
  assign _T_4986 = _T_4978 + _T_4985; // @[Bitwise.scala 48:55:@2923.4]
  assign _T_4987 = _T_4972 + _T_4986; // @[Bitwise.scala 48:55:@2924.4]
  assign _T_5051 = _T_2230[30:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@2989.4]
  assign _T_5052 = _T_5051[0]; // @[Bitwise.scala 50:65:@2990.4]
  assign _T_5053 = _T_5051[1]; // @[Bitwise.scala 50:65:@2991.4]
  assign _T_5054 = _T_5051[2]; // @[Bitwise.scala 50:65:@2992.4]
  assign _T_5055 = _T_5051[3]; // @[Bitwise.scala 50:65:@2993.4]
  assign _T_5056 = _T_5051[4]; // @[Bitwise.scala 50:65:@2994.4]
  assign _T_5057 = _T_5051[5]; // @[Bitwise.scala 50:65:@2995.4]
  assign _T_5058 = _T_5051[6]; // @[Bitwise.scala 50:65:@2996.4]
  assign _T_5059 = _T_5051[7]; // @[Bitwise.scala 50:65:@2997.4]
  assign _T_5060 = _T_5051[8]; // @[Bitwise.scala 50:65:@2998.4]
  assign _T_5061 = _T_5051[9]; // @[Bitwise.scala 50:65:@2999.4]
  assign _T_5062 = _T_5051[10]; // @[Bitwise.scala 50:65:@3000.4]
  assign _T_5063 = _T_5051[11]; // @[Bitwise.scala 50:65:@3001.4]
  assign _T_5064 = _T_5051[12]; // @[Bitwise.scala 50:65:@3002.4]
  assign _T_5065 = _T_5051[13]; // @[Bitwise.scala 50:65:@3003.4]
  assign _T_5066 = _T_5051[14]; // @[Bitwise.scala 50:65:@3004.4]
  assign _T_5067 = _T_5051[15]; // @[Bitwise.scala 50:65:@3005.4]
  assign _T_5068 = _T_5051[16]; // @[Bitwise.scala 50:65:@3006.4]
  assign _T_5069 = _T_5051[17]; // @[Bitwise.scala 50:65:@3007.4]
  assign _T_5070 = _T_5051[18]; // @[Bitwise.scala 50:65:@3008.4]
  assign _T_5071 = _T_5051[19]; // @[Bitwise.scala 50:65:@3009.4]
  assign _T_5072 = _T_5051[20]; // @[Bitwise.scala 50:65:@3010.4]
  assign _T_5073 = _T_5051[21]; // @[Bitwise.scala 50:65:@3011.4]
  assign _T_5074 = _T_5051[22]; // @[Bitwise.scala 50:65:@3012.4]
  assign _T_5075 = _T_5051[23]; // @[Bitwise.scala 50:65:@3013.4]
  assign _T_5076 = _T_5051[24]; // @[Bitwise.scala 50:65:@3014.4]
  assign _T_5077 = _T_5051[25]; // @[Bitwise.scala 50:65:@3015.4]
  assign _T_5078 = _T_5051[26]; // @[Bitwise.scala 50:65:@3016.4]
  assign _T_5079 = _T_5051[27]; // @[Bitwise.scala 50:65:@3017.4]
  assign _T_5080 = _T_5051[28]; // @[Bitwise.scala 50:65:@3018.4]
  assign _T_5081 = _T_5051[29]; // @[Bitwise.scala 50:65:@3019.4]
  assign _T_5082 = _T_5051[30]; // @[Bitwise.scala 50:65:@3020.4]
  assign _T_5083 = _T_5053 + _T_5054; // @[Bitwise.scala 48:55:@3021.4]
  assign _GEN_655 = {{1'd0}, _T_5052}; // @[Bitwise.scala 48:55:@3022.4]
  assign _T_5084 = _GEN_655 + _T_5083; // @[Bitwise.scala 48:55:@3022.4]
  assign _T_5085 = _T_5055 + _T_5056; // @[Bitwise.scala 48:55:@3023.4]
  assign _T_5086 = _T_5057 + _T_5058; // @[Bitwise.scala 48:55:@3024.4]
  assign _T_5087 = _T_5085 + _T_5086; // @[Bitwise.scala 48:55:@3025.4]
  assign _T_5088 = _T_5084 + _T_5087; // @[Bitwise.scala 48:55:@3026.4]
  assign _T_5089 = _T_5059 + _T_5060; // @[Bitwise.scala 48:55:@3027.4]
  assign _T_5090 = _T_5061 + _T_5062; // @[Bitwise.scala 48:55:@3028.4]
  assign _T_5091 = _T_5089 + _T_5090; // @[Bitwise.scala 48:55:@3029.4]
  assign _T_5092 = _T_5063 + _T_5064; // @[Bitwise.scala 48:55:@3030.4]
  assign _T_5093 = _T_5065 + _T_5066; // @[Bitwise.scala 48:55:@3031.4]
  assign _T_5094 = _T_5092 + _T_5093; // @[Bitwise.scala 48:55:@3032.4]
  assign _T_5095 = _T_5091 + _T_5094; // @[Bitwise.scala 48:55:@3033.4]
  assign _T_5096 = _T_5088 + _T_5095; // @[Bitwise.scala 48:55:@3034.4]
  assign _T_5097 = _T_5067 + _T_5068; // @[Bitwise.scala 48:55:@3035.4]
  assign _T_5098 = _T_5069 + _T_5070; // @[Bitwise.scala 48:55:@3036.4]
  assign _T_5099 = _T_5097 + _T_5098; // @[Bitwise.scala 48:55:@3037.4]
  assign _T_5100 = _T_5071 + _T_5072; // @[Bitwise.scala 48:55:@3038.4]
  assign _T_5101 = _T_5073 + _T_5074; // @[Bitwise.scala 48:55:@3039.4]
  assign _T_5102 = _T_5100 + _T_5101; // @[Bitwise.scala 48:55:@3040.4]
  assign _T_5103 = _T_5099 + _T_5102; // @[Bitwise.scala 48:55:@3041.4]
  assign _T_5104 = _T_5075 + _T_5076; // @[Bitwise.scala 48:55:@3042.4]
  assign _T_5105 = _T_5077 + _T_5078; // @[Bitwise.scala 48:55:@3043.4]
  assign _T_5106 = _T_5104 + _T_5105; // @[Bitwise.scala 48:55:@3044.4]
  assign _T_5107 = _T_5079 + _T_5080; // @[Bitwise.scala 48:55:@3045.4]
  assign _T_5108 = _T_5081 + _T_5082; // @[Bitwise.scala 48:55:@3046.4]
  assign _T_5109 = _T_5107 + _T_5108; // @[Bitwise.scala 48:55:@3047.4]
  assign _T_5110 = _T_5106 + _T_5109; // @[Bitwise.scala 48:55:@3048.4]
  assign _T_5111 = _T_5103 + _T_5110; // @[Bitwise.scala 48:55:@3049.4]
  assign _T_5112 = _T_5096 + _T_5111; // @[Bitwise.scala 48:55:@3050.4]
  assign _T_5176 = _T_2230[31:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3115.4]
  assign _T_5177 = _T_5176[0]; // @[Bitwise.scala 50:65:@3116.4]
  assign _T_5178 = _T_5176[1]; // @[Bitwise.scala 50:65:@3117.4]
  assign _T_5179 = _T_5176[2]; // @[Bitwise.scala 50:65:@3118.4]
  assign _T_5180 = _T_5176[3]; // @[Bitwise.scala 50:65:@3119.4]
  assign _T_5181 = _T_5176[4]; // @[Bitwise.scala 50:65:@3120.4]
  assign _T_5182 = _T_5176[5]; // @[Bitwise.scala 50:65:@3121.4]
  assign _T_5183 = _T_5176[6]; // @[Bitwise.scala 50:65:@3122.4]
  assign _T_5184 = _T_5176[7]; // @[Bitwise.scala 50:65:@3123.4]
  assign _T_5185 = _T_5176[8]; // @[Bitwise.scala 50:65:@3124.4]
  assign _T_5186 = _T_5176[9]; // @[Bitwise.scala 50:65:@3125.4]
  assign _T_5187 = _T_5176[10]; // @[Bitwise.scala 50:65:@3126.4]
  assign _T_5188 = _T_5176[11]; // @[Bitwise.scala 50:65:@3127.4]
  assign _T_5189 = _T_5176[12]; // @[Bitwise.scala 50:65:@3128.4]
  assign _T_5190 = _T_5176[13]; // @[Bitwise.scala 50:65:@3129.4]
  assign _T_5191 = _T_5176[14]; // @[Bitwise.scala 50:65:@3130.4]
  assign _T_5192 = _T_5176[15]; // @[Bitwise.scala 50:65:@3131.4]
  assign _T_5193 = _T_5176[16]; // @[Bitwise.scala 50:65:@3132.4]
  assign _T_5194 = _T_5176[17]; // @[Bitwise.scala 50:65:@3133.4]
  assign _T_5195 = _T_5176[18]; // @[Bitwise.scala 50:65:@3134.4]
  assign _T_5196 = _T_5176[19]; // @[Bitwise.scala 50:65:@3135.4]
  assign _T_5197 = _T_5176[20]; // @[Bitwise.scala 50:65:@3136.4]
  assign _T_5198 = _T_5176[21]; // @[Bitwise.scala 50:65:@3137.4]
  assign _T_5199 = _T_5176[22]; // @[Bitwise.scala 50:65:@3138.4]
  assign _T_5200 = _T_5176[23]; // @[Bitwise.scala 50:65:@3139.4]
  assign _T_5201 = _T_5176[24]; // @[Bitwise.scala 50:65:@3140.4]
  assign _T_5202 = _T_5176[25]; // @[Bitwise.scala 50:65:@3141.4]
  assign _T_5203 = _T_5176[26]; // @[Bitwise.scala 50:65:@3142.4]
  assign _T_5204 = _T_5176[27]; // @[Bitwise.scala 50:65:@3143.4]
  assign _T_5205 = _T_5176[28]; // @[Bitwise.scala 50:65:@3144.4]
  assign _T_5206 = _T_5176[29]; // @[Bitwise.scala 50:65:@3145.4]
  assign _T_5207 = _T_5176[30]; // @[Bitwise.scala 50:65:@3146.4]
  assign _T_5208 = _T_5176[31]; // @[Bitwise.scala 50:65:@3147.4]
  assign _T_5209 = _T_5177 + _T_5178; // @[Bitwise.scala 48:55:@3148.4]
  assign _T_5210 = _T_5179 + _T_5180; // @[Bitwise.scala 48:55:@3149.4]
  assign _T_5211 = _T_5209 + _T_5210; // @[Bitwise.scala 48:55:@3150.4]
  assign _T_5212 = _T_5181 + _T_5182; // @[Bitwise.scala 48:55:@3151.4]
  assign _T_5213 = _T_5183 + _T_5184; // @[Bitwise.scala 48:55:@3152.4]
  assign _T_5214 = _T_5212 + _T_5213; // @[Bitwise.scala 48:55:@3153.4]
  assign _T_5215 = _T_5211 + _T_5214; // @[Bitwise.scala 48:55:@3154.4]
  assign _T_5216 = _T_5185 + _T_5186; // @[Bitwise.scala 48:55:@3155.4]
  assign _T_5217 = _T_5187 + _T_5188; // @[Bitwise.scala 48:55:@3156.4]
  assign _T_5218 = _T_5216 + _T_5217; // @[Bitwise.scala 48:55:@3157.4]
  assign _T_5219 = _T_5189 + _T_5190; // @[Bitwise.scala 48:55:@3158.4]
  assign _T_5220 = _T_5191 + _T_5192; // @[Bitwise.scala 48:55:@3159.4]
  assign _T_5221 = _T_5219 + _T_5220; // @[Bitwise.scala 48:55:@3160.4]
  assign _T_5222 = _T_5218 + _T_5221; // @[Bitwise.scala 48:55:@3161.4]
  assign _T_5223 = _T_5215 + _T_5222; // @[Bitwise.scala 48:55:@3162.4]
  assign _T_5224 = _T_5193 + _T_5194; // @[Bitwise.scala 48:55:@3163.4]
  assign _T_5225 = _T_5195 + _T_5196; // @[Bitwise.scala 48:55:@3164.4]
  assign _T_5226 = _T_5224 + _T_5225; // @[Bitwise.scala 48:55:@3165.4]
  assign _T_5227 = _T_5197 + _T_5198; // @[Bitwise.scala 48:55:@3166.4]
  assign _T_5228 = _T_5199 + _T_5200; // @[Bitwise.scala 48:55:@3167.4]
  assign _T_5229 = _T_5227 + _T_5228; // @[Bitwise.scala 48:55:@3168.4]
  assign _T_5230 = _T_5226 + _T_5229; // @[Bitwise.scala 48:55:@3169.4]
  assign _T_5231 = _T_5201 + _T_5202; // @[Bitwise.scala 48:55:@3170.4]
  assign _T_5232 = _T_5203 + _T_5204; // @[Bitwise.scala 48:55:@3171.4]
  assign _T_5233 = _T_5231 + _T_5232; // @[Bitwise.scala 48:55:@3172.4]
  assign _T_5234 = _T_5205 + _T_5206; // @[Bitwise.scala 48:55:@3173.4]
  assign _T_5235 = _T_5207 + _T_5208; // @[Bitwise.scala 48:55:@3174.4]
  assign _T_5236 = _T_5234 + _T_5235; // @[Bitwise.scala 48:55:@3175.4]
  assign _T_5237 = _T_5233 + _T_5236; // @[Bitwise.scala 48:55:@3176.4]
  assign _T_5238 = _T_5230 + _T_5237; // @[Bitwise.scala 48:55:@3177.4]
  assign _T_5239 = _T_5223 + _T_5238; // @[Bitwise.scala 48:55:@3178.4]
  assign _T_5303 = _T_2230[32:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3243.4]
  assign _T_5304 = _T_5303[0]; // @[Bitwise.scala 50:65:@3244.4]
  assign _T_5305 = _T_5303[1]; // @[Bitwise.scala 50:65:@3245.4]
  assign _T_5306 = _T_5303[2]; // @[Bitwise.scala 50:65:@3246.4]
  assign _T_5307 = _T_5303[3]; // @[Bitwise.scala 50:65:@3247.4]
  assign _T_5308 = _T_5303[4]; // @[Bitwise.scala 50:65:@3248.4]
  assign _T_5309 = _T_5303[5]; // @[Bitwise.scala 50:65:@3249.4]
  assign _T_5310 = _T_5303[6]; // @[Bitwise.scala 50:65:@3250.4]
  assign _T_5311 = _T_5303[7]; // @[Bitwise.scala 50:65:@3251.4]
  assign _T_5312 = _T_5303[8]; // @[Bitwise.scala 50:65:@3252.4]
  assign _T_5313 = _T_5303[9]; // @[Bitwise.scala 50:65:@3253.4]
  assign _T_5314 = _T_5303[10]; // @[Bitwise.scala 50:65:@3254.4]
  assign _T_5315 = _T_5303[11]; // @[Bitwise.scala 50:65:@3255.4]
  assign _T_5316 = _T_5303[12]; // @[Bitwise.scala 50:65:@3256.4]
  assign _T_5317 = _T_5303[13]; // @[Bitwise.scala 50:65:@3257.4]
  assign _T_5318 = _T_5303[14]; // @[Bitwise.scala 50:65:@3258.4]
  assign _T_5319 = _T_5303[15]; // @[Bitwise.scala 50:65:@3259.4]
  assign _T_5320 = _T_5303[16]; // @[Bitwise.scala 50:65:@3260.4]
  assign _T_5321 = _T_5303[17]; // @[Bitwise.scala 50:65:@3261.4]
  assign _T_5322 = _T_5303[18]; // @[Bitwise.scala 50:65:@3262.4]
  assign _T_5323 = _T_5303[19]; // @[Bitwise.scala 50:65:@3263.4]
  assign _T_5324 = _T_5303[20]; // @[Bitwise.scala 50:65:@3264.4]
  assign _T_5325 = _T_5303[21]; // @[Bitwise.scala 50:65:@3265.4]
  assign _T_5326 = _T_5303[22]; // @[Bitwise.scala 50:65:@3266.4]
  assign _T_5327 = _T_5303[23]; // @[Bitwise.scala 50:65:@3267.4]
  assign _T_5328 = _T_5303[24]; // @[Bitwise.scala 50:65:@3268.4]
  assign _T_5329 = _T_5303[25]; // @[Bitwise.scala 50:65:@3269.4]
  assign _T_5330 = _T_5303[26]; // @[Bitwise.scala 50:65:@3270.4]
  assign _T_5331 = _T_5303[27]; // @[Bitwise.scala 50:65:@3271.4]
  assign _T_5332 = _T_5303[28]; // @[Bitwise.scala 50:65:@3272.4]
  assign _T_5333 = _T_5303[29]; // @[Bitwise.scala 50:65:@3273.4]
  assign _T_5334 = _T_5303[30]; // @[Bitwise.scala 50:65:@3274.4]
  assign _T_5335 = _T_5303[31]; // @[Bitwise.scala 50:65:@3275.4]
  assign _T_5336 = _T_5303[32]; // @[Bitwise.scala 50:65:@3276.4]
  assign _T_5337 = _T_5304 + _T_5305; // @[Bitwise.scala 48:55:@3277.4]
  assign _T_5338 = _T_5306 + _T_5307; // @[Bitwise.scala 48:55:@3278.4]
  assign _T_5339 = _T_5337 + _T_5338; // @[Bitwise.scala 48:55:@3279.4]
  assign _T_5340 = _T_5308 + _T_5309; // @[Bitwise.scala 48:55:@3280.4]
  assign _T_5341 = _T_5310 + _T_5311; // @[Bitwise.scala 48:55:@3281.4]
  assign _T_5342 = _T_5340 + _T_5341; // @[Bitwise.scala 48:55:@3282.4]
  assign _T_5343 = _T_5339 + _T_5342; // @[Bitwise.scala 48:55:@3283.4]
  assign _T_5344 = _T_5312 + _T_5313; // @[Bitwise.scala 48:55:@3284.4]
  assign _T_5345 = _T_5314 + _T_5315; // @[Bitwise.scala 48:55:@3285.4]
  assign _T_5346 = _T_5344 + _T_5345; // @[Bitwise.scala 48:55:@3286.4]
  assign _T_5347 = _T_5316 + _T_5317; // @[Bitwise.scala 48:55:@3287.4]
  assign _T_5348 = _T_5318 + _T_5319; // @[Bitwise.scala 48:55:@3288.4]
  assign _T_5349 = _T_5347 + _T_5348; // @[Bitwise.scala 48:55:@3289.4]
  assign _T_5350 = _T_5346 + _T_5349; // @[Bitwise.scala 48:55:@3290.4]
  assign _T_5351 = _T_5343 + _T_5350; // @[Bitwise.scala 48:55:@3291.4]
  assign _T_5352 = _T_5320 + _T_5321; // @[Bitwise.scala 48:55:@3292.4]
  assign _T_5353 = _T_5322 + _T_5323; // @[Bitwise.scala 48:55:@3293.4]
  assign _T_5354 = _T_5352 + _T_5353; // @[Bitwise.scala 48:55:@3294.4]
  assign _T_5355 = _T_5324 + _T_5325; // @[Bitwise.scala 48:55:@3295.4]
  assign _T_5356 = _T_5326 + _T_5327; // @[Bitwise.scala 48:55:@3296.4]
  assign _T_5357 = _T_5355 + _T_5356; // @[Bitwise.scala 48:55:@3297.4]
  assign _T_5358 = _T_5354 + _T_5357; // @[Bitwise.scala 48:55:@3298.4]
  assign _T_5359 = _T_5328 + _T_5329; // @[Bitwise.scala 48:55:@3299.4]
  assign _T_5360 = _T_5330 + _T_5331; // @[Bitwise.scala 48:55:@3300.4]
  assign _T_5361 = _T_5359 + _T_5360; // @[Bitwise.scala 48:55:@3301.4]
  assign _T_5362 = _T_5332 + _T_5333; // @[Bitwise.scala 48:55:@3302.4]
  assign _T_5363 = _T_5335 + _T_5336; // @[Bitwise.scala 48:55:@3303.4]
  assign _GEN_656 = {{1'd0}, _T_5334}; // @[Bitwise.scala 48:55:@3304.4]
  assign _T_5364 = _GEN_656 + _T_5363; // @[Bitwise.scala 48:55:@3304.4]
  assign _GEN_657 = {{1'd0}, _T_5362}; // @[Bitwise.scala 48:55:@3305.4]
  assign _T_5365 = _GEN_657 + _T_5364; // @[Bitwise.scala 48:55:@3305.4]
  assign _GEN_658 = {{1'd0}, _T_5361}; // @[Bitwise.scala 48:55:@3306.4]
  assign _T_5366 = _GEN_658 + _T_5365; // @[Bitwise.scala 48:55:@3306.4]
  assign _GEN_659 = {{1'd0}, _T_5358}; // @[Bitwise.scala 48:55:@3307.4]
  assign _T_5367 = _GEN_659 + _T_5366; // @[Bitwise.scala 48:55:@3307.4]
  assign _GEN_660 = {{1'd0}, _T_5351}; // @[Bitwise.scala 48:55:@3308.4]
  assign _T_5368 = _GEN_660 + _T_5367; // @[Bitwise.scala 48:55:@3308.4]
  assign _T_5432 = _T_2230[33:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3373.4]
  assign _T_5433 = _T_5432[0]; // @[Bitwise.scala 50:65:@3374.4]
  assign _T_5434 = _T_5432[1]; // @[Bitwise.scala 50:65:@3375.4]
  assign _T_5435 = _T_5432[2]; // @[Bitwise.scala 50:65:@3376.4]
  assign _T_5436 = _T_5432[3]; // @[Bitwise.scala 50:65:@3377.4]
  assign _T_5437 = _T_5432[4]; // @[Bitwise.scala 50:65:@3378.4]
  assign _T_5438 = _T_5432[5]; // @[Bitwise.scala 50:65:@3379.4]
  assign _T_5439 = _T_5432[6]; // @[Bitwise.scala 50:65:@3380.4]
  assign _T_5440 = _T_5432[7]; // @[Bitwise.scala 50:65:@3381.4]
  assign _T_5441 = _T_5432[8]; // @[Bitwise.scala 50:65:@3382.4]
  assign _T_5442 = _T_5432[9]; // @[Bitwise.scala 50:65:@3383.4]
  assign _T_5443 = _T_5432[10]; // @[Bitwise.scala 50:65:@3384.4]
  assign _T_5444 = _T_5432[11]; // @[Bitwise.scala 50:65:@3385.4]
  assign _T_5445 = _T_5432[12]; // @[Bitwise.scala 50:65:@3386.4]
  assign _T_5446 = _T_5432[13]; // @[Bitwise.scala 50:65:@3387.4]
  assign _T_5447 = _T_5432[14]; // @[Bitwise.scala 50:65:@3388.4]
  assign _T_5448 = _T_5432[15]; // @[Bitwise.scala 50:65:@3389.4]
  assign _T_5449 = _T_5432[16]; // @[Bitwise.scala 50:65:@3390.4]
  assign _T_5450 = _T_5432[17]; // @[Bitwise.scala 50:65:@3391.4]
  assign _T_5451 = _T_5432[18]; // @[Bitwise.scala 50:65:@3392.4]
  assign _T_5452 = _T_5432[19]; // @[Bitwise.scala 50:65:@3393.4]
  assign _T_5453 = _T_5432[20]; // @[Bitwise.scala 50:65:@3394.4]
  assign _T_5454 = _T_5432[21]; // @[Bitwise.scala 50:65:@3395.4]
  assign _T_5455 = _T_5432[22]; // @[Bitwise.scala 50:65:@3396.4]
  assign _T_5456 = _T_5432[23]; // @[Bitwise.scala 50:65:@3397.4]
  assign _T_5457 = _T_5432[24]; // @[Bitwise.scala 50:65:@3398.4]
  assign _T_5458 = _T_5432[25]; // @[Bitwise.scala 50:65:@3399.4]
  assign _T_5459 = _T_5432[26]; // @[Bitwise.scala 50:65:@3400.4]
  assign _T_5460 = _T_5432[27]; // @[Bitwise.scala 50:65:@3401.4]
  assign _T_5461 = _T_5432[28]; // @[Bitwise.scala 50:65:@3402.4]
  assign _T_5462 = _T_5432[29]; // @[Bitwise.scala 50:65:@3403.4]
  assign _T_5463 = _T_5432[30]; // @[Bitwise.scala 50:65:@3404.4]
  assign _T_5464 = _T_5432[31]; // @[Bitwise.scala 50:65:@3405.4]
  assign _T_5465 = _T_5432[32]; // @[Bitwise.scala 50:65:@3406.4]
  assign _T_5466 = _T_5432[33]; // @[Bitwise.scala 50:65:@3407.4]
  assign _T_5467 = _T_5433 + _T_5434; // @[Bitwise.scala 48:55:@3408.4]
  assign _T_5468 = _T_5435 + _T_5436; // @[Bitwise.scala 48:55:@3409.4]
  assign _T_5469 = _T_5467 + _T_5468; // @[Bitwise.scala 48:55:@3410.4]
  assign _T_5470 = _T_5437 + _T_5438; // @[Bitwise.scala 48:55:@3411.4]
  assign _T_5471 = _T_5439 + _T_5440; // @[Bitwise.scala 48:55:@3412.4]
  assign _T_5472 = _T_5470 + _T_5471; // @[Bitwise.scala 48:55:@3413.4]
  assign _T_5473 = _T_5469 + _T_5472; // @[Bitwise.scala 48:55:@3414.4]
  assign _T_5474 = _T_5441 + _T_5442; // @[Bitwise.scala 48:55:@3415.4]
  assign _T_5475 = _T_5443 + _T_5444; // @[Bitwise.scala 48:55:@3416.4]
  assign _T_5476 = _T_5474 + _T_5475; // @[Bitwise.scala 48:55:@3417.4]
  assign _T_5477 = _T_5445 + _T_5446; // @[Bitwise.scala 48:55:@3418.4]
  assign _T_5478 = _T_5448 + _T_5449; // @[Bitwise.scala 48:55:@3419.4]
  assign _GEN_661 = {{1'd0}, _T_5447}; // @[Bitwise.scala 48:55:@3420.4]
  assign _T_5479 = _GEN_661 + _T_5478; // @[Bitwise.scala 48:55:@3420.4]
  assign _GEN_662 = {{1'd0}, _T_5477}; // @[Bitwise.scala 48:55:@3421.4]
  assign _T_5480 = _GEN_662 + _T_5479; // @[Bitwise.scala 48:55:@3421.4]
  assign _GEN_663 = {{1'd0}, _T_5476}; // @[Bitwise.scala 48:55:@3422.4]
  assign _T_5481 = _GEN_663 + _T_5480; // @[Bitwise.scala 48:55:@3422.4]
  assign _GEN_664 = {{1'd0}, _T_5473}; // @[Bitwise.scala 48:55:@3423.4]
  assign _T_5482 = _GEN_664 + _T_5481; // @[Bitwise.scala 48:55:@3423.4]
  assign _T_5483 = _T_5450 + _T_5451; // @[Bitwise.scala 48:55:@3424.4]
  assign _T_5484 = _T_5452 + _T_5453; // @[Bitwise.scala 48:55:@3425.4]
  assign _T_5485 = _T_5483 + _T_5484; // @[Bitwise.scala 48:55:@3426.4]
  assign _T_5486 = _T_5454 + _T_5455; // @[Bitwise.scala 48:55:@3427.4]
  assign _T_5487 = _T_5456 + _T_5457; // @[Bitwise.scala 48:55:@3428.4]
  assign _T_5488 = _T_5486 + _T_5487; // @[Bitwise.scala 48:55:@3429.4]
  assign _T_5489 = _T_5485 + _T_5488; // @[Bitwise.scala 48:55:@3430.4]
  assign _T_5490 = _T_5458 + _T_5459; // @[Bitwise.scala 48:55:@3431.4]
  assign _T_5491 = _T_5460 + _T_5461; // @[Bitwise.scala 48:55:@3432.4]
  assign _T_5492 = _T_5490 + _T_5491; // @[Bitwise.scala 48:55:@3433.4]
  assign _T_5493 = _T_5462 + _T_5463; // @[Bitwise.scala 48:55:@3434.4]
  assign _T_5494 = _T_5465 + _T_5466; // @[Bitwise.scala 48:55:@3435.4]
  assign _GEN_665 = {{1'd0}, _T_5464}; // @[Bitwise.scala 48:55:@3436.4]
  assign _T_5495 = _GEN_665 + _T_5494; // @[Bitwise.scala 48:55:@3436.4]
  assign _GEN_666 = {{1'd0}, _T_5493}; // @[Bitwise.scala 48:55:@3437.4]
  assign _T_5496 = _GEN_666 + _T_5495; // @[Bitwise.scala 48:55:@3437.4]
  assign _GEN_667 = {{1'd0}, _T_5492}; // @[Bitwise.scala 48:55:@3438.4]
  assign _T_5497 = _GEN_667 + _T_5496; // @[Bitwise.scala 48:55:@3438.4]
  assign _GEN_668 = {{1'd0}, _T_5489}; // @[Bitwise.scala 48:55:@3439.4]
  assign _T_5498 = _GEN_668 + _T_5497; // @[Bitwise.scala 48:55:@3439.4]
  assign _T_5499 = _T_5482 + _T_5498; // @[Bitwise.scala 48:55:@3440.4]
  assign _T_5563 = _T_2230[34:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3505.4]
  assign _T_5564 = _T_5563[0]; // @[Bitwise.scala 50:65:@3506.4]
  assign _T_5565 = _T_5563[1]; // @[Bitwise.scala 50:65:@3507.4]
  assign _T_5566 = _T_5563[2]; // @[Bitwise.scala 50:65:@3508.4]
  assign _T_5567 = _T_5563[3]; // @[Bitwise.scala 50:65:@3509.4]
  assign _T_5568 = _T_5563[4]; // @[Bitwise.scala 50:65:@3510.4]
  assign _T_5569 = _T_5563[5]; // @[Bitwise.scala 50:65:@3511.4]
  assign _T_5570 = _T_5563[6]; // @[Bitwise.scala 50:65:@3512.4]
  assign _T_5571 = _T_5563[7]; // @[Bitwise.scala 50:65:@3513.4]
  assign _T_5572 = _T_5563[8]; // @[Bitwise.scala 50:65:@3514.4]
  assign _T_5573 = _T_5563[9]; // @[Bitwise.scala 50:65:@3515.4]
  assign _T_5574 = _T_5563[10]; // @[Bitwise.scala 50:65:@3516.4]
  assign _T_5575 = _T_5563[11]; // @[Bitwise.scala 50:65:@3517.4]
  assign _T_5576 = _T_5563[12]; // @[Bitwise.scala 50:65:@3518.4]
  assign _T_5577 = _T_5563[13]; // @[Bitwise.scala 50:65:@3519.4]
  assign _T_5578 = _T_5563[14]; // @[Bitwise.scala 50:65:@3520.4]
  assign _T_5579 = _T_5563[15]; // @[Bitwise.scala 50:65:@3521.4]
  assign _T_5580 = _T_5563[16]; // @[Bitwise.scala 50:65:@3522.4]
  assign _T_5581 = _T_5563[17]; // @[Bitwise.scala 50:65:@3523.4]
  assign _T_5582 = _T_5563[18]; // @[Bitwise.scala 50:65:@3524.4]
  assign _T_5583 = _T_5563[19]; // @[Bitwise.scala 50:65:@3525.4]
  assign _T_5584 = _T_5563[20]; // @[Bitwise.scala 50:65:@3526.4]
  assign _T_5585 = _T_5563[21]; // @[Bitwise.scala 50:65:@3527.4]
  assign _T_5586 = _T_5563[22]; // @[Bitwise.scala 50:65:@3528.4]
  assign _T_5587 = _T_5563[23]; // @[Bitwise.scala 50:65:@3529.4]
  assign _T_5588 = _T_5563[24]; // @[Bitwise.scala 50:65:@3530.4]
  assign _T_5589 = _T_5563[25]; // @[Bitwise.scala 50:65:@3531.4]
  assign _T_5590 = _T_5563[26]; // @[Bitwise.scala 50:65:@3532.4]
  assign _T_5591 = _T_5563[27]; // @[Bitwise.scala 50:65:@3533.4]
  assign _T_5592 = _T_5563[28]; // @[Bitwise.scala 50:65:@3534.4]
  assign _T_5593 = _T_5563[29]; // @[Bitwise.scala 50:65:@3535.4]
  assign _T_5594 = _T_5563[30]; // @[Bitwise.scala 50:65:@3536.4]
  assign _T_5595 = _T_5563[31]; // @[Bitwise.scala 50:65:@3537.4]
  assign _T_5596 = _T_5563[32]; // @[Bitwise.scala 50:65:@3538.4]
  assign _T_5597 = _T_5563[33]; // @[Bitwise.scala 50:65:@3539.4]
  assign _T_5598 = _T_5563[34]; // @[Bitwise.scala 50:65:@3540.4]
  assign _T_5599 = _T_5564 + _T_5565; // @[Bitwise.scala 48:55:@3541.4]
  assign _T_5600 = _T_5566 + _T_5567; // @[Bitwise.scala 48:55:@3542.4]
  assign _T_5601 = _T_5599 + _T_5600; // @[Bitwise.scala 48:55:@3543.4]
  assign _T_5602 = _T_5568 + _T_5569; // @[Bitwise.scala 48:55:@3544.4]
  assign _T_5603 = _T_5570 + _T_5571; // @[Bitwise.scala 48:55:@3545.4]
  assign _T_5604 = _T_5602 + _T_5603; // @[Bitwise.scala 48:55:@3546.4]
  assign _T_5605 = _T_5601 + _T_5604; // @[Bitwise.scala 48:55:@3547.4]
  assign _T_5606 = _T_5572 + _T_5573; // @[Bitwise.scala 48:55:@3548.4]
  assign _T_5607 = _T_5574 + _T_5575; // @[Bitwise.scala 48:55:@3549.4]
  assign _T_5608 = _T_5606 + _T_5607; // @[Bitwise.scala 48:55:@3550.4]
  assign _T_5609 = _T_5576 + _T_5577; // @[Bitwise.scala 48:55:@3551.4]
  assign _T_5610 = _T_5579 + _T_5580; // @[Bitwise.scala 48:55:@3552.4]
  assign _GEN_669 = {{1'd0}, _T_5578}; // @[Bitwise.scala 48:55:@3553.4]
  assign _T_5611 = _GEN_669 + _T_5610; // @[Bitwise.scala 48:55:@3553.4]
  assign _GEN_670 = {{1'd0}, _T_5609}; // @[Bitwise.scala 48:55:@3554.4]
  assign _T_5612 = _GEN_670 + _T_5611; // @[Bitwise.scala 48:55:@3554.4]
  assign _GEN_671 = {{1'd0}, _T_5608}; // @[Bitwise.scala 48:55:@3555.4]
  assign _T_5613 = _GEN_671 + _T_5612; // @[Bitwise.scala 48:55:@3555.4]
  assign _GEN_672 = {{1'd0}, _T_5605}; // @[Bitwise.scala 48:55:@3556.4]
  assign _T_5614 = _GEN_672 + _T_5613; // @[Bitwise.scala 48:55:@3556.4]
  assign _T_5615 = _T_5581 + _T_5582; // @[Bitwise.scala 48:55:@3557.4]
  assign _T_5616 = _T_5583 + _T_5584; // @[Bitwise.scala 48:55:@3558.4]
  assign _T_5617 = _T_5615 + _T_5616; // @[Bitwise.scala 48:55:@3559.4]
  assign _T_5618 = _T_5585 + _T_5586; // @[Bitwise.scala 48:55:@3560.4]
  assign _T_5619 = _T_5588 + _T_5589; // @[Bitwise.scala 48:55:@3561.4]
  assign _GEN_673 = {{1'd0}, _T_5587}; // @[Bitwise.scala 48:55:@3562.4]
  assign _T_5620 = _GEN_673 + _T_5619; // @[Bitwise.scala 48:55:@3562.4]
  assign _GEN_674 = {{1'd0}, _T_5618}; // @[Bitwise.scala 48:55:@3563.4]
  assign _T_5621 = _GEN_674 + _T_5620; // @[Bitwise.scala 48:55:@3563.4]
  assign _GEN_675 = {{1'd0}, _T_5617}; // @[Bitwise.scala 48:55:@3564.4]
  assign _T_5622 = _GEN_675 + _T_5621; // @[Bitwise.scala 48:55:@3564.4]
  assign _T_5623 = _T_5590 + _T_5591; // @[Bitwise.scala 48:55:@3565.4]
  assign _T_5624 = _T_5592 + _T_5593; // @[Bitwise.scala 48:55:@3566.4]
  assign _T_5625 = _T_5623 + _T_5624; // @[Bitwise.scala 48:55:@3567.4]
  assign _T_5626 = _T_5594 + _T_5595; // @[Bitwise.scala 48:55:@3568.4]
  assign _T_5627 = _T_5597 + _T_5598; // @[Bitwise.scala 48:55:@3569.4]
  assign _GEN_676 = {{1'd0}, _T_5596}; // @[Bitwise.scala 48:55:@3570.4]
  assign _T_5628 = _GEN_676 + _T_5627; // @[Bitwise.scala 48:55:@3570.4]
  assign _GEN_677 = {{1'd0}, _T_5626}; // @[Bitwise.scala 48:55:@3571.4]
  assign _T_5629 = _GEN_677 + _T_5628; // @[Bitwise.scala 48:55:@3571.4]
  assign _GEN_678 = {{1'd0}, _T_5625}; // @[Bitwise.scala 48:55:@3572.4]
  assign _T_5630 = _GEN_678 + _T_5629; // @[Bitwise.scala 48:55:@3572.4]
  assign _T_5631 = _T_5622 + _T_5630; // @[Bitwise.scala 48:55:@3573.4]
  assign _T_5632 = _T_5614 + _T_5631; // @[Bitwise.scala 48:55:@3574.4]
  assign _T_5696 = _T_2230[35:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3639.4]
  assign _T_5697 = _T_5696[0]; // @[Bitwise.scala 50:65:@3640.4]
  assign _T_5698 = _T_5696[1]; // @[Bitwise.scala 50:65:@3641.4]
  assign _T_5699 = _T_5696[2]; // @[Bitwise.scala 50:65:@3642.4]
  assign _T_5700 = _T_5696[3]; // @[Bitwise.scala 50:65:@3643.4]
  assign _T_5701 = _T_5696[4]; // @[Bitwise.scala 50:65:@3644.4]
  assign _T_5702 = _T_5696[5]; // @[Bitwise.scala 50:65:@3645.4]
  assign _T_5703 = _T_5696[6]; // @[Bitwise.scala 50:65:@3646.4]
  assign _T_5704 = _T_5696[7]; // @[Bitwise.scala 50:65:@3647.4]
  assign _T_5705 = _T_5696[8]; // @[Bitwise.scala 50:65:@3648.4]
  assign _T_5706 = _T_5696[9]; // @[Bitwise.scala 50:65:@3649.4]
  assign _T_5707 = _T_5696[10]; // @[Bitwise.scala 50:65:@3650.4]
  assign _T_5708 = _T_5696[11]; // @[Bitwise.scala 50:65:@3651.4]
  assign _T_5709 = _T_5696[12]; // @[Bitwise.scala 50:65:@3652.4]
  assign _T_5710 = _T_5696[13]; // @[Bitwise.scala 50:65:@3653.4]
  assign _T_5711 = _T_5696[14]; // @[Bitwise.scala 50:65:@3654.4]
  assign _T_5712 = _T_5696[15]; // @[Bitwise.scala 50:65:@3655.4]
  assign _T_5713 = _T_5696[16]; // @[Bitwise.scala 50:65:@3656.4]
  assign _T_5714 = _T_5696[17]; // @[Bitwise.scala 50:65:@3657.4]
  assign _T_5715 = _T_5696[18]; // @[Bitwise.scala 50:65:@3658.4]
  assign _T_5716 = _T_5696[19]; // @[Bitwise.scala 50:65:@3659.4]
  assign _T_5717 = _T_5696[20]; // @[Bitwise.scala 50:65:@3660.4]
  assign _T_5718 = _T_5696[21]; // @[Bitwise.scala 50:65:@3661.4]
  assign _T_5719 = _T_5696[22]; // @[Bitwise.scala 50:65:@3662.4]
  assign _T_5720 = _T_5696[23]; // @[Bitwise.scala 50:65:@3663.4]
  assign _T_5721 = _T_5696[24]; // @[Bitwise.scala 50:65:@3664.4]
  assign _T_5722 = _T_5696[25]; // @[Bitwise.scala 50:65:@3665.4]
  assign _T_5723 = _T_5696[26]; // @[Bitwise.scala 50:65:@3666.4]
  assign _T_5724 = _T_5696[27]; // @[Bitwise.scala 50:65:@3667.4]
  assign _T_5725 = _T_5696[28]; // @[Bitwise.scala 50:65:@3668.4]
  assign _T_5726 = _T_5696[29]; // @[Bitwise.scala 50:65:@3669.4]
  assign _T_5727 = _T_5696[30]; // @[Bitwise.scala 50:65:@3670.4]
  assign _T_5728 = _T_5696[31]; // @[Bitwise.scala 50:65:@3671.4]
  assign _T_5729 = _T_5696[32]; // @[Bitwise.scala 50:65:@3672.4]
  assign _T_5730 = _T_5696[33]; // @[Bitwise.scala 50:65:@3673.4]
  assign _T_5731 = _T_5696[34]; // @[Bitwise.scala 50:65:@3674.4]
  assign _T_5732 = _T_5696[35]; // @[Bitwise.scala 50:65:@3675.4]
  assign _T_5733 = _T_5697 + _T_5698; // @[Bitwise.scala 48:55:@3676.4]
  assign _T_5734 = _T_5699 + _T_5700; // @[Bitwise.scala 48:55:@3677.4]
  assign _T_5735 = _T_5733 + _T_5734; // @[Bitwise.scala 48:55:@3678.4]
  assign _T_5736 = _T_5701 + _T_5702; // @[Bitwise.scala 48:55:@3679.4]
  assign _T_5737 = _T_5704 + _T_5705; // @[Bitwise.scala 48:55:@3680.4]
  assign _GEN_679 = {{1'd0}, _T_5703}; // @[Bitwise.scala 48:55:@3681.4]
  assign _T_5738 = _GEN_679 + _T_5737; // @[Bitwise.scala 48:55:@3681.4]
  assign _GEN_680 = {{1'd0}, _T_5736}; // @[Bitwise.scala 48:55:@3682.4]
  assign _T_5739 = _GEN_680 + _T_5738; // @[Bitwise.scala 48:55:@3682.4]
  assign _GEN_681 = {{1'd0}, _T_5735}; // @[Bitwise.scala 48:55:@3683.4]
  assign _T_5740 = _GEN_681 + _T_5739; // @[Bitwise.scala 48:55:@3683.4]
  assign _T_5741 = _T_5706 + _T_5707; // @[Bitwise.scala 48:55:@3684.4]
  assign _T_5742 = _T_5708 + _T_5709; // @[Bitwise.scala 48:55:@3685.4]
  assign _T_5743 = _T_5741 + _T_5742; // @[Bitwise.scala 48:55:@3686.4]
  assign _T_5744 = _T_5710 + _T_5711; // @[Bitwise.scala 48:55:@3687.4]
  assign _T_5745 = _T_5713 + _T_5714; // @[Bitwise.scala 48:55:@3688.4]
  assign _GEN_682 = {{1'd0}, _T_5712}; // @[Bitwise.scala 48:55:@3689.4]
  assign _T_5746 = _GEN_682 + _T_5745; // @[Bitwise.scala 48:55:@3689.4]
  assign _GEN_683 = {{1'd0}, _T_5744}; // @[Bitwise.scala 48:55:@3690.4]
  assign _T_5747 = _GEN_683 + _T_5746; // @[Bitwise.scala 48:55:@3690.4]
  assign _GEN_684 = {{1'd0}, _T_5743}; // @[Bitwise.scala 48:55:@3691.4]
  assign _T_5748 = _GEN_684 + _T_5747; // @[Bitwise.scala 48:55:@3691.4]
  assign _T_5749 = _T_5740 + _T_5748; // @[Bitwise.scala 48:55:@3692.4]
  assign _T_5750 = _T_5715 + _T_5716; // @[Bitwise.scala 48:55:@3693.4]
  assign _T_5751 = _T_5717 + _T_5718; // @[Bitwise.scala 48:55:@3694.4]
  assign _T_5752 = _T_5750 + _T_5751; // @[Bitwise.scala 48:55:@3695.4]
  assign _T_5753 = _T_5719 + _T_5720; // @[Bitwise.scala 48:55:@3696.4]
  assign _T_5754 = _T_5722 + _T_5723; // @[Bitwise.scala 48:55:@3697.4]
  assign _GEN_685 = {{1'd0}, _T_5721}; // @[Bitwise.scala 48:55:@3698.4]
  assign _T_5755 = _GEN_685 + _T_5754; // @[Bitwise.scala 48:55:@3698.4]
  assign _GEN_686 = {{1'd0}, _T_5753}; // @[Bitwise.scala 48:55:@3699.4]
  assign _T_5756 = _GEN_686 + _T_5755; // @[Bitwise.scala 48:55:@3699.4]
  assign _GEN_687 = {{1'd0}, _T_5752}; // @[Bitwise.scala 48:55:@3700.4]
  assign _T_5757 = _GEN_687 + _T_5756; // @[Bitwise.scala 48:55:@3700.4]
  assign _T_5758 = _T_5724 + _T_5725; // @[Bitwise.scala 48:55:@3701.4]
  assign _T_5759 = _T_5726 + _T_5727; // @[Bitwise.scala 48:55:@3702.4]
  assign _T_5760 = _T_5758 + _T_5759; // @[Bitwise.scala 48:55:@3703.4]
  assign _T_5761 = _T_5728 + _T_5729; // @[Bitwise.scala 48:55:@3704.4]
  assign _T_5762 = _T_5731 + _T_5732; // @[Bitwise.scala 48:55:@3705.4]
  assign _GEN_688 = {{1'd0}, _T_5730}; // @[Bitwise.scala 48:55:@3706.4]
  assign _T_5763 = _GEN_688 + _T_5762; // @[Bitwise.scala 48:55:@3706.4]
  assign _GEN_689 = {{1'd0}, _T_5761}; // @[Bitwise.scala 48:55:@3707.4]
  assign _T_5764 = _GEN_689 + _T_5763; // @[Bitwise.scala 48:55:@3707.4]
  assign _GEN_690 = {{1'd0}, _T_5760}; // @[Bitwise.scala 48:55:@3708.4]
  assign _T_5765 = _GEN_690 + _T_5764; // @[Bitwise.scala 48:55:@3708.4]
  assign _T_5766 = _T_5757 + _T_5765; // @[Bitwise.scala 48:55:@3709.4]
  assign _T_5767 = _T_5749 + _T_5766; // @[Bitwise.scala 48:55:@3710.4]
  assign _T_5831 = _T_2230[36:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3775.4]
  assign _T_5832 = _T_5831[0]; // @[Bitwise.scala 50:65:@3776.4]
  assign _T_5833 = _T_5831[1]; // @[Bitwise.scala 50:65:@3777.4]
  assign _T_5834 = _T_5831[2]; // @[Bitwise.scala 50:65:@3778.4]
  assign _T_5835 = _T_5831[3]; // @[Bitwise.scala 50:65:@3779.4]
  assign _T_5836 = _T_5831[4]; // @[Bitwise.scala 50:65:@3780.4]
  assign _T_5837 = _T_5831[5]; // @[Bitwise.scala 50:65:@3781.4]
  assign _T_5838 = _T_5831[6]; // @[Bitwise.scala 50:65:@3782.4]
  assign _T_5839 = _T_5831[7]; // @[Bitwise.scala 50:65:@3783.4]
  assign _T_5840 = _T_5831[8]; // @[Bitwise.scala 50:65:@3784.4]
  assign _T_5841 = _T_5831[9]; // @[Bitwise.scala 50:65:@3785.4]
  assign _T_5842 = _T_5831[10]; // @[Bitwise.scala 50:65:@3786.4]
  assign _T_5843 = _T_5831[11]; // @[Bitwise.scala 50:65:@3787.4]
  assign _T_5844 = _T_5831[12]; // @[Bitwise.scala 50:65:@3788.4]
  assign _T_5845 = _T_5831[13]; // @[Bitwise.scala 50:65:@3789.4]
  assign _T_5846 = _T_5831[14]; // @[Bitwise.scala 50:65:@3790.4]
  assign _T_5847 = _T_5831[15]; // @[Bitwise.scala 50:65:@3791.4]
  assign _T_5848 = _T_5831[16]; // @[Bitwise.scala 50:65:@3792.4]
  assign _T_5849 = _T_5831[17]; // @[Bitwise.scala 50:65:@3793.4]
  assign _T_5850 = _T_5831[18]; // @[Bitwise.scala 50:65:@3794.4]
  assign _T_5851 = _T_5831[19]; // @[Bitwise.scala 50:65:@3795.4]
  assign _T_5852 = _T_5831[20]; // @[Bitwise.scala 50:65:@3796.4]
  assign _T_5853 = _T_5831[21]; // @[Bitwise.scala 50:65:@3797.4]
  assign _T_5854 = _T_5831[22]; // @[Bitwise.scala 50:65:@3798.4]
  assign _T_5855 = _T_5831[23]; // @[Bitwise.scala 50:65:@3799.4]
  assign _T_5856 = _T_5831[24]; // @[Bitwise.scala 50:65:@3800.4]
  assign _T_5857 = _T_5831[25]; // @[Bitwise.scala 50:65:@3801.4]
  assign _T_5858 = _T_5831[26]; // @[Bitwise.scala 50:65:@3802.4]
  assign _T_5859 = _T_5831[27]; // @[Bitwise.scala 50:65:@3803.4]
  assign _T_5860 = _T_5831[28]; // @[Bitwise.scala 50:65:@3804.4]
  assign _T_5861 = _T_5831[29]; // @[Bitwise.scala 50:65:@3805.4]
  assign _T_5862 = _T_5831[30]; // @[Bitwise.scala 50:65:@3806.4]
  assign _T_5863 = _T_5831[31]; // @[Bitwise.scala 50:65:@3807.4]
  assign _T_5864 = _T_5831[32]; // @[Bitwise.scala 50:65:@3808.4]
  assign _T_5865 = _T_5831[33]; // @[Bitwise.scala 50:65:@3809.4]
  assign _T_5866 = _T_5831[34]; // @[Bitwise.scala 50:65:@3810.4]
  assign _T_5867 = _T_5831[35]; // @[Bitwise.scala 50:65:@3811.4]
  assign _T_5868 = _T_5831[36]; // @[Bitwise.scala 50:65:@3812.4]
  assign _T_5869 = _T_5832 + _T_5833; // @[Bitwise.scala 48:55:@3813.4]
  assign _T_5870 = _T_5834 + _T_5835; // @[Bitwise.scala 48:55:@3814.4]
  assign _T_5871 = _T_5869 + _T_5870; // @[Bitwise.scala 48:55:@3815.4]
  assign _T_5872 = _T_5836 + _T_5837; // @[Bitwise.scala 48:55:@3816.4]
  assign _T_5873 = _T_5839 + _T_5840; // @[Bitwise.scala 48:55:@3817.4]
  assign _GEN_691 = {{1'd0}, _T_5838}; // @[Bitwise.scala 48:55:@3818.4]
  assign _T_5874 = _GEN_691 + _T_5873; // @[Bitwise.scala 48:55:@3818.4]
  assign _GEN_692 = {{1'd0}, _T_5872}; // @[Bitwise.scala 48:55:@3819.4]
  assign _T_5875 = _GEN_692 + _T_5874; // @[Bitwise.scala 48:55:@3819.4]
  assign _GEN_693 = {{1'd0}, _T_5871}; // @[Bitwise.scala 48:55:@3820.4]
  assign _T_5876 = _GEN_693 + _T_5875; // @[Bitwise.scala 48:55:@3820.4]
  assign _T_5877 = _T_5841 + _T_5842; // @[Bitwise.scala 48:55:@3821.4]
  assign _T_5878 = _T_5843 + _T_5844; // @[Bitwise.scala 48:55:@3822.4]
  assign _T_5879 = _T_5877 + _T_5878; // @[Bitwise.scala 48:55:@3823.4]
  assign _T_5880 = _T_5845 + _T_5846; // @[Bitwise.scala 48:55:@3824.4]
  assign _T_5881 = _T_5848 + _T_5849; // @[Bitwise.scala 48:55:@3825.4]
  assign _GEN_694 = {{1'd0}, _T_5847}; // @[Bitwise.scala 48:55:@3826.4]
  assign _T_5882 = _GEN_694 + _T_5881; // @[Bitwise.scala 48:55:@3826.4]
  assign _GEN_695 = {{1'd0}, _T_5880}; // @[Bitwise.scala 48:55:@3827.4]
  assign _T_5883 = _GEN_695 + _T_5882; // @[Bitwise.scala 48:55:@3827.4]
  assign _GEN_696 = {{1'd0}, _T_5879}; // @[Bitwise.scala 48:55:@3828.4]
  assign _T_5884 = _GEN_696 + _T_5883; // @[Bitwise.scala 48:55:@3828.4]
  assign _T_5885 = _T_5876 + _T_5884; // @[Bitwise.scala 48:55:@3829.4]
  assign _T_5886 = _T_5850 + _T_5851; // @[Bitwise.scala 48:55:@3830.4]
  assign _T_5887 = _T_5852 + _T_5853; // @[Bitwise.scala 48:55:@3831.4]
  assign _T_5888 = _T_5886 + _T_5887; // @[Bitwise.scala 48:55:@3832.4]
  assign _T_5889 = _T_5854 + _T_5855; // @[Bitwise.scala 48:55:@3833.4]
  assign _T_5890 = _T_5857 + _T_5858; // @[Bitwise.scala 48:55:@3834.4]
  assign _GEN_697 = {{1'd0}, _T_5856}; // @[Bitwise.scala 48:55:@3835.4]
  assign _T_5891 = _GEN_697 + _T_5890; // @[Bitwise.scala 48:55:@3835.4]
  assign _GEN_698 = {{1'd0}, _T_5889}; // @[Bitwise.scala 48:55:@3836.4]
  assign _T_5892 = _GEN_698 + _T_5891; // @[Bitwise.scala 48:55:@3836.4]
  assign _GEN_699 = {{1'd0}, _T_5888}; // @[Bitwise.scala 48:55:@3837.4]
  assign _T_5893 = _GEN_699 + _T_5892; // @[Bitwise.scala 48:55:@3837.4]
  assign _T_5894 = _T_5859 + _T_5860; // @[Bitwise.scala 48:55:@3838.4]
  assign _T_5895 = _T_5862 + _T_5863; // @[Bitwise.scala 48:55:@3839.4]
  assign _GEN_700 = {{1'd0}, _T_5861}; // @[Bitwise.scala 48:55:@3840.4]
  assign _T_5896 = _GEN_700 + _T_5895; // @[Bitwise.scala 48:55:@3840.4]
  assign _GEN_701 = {{1'd0}, _T_5894}; // @[Bitwise.scala 48:55:@3841.4]
  assign _T_5897 = _GEN_701 + _T_5896; // @[Bitwise.scala 48:55:@3841.4]
  assign _T_5898 = _T_5864 + _T_5865; // @[Bitwise.scala 48:55:@3842.4]
  assign _T_5899 = _T_5867 + _T_5868; // @[Bitwise.scala 48:55:@3843.4]
  assign _GEN_702 = {{1'd0}, _T_5866}; // @[Bitwise.scala 48:55:@3844.4]
  assign _T_5900 = _GEN_702 + _T_5899; // @[Bitwise.scala 48:55:@3844.4]
  assign _GEN_703 = {{1'd0}, _T_5898}; // @[Bitwise.scala 48:55:@3845.4]
  assign _T_5901 = _GEN_703 + _T_5900; // @[Bitwise.scala 48:55:@3845.4]
  assign _T_5902 = _T_5897 + _T_5901; // @[Bitwise.scala 48:55:@3846.4]
  assign _T_5903 = _T_5893 + _T_5902; // @[Bitwise.scala 48:55:@3847.4]
  assign _T_5904 = _T_5885 + _T_5903; // @[Bitwise.scala 48:55:@3848.4]
  assign _T_5968 = _T_2230[37:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@3913.4]
  assign _T_5969 = _T_5968[0]; // @[Bitwise.scala 50:65:@3914.4]
  assign _T_5970 = _T_5968[1]; // @[Bitwise.scala 50:65:@3915.4]
  assign _T_5971 = _T_5968[2]; // @[Bitwise.scala 50:65:@3916.4]
  assign _T_5972 = _T_5968[3]; // @[Bitwise.scala 50:65:@3917.4]
  assign _T_5973 = _T_5968[4]; // @[Bitwise.scala 50:65:@3918.4]
  assign _T_5974 = _T_5968[5]; // @[Bitwise.scala 50:65:@3919.4]
  assign _T_5975 = _T_5968[6]; // @[Bitwise.scala 50:65:@3920.4]
  assign _T_5976 = _T_5968[7]; // @[Bitwise.scala 50:65:@3921.4]
  assign _T_5977 = _T_5968[8]; // @[Bitwise.scala 50:65:@3922.4]
  assign _T_5978 = _T_5968[9]; // @[Bitwise.scala 50:65:@3923.4]
  assign _T_5979 = _T_5968[10]; // @[Bitwise.scala 50:65:@3924.4]
  assign _T_5980 = _T_5968[11]; // @[Bitwise.scala 50:65:@3925.4]
  assign _T_5981 = _T_5968[12]; // @[Bitwise.scala 50:65:@3926.4]
  assign _T_5982 = _T_5968[13]; // @[Bitwise.scala 50:65:@3927.4]
  assign _T_5983 = _T_5968[14]; // @[Bitwise.scala 50:65:@3928.4]
  assign _T_5984 = _T_5968[15]; // @[Bitwise.scala 50:65:@3929.4]
  assign _T_5985 = _T_5968[16]; // @[Bitwise.scala 50:65:@3930.4]
  assign _T_5986 = _T_5968[17]; // @[Bitwise.scala 50:65:@3931.4]
  assign _T_5987 = _T_5968[18]; // @[Bitwise.scala 50:65:@3932.4]
  assign _T_5988 = _T_5968[19]; // @[Bitwise.scala 50:65:@3933.4]
  assign _T_5989 = _T_5968[20]; // @[Bitwise.scala 50:65:@3934.4]
  assign _T_5990 = _T_5968[21]; // @[Bitwise.scala 50:65:@3935.4]
  assign _T_5991 = _T_5968[22]; // @[Bitwise.scala 50:65:@3936.4]
  assign _T_5992 = _T_5968[23]; // @[Bitwise.scala 50:65:@3937.4]
  assign _T_5993 = _T_5968[24]; // @[Bitwise.scala 50:65:@3938.4]
  assign _T_5994 = _T_5968[25]; // @[Bitwise.scala 50:65:@3939.4]
  assign _T_5995 = _T_5968[26]; // @[Bitwise.scala 50:65:@3940.4]
  assign _T_5996 = _T_5968[27]; // @[Bitwise.scala 50:65:@3941.4]
  assign _T_5997 = _T_5968[28]; // @[Bitwise.scala 50:65:@3942.4]
  assign _T_5998 = _T_5968[29]; // @[Bitwise.scala 50:65:@3943.4]
  assign _T_5999 = _T_5968[30]; // @[Bitwise.scala 50:65:@3944.4]
  assign _T_6000 = _T_5968[31]; // @[Bitwise.scala 50:65:@3945.4]
  assign _T_6001 = _T_5968[32]; // @[Bitwise.scala 50:65:@3946.4]
  assign _T_6002 = _T_5968[33]; // @[Bitwise.scala 50:65:@3947.4]
  assign _T_6003 = _T_5968[34]; // @[Bitwise.scala 50:65:@3948.4]
  assign _T_6004 = _T_5968[35]; // @[Bitwise.scala 50:65:@3949.4]
  assign _T_6005 = _T_5968[36]; // @[Bitwise.scala 50:65:@3950.4]
  assign _T_6006 = _T_5968[37]; // @[Bitwise.scala 50:65:@3951.4]
  assign _T_6007 = _T_5969 + _T_5970; // @[Bitwise.scala 48:55:@3952.4]
  assign _T_6008 = _T_5971 + _T_5972; // @[Bitwise.scala 48:55:@3953.4]
  assign _T_6009 = _T_6007 + _T_6008; // @[Bitwise.scala 48:55:@3954.4]
  assign _T_6010 = _T_5973 + _T_5974; // @[Bitwise.scala 48:55:@3955.4]
  assign _T_6011 = _T_5976 + _T_5977; // @[Bitwise.scala 48:55:@3956.4]
  assign _GEN_704 = {{1'd0}, _T_5975}; // @[Bitwise.scala 48:55:@3957.4]
  assign _T_6012 = _GEN_704 + _T_6011; // @[Bitwise.scala 48:55:@3957.4]
  assign _GEN_705 = {{1'd0}, _T_6010}; // @[Bitwise.scala 48:55:@3958.4]
  assign _T_6013 = _GEN_705 + _T_6012; // @[Bitwise.scala 48:55:@3958.4]
  assign _GEN_706 = {{1'd0}, _T_6009}; // @[Bitwise.scala 48:55:@3959.4]
  assign _T_6014 = _GEN_706 + _T_6013; // @[Bitwise.scala 48:55:@3959.4]
  assign _T_6015 = _T_5978 + _T_5979; // @[Bitwise.scala 48:55:@3960.4]
  assign _T_6016 = _T_5981 + _T_5982; // @[Bitwise.scala 48:55:@3961.4]
  assign _GEN_707 = {{1'd0}, _T_5980}; // @[Bitwise.scala 48:55:@3962.4]
  assign _T_6017 = _GEN_707 + _T_6016; // @[Bitwise.scala 48:55:@3962.4]
  assign _GEN_708 = {{1'd0}, _T_6015}; // @[Bitwise.scala 48:55:@3963.4]
  assign _T_6018 = _GEN_708 + _T_6017; // @[Bitwise.scala 48:55:@3963.4]
  assign _T_6019 = _T_5983 + _T_5984; // @[Bitwise.scala 48:55:@3964.4]
  assign _T_6020 = _T_5986 + _T_5987; // @[Bitwise.scala 48:55:@3965.4]
  assign _GEN_709 = {{1'd0}, _T_5985}; // @[Bitwise.scala 48:55:@3966.4]
  assign _T_6021 = _GEN_709 + _T_6020; // @[Bitwise.scala 48:55:@3966.4]
  assign _GEN_710 = {{1'd0}, _T_6019}; // @[Bitwise.scala 48:55:@3967.4]
  assign _T_6022 = _GEN_710 + _T_6021; // @[Bitwise.scala 48:55:@3967.4]
  assign _T_6023 = _T_6018 + _T_6022; // @[Bitwise.scala 48:55:@3968.4]
  assign _T_6024 = _T_6014 + _T_6023; // @[Bitwise.scala 48:55:@3969.4]
  assign _T_6025 = _T_5988 + _T_5989; // @[Bitwise.scala 48:55:@3970.4]
  assign _T_6026 = _T_5990 + _T_5991; // @[Bitwise.scala 48:55:@3971.4]
  assign _T_6027 = _T_6025 + _T_6026; // @[Bitwise.scala 48:55:@3972.4]
  assign _T_6028 = _T_5992 + _T_5993; // @[Bitwise.scala 48:55:@3973.4]
  assign _T_6029 = _T_5995 + _T_5996; // @[Bitwise.scala 48:55:@3974.4]
  assign _GEN_711 = {{1'd0}, _T_5994}; // @[Bitwise.scala 48:55:@3975.4]
  assign _T_6030 = _GEN_711 + _T_6029; // @[Bitwise.scala 48:55:@3975.4]
  assign _GEN_712 = {{1'd0}, _T_6028}; // @[Bitwise.scala 48:55:@3976.4]
  assign _T_6031 = _GEN_712 + _T_6030; // @[Bitwise.scala 48:55:@3976.4]
  assign _GEN_713 = {{1'd0}, _T_6027}; // @[Bitwise.scala 48:55:@3977.4]
  assign _T_6032 = _GEN_713 + _T_6031; // @[Bitwise.scala 48:55:@3977.4]
  assign _T_6033 = _T_5997 + _T_5998; // @[Bitwise.scala 48:55:@3978.4]
  assign _T_6034 = _T_6000 + _T_6001; // @[Bitwise.scala 48:55:@3979.4]
  assign _GEN_714 = {{1'd0}, _T_5999}; // @[Bitwise.scala 48:55:@3980.4]
  assign _T_6035 = _GEN_714 + _T_6034; // @[Bitwise.scala 48:55:@3980.4]
  assign _GEN_715 = {{1'd0}, _T_6033}; // @[Bitwise.scala 48:55:@3981.4]
  assign _T_6036 = _GEN_715 + _T_6035; // @[Bitwise.scala 48:55:@3981.4]
  assign _T_6037 = _T_6002 + _T_6003; // @[Bitwise.scala 48:55:@3982.4]
  assign _T_6038 = _T_6005 + _T_6006; // @[Bitwise.scala 48:55:@3983.4]
  assign _GEN_716 = {{1'd0}, _T_6004}; // @[Bitwise.scala 48:55:@3984.4]
  assign _T_6039 = _GEN_716 + _T_6038; // @[Bitwise.scala 48:55:@3984.4]
  assign _GEN_717 = {{1'd0}, _T_6037}; // @[Bitwise.scala 48:55:@3985.4]
  assign _T_6040 = _GEN_717 + _T_6039; // @[Bitwise.scala 48:55:@3985.4]
  assign _T_6041 = _T_6036 + _T_6040; // @[Bitwise.scala 48:55:@3986.4]
  assign _T_6042 = _T_6032 + _T_6041; // @[Bitwise.scala 48:55:@3987.4]
  assign _T_6043 = _T_6024 + _T_6042; // @[Bitwise.scala 48:55:@3988.4]
  assign _T_6107 = _T_2230[38:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4053.4]
  assign _T_6108 = _T_6107[0]; // @[Bitwise.scala 50:65:@4054.4]
  assign _T_6109 = _T_6107[1]; // @[Bitwise.scala 50:65:@4055.4]
  assign _T_6110 = _T_6107[2]; // @[Bitwise.scala 50:65:@4056.4]
  assign _T_6111 = _T_6107[3]; // @[Bitwise.scala 50:65:@4057.4]
  assign _T_6112 = _T_6107[4]; // @[Bitwise.scala 50:65:@4058.4]
  assign _T_6113 = _T_6107[5]; // @[Bitwise.scala 50:65:@4059.4]
  assign _T_6114 = _T_6107[6]; // @[Bitwise.scala 50:65:@4060.4]
  assign _T_6115 = _T_6107[7]; // @[Bitwise.scala 50:65:@4061.4]
  assign _T_6116 = _T_6107[8]; // @[Bitwise.scala 50:65:@4062.4]
  assign _T_6117 = _T_6107[9]; // @[Bitwise.scala 50:65:@4063.4]
  assign _T_6118 = _T_6107[10]; // @[Bitwise.scala 50:65:@4064.4]
  assign _T_6119 = _T_6107[11]; // @[Bitwise.scala 50:65:@4065.4]
  assign _T_6120 = _T_6107[12]; // @[Bitwise.scala 50:65:@4066.4]
  assign _T_6121 = _T_6107[13]; // @[Bitwise.scala 50:65:@4067.4]
  assign _T_6122 = _T_6107[14]; // @[Bitwise.scala 50:65:@4068.4]
  assign _T_6123 = _T_6107[15]; // @[Bitwise.scala 50:65:@4069.4]
  assign _T_6124 = _T_6107[16]; // @[Bitwise.scala 50:65:@4070.4]
  assign _T_6125 = _T_6107[17]; // @[Bitwise.scala 50:65:@4071.4]
  assign _T_6126 = _T_6107[18]; // @[Bitwise.scala 50:65:@4072.4]
  assign _T_6127 = _T_6107[19]; // @[Bitwise.scala 50:65:@4073.4]
  assign _T_6128 = _T_6107[20]; // @[Bitwise.scala 50:65:@4074.4]
  assign _T_6129 = _T_6107[21]; // @[Bitwise.scala 50:65:@4075.4]
  assign _T_6130 = _T_6107[22]; // @[Bitwise.scala 50:65:@4076.4]
  assign _T_6131 = _T_6107[23]; // @[Bitwise.scala 50:65:@4077.4]
  assign _T_6132 = _T_6107[24]; // @[Bitwise.scala 50:65:@4078.4]
  assign _T_6133 = _T_6107[25]; // @[Bitwise.scala 50:65:@4079.4]
  assign _T_6134 = _T_6107[26]; // @[Bitwise.scala 50:65:@4080.4]
  assign _T_6135 = _T_6107[27]; // @[Bitwise.scala 50:65:@4081.4]
  assign _T_6136 = _T_6107[28]; // @[Bitwise.scala 50:65:@4082.4]
  assign _T_6137 = _T_6107[29]; // @[Bitwise.scala 50:65:@4083.4]
  assign _T_6138 = _T_6107[30]; // @[Bitwise.scala 50:65:@4084.4]
  assign _T_6139 = _T_6107[31]; // @[Bitwise.scala 50:65:@4085.4]
  assign _T_6140 = _T_6107[32]; // @[Bitwise.scala 50:65:@4086.4]
  assign _T_6141 = _T_6107[33]; // @[Bitwise.scala 50:65:@4087.4]
  assign _T_6142 = _T_6107[34]; // @[Bitwise.scala 50:65:@4088.4]
  assign _T_6143 = _T_6107[35]; // @[Bitwise.scala 50:65:@4089.4]
  assign _T_6144 = _T_6107[36]; // @[Bitwise.scala 50:65:@4090.4]
  assign _T_6145 = _T_6107[37]; // @[Bitwise.scala 50:65:@4091.4]
  assign _T_6146 = _T_6107[38]; // @[Bitwise.scala 50:65:@4092.4]
  assign _T_6147 = _T_6108 + _T_6109; // @[Bitwise.scala 48:55:@4093.4]
  assign _T_6148 = _T_6110 + _T_6111; // @[Bitwise.scala 48:55:@4094.4]
  assign _T_6149 = _T_6147 + _T_6148; // @[Bitwise.scala 48:55:@4095.4]
  assign _T_6150 = _T_6112 + _T_6113; // @[Bitwise.scala 48:55:@4096.4]
  assign _T_6151 = _T_6115 + _T_6116; // @[Bitwise.scala 48:55:@4097.4]
  assign _GEN_718 = {{1'd0}, _T_6114}; // @[Bitwise.scala 48:55:@4098.4]
  assign _T_6152 = _GEN_718 + _T_6151; // @[Bitwise.scala 48:55:@4098.4]
  assign _GEN_719 = {{1'd0}, _T_6150}; // @[Bitwise.scala 48:55:@4099.4]
  assign _T_6153 = _GEN_719 + _T_6152; // @[Bitwise.scala 48:55:@4099.4]
  assign _GEN_720 = {{1'd0}, _T_6149}; // @[Bitwise.scala 48:55:@4100.4]
  assign _T_6154 = _GEN_720 + _T_6153; // @[Bitwise.scala 48:55:@4100.4]
  assign _T_6155 = _T_6117 + _T_6118; // @[Bitwise.scala 48:55:@4101.4]
  assign _T_6156 = _T_6120 + _T_6121; // @[Bitwise.scala 48:55:@4102.4]
  assign _GEN_721 = {{1'd0}, _T_6119}; // @[Bitwise.scala 48:55:@4103.4]
  assign _T_6157 = _GEN_721 + _T_6156; // @[Bitwise.scala 48:55:@4103.4]
  assign _GEN_722 = {{1'd0}, _T_6155}; // @[Bitwise.scala 48:55:@4104.4]
  assign _T_6158 = _GEN_722 + _T_6157; // @[Bitwise.scala 48:55:@4104.4]
  assign _T_6159 = _T_6122 + _T_6123; // @[Bitwise.scala 48:55:@4105.4]
  assign _T_6160 = _T_6125 + _T_6126; // @[Bitwise.scala 48:55:@4106.4]
  assign _GEN_723 = {{1'd0}, _T_6124}; // @[Bitwise.scala 48:55:@4107.4]
  assign _T_6161 = _GEN_723 + _T_6160; // @[Bitwise.scala 48:55:@4107.4]
  assign _GEN_724 = {{1'd0}, _T_6159}; // @[Bitwise.scala 48:55:@4108.4]
  assign _T_6162 = _GEN_724 + _T_6161; // @[Bitwise.scala 48:55:@4108.4]
  assign _T_6163 = _T_6158 + _T_6162; // @[Bitwise.scala 48:55:@4109.4]
  assign _T_6164 = _T_6154 + _T_6163; // @[Bitwise.scala 48:55:@4110.4]
  assign _T_6165 = _T_6127 + _T_6128; // @[Bitwise.scala 48:55:@4111.4]
  assign _T_6166 = _T_6130 + _T_6131; // @[Bitwise.scala 48:55:@4112.4]
  assign _GEN_725 = {{1'd0}, _T_6129}; // @[Bitwise.scala 48:55:@4113.4]
  assign _T_6167 = _GEN_725 + _T_6166; // @[Bitwise.scala 48:55:@4113.4]
  assign _GEN_726 = {{1'd0}, _T_6165}; // @[Bitwise.scala 48:55:@4114.4]
  assign _T_6168 = _GEN_726 + _T_6167; // @[Bitwise.scala 48:55:@4114.4]
  assign _T_6169 = _T_6132 + _T_6133; // @[Bitwise.scala 48:55:@4115.4]
  assign _T_6170 = _T_6135 + _T_6136; // @[Bitwise.scala 48:55:@4116.4]
  assign _GEN_727 = {{1'd0}, _T_6134}; // @[Bitwise.scala 48:55:@4117.4]
  assign _T_6171 = _GEN_727 + _T_6170; // @[Bitwise.scala 48:55:@4117.4]
  assign _GEN_728 = {{1'd0}, _T_6169}; // @[Bitwise.scala 48:55:@4118.4]
  assign _T_6172 = _GEN_728 + _T_6171; // @[Bitwise.scala 48:55:@4118.4]
  assign _T_6173 = _T_6168 + _T_6172; // @[Bitwise.scala 48:55:@4119.4]
  assign _T_6174 = _T_6137 + _T_6138; // @[Bitwise.scala 48:55:@4120.4]
  assign _T_6175 = _T_6140 + _T_6141; // @[Bitwise.scala 48:55:@4121.4]
  assign _GEN_729 = {{1'd0}, _T_6139}; // @[Bitwise.scala 48:55:@4122.4]
  assign _T_6176 = _GEN_729 + _T_6175; // @[Bitwise.scala 48:55:@4122.4]
  assign _GEN_730 = {{1'd0}, _T_6174}; // @[Bitwise.scala 48:55:@4123.4]
  assign _T_6177 = _GEN_730 + _T_6176; // @[Bitwise.scala 48:55:@4123.4]
  assign _T_6178 = _T_6142 + _T_6143; // @[Bitwise.scala 48:55:@4124.4]
  assign _T_6179 = _T_6145 + _T_6146; // @[Bitwise.scala 48:55:@4125.4]
  assign _GEN_731 = {{1'd0}, _T_6144}; // @[Bitwise.scala 48:55:@4126.4]
  assign _T_6180 = _GEN_731 + _T_6179; // @[Bitwise.scala 48:55:@4126.4]
  assign _GEN_732 = {{1'd0}, _T_6178}; // @[Bitwise.scala 48:55:@4127.4]
  assign _T_6181 = _GEN_732 + _T_6180; // @[Bitwise.scala 48:55:@4127.4]
  assign _T_6182 = _T_6177 + _T_6181; // @[Bitwise.scala 48:55:@4128.4]
  assign _T_6183 = _T_6173 + _T_6182; // @[Bitwise.scala 48:55:@4129.4]
  assign _T_6184 = _T_6164 + _T_6183; // @[Bitwise.scala 48:55:@4130.4]
  assign _T_6248 = _T_2230[39:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4195.4]
  assign _T_6249 = _T_6248[0]; // @[Bitwise.scala 50:65:@4196.4]
  assign _T_6250 = _T_6248[1]; // @[Bitwise.scala 50:65:@4197.4]
  assign _T_6251 = _T_6248[2]; // @[Bitwise.scala 50:65:@4198.4]
  assign _T_6252 = _T_6248[3]; // @[Bitwise.scala 50:65:@4199.4]
  assign _T_6253 = _T_6248[4]; // @[Bitwise.scala 50:65:@4200.4]
  assign _T_6254 = _T_6248[5]; // @[Bitwise.scala 50:65:@4201.4]
  assign _T_6255 = _T_6248[6]; // @[Bitwise.scala 50:65:@4202.4]
  assign _T_6256 = _T_6248[7]; // @[Bitwise.scala 50:65:@4203.4]
  assign _T_6257 = _T_6248[8]; // @[Bitwise.scala 50:65:@4204.4]
  assign _T_6258 = _T_6248[9]; // @[Bitwise.scala 50:65:@4205.4]
  assign _T_6259 = _T_6248[10]; // @[Bitwise.scala 50:65:@4206.4]
  assign _T_6260 = _T_6248[11]; // @[Bitwise.scala 50:65:@4207.4]
  assign _T_6261 = _T_6248[12]; // @[Bitwise.scala 50:65:@4208.4]
  assign _T_6262 = _T_6248[13]; // @[Bitwise.scala 50:65:@4209.4]
  assign _T_6263 = _T_6248[14]; // @[Bitwise.scala 50:65:@4210.4]
  assign _T_6264 = _T_6248[15]; // @[Bitwise.scala 50:65:@4211.4]
  assign _T_6265 = _T_6248[16]; // @[Bitwise.scala 50:65:@4212.4]
  assign _T_6266 = _T_6248[17]; // @[Bitwise.scala 50:65:@4213.4]
  assign _T_6267 = _T_6248[18]; // @[Bitwise.scala 50:65:@4214.4]
  assign _T_6268 = _T_6248[19]; // @[Bitwise.scala 50:65:@4215.4]
  assign _T_6269 = _T_6248[20]; // @[Bitwise.scala 50:65:@4216.4]
  assign _T_6270 = _T_6248[21]; // @[Bitwise.scala 50:65:@4217.4]
  assign _T_6271 = _T_6248[22]; // @[Bitwise.scala 50:65:@4218.4]
  assign _T_6272 = _T_6248[23]; // @[Bitwise.scala 50:65:@4219.4]
  assign _T_6273 = _T_6248[24]; // @[Bitwise.scala 50:65:@4220.4]
  assign _T_6274 = _T_6248[25]; // @[Bitwise.scala 50:65:@4221.4]
  assign _T_6275 = _T_6248[26]; // @[Bitwise.scala 50:65:@4222.4]
  assign _T_6276 = _T_6248[27]; // @[Bitwise.scala 50:65:@4223.4]
  assign _T_6277 = _T_6248[28]; // @[Bitwise.scala 50:65:@4224.4]
  assign _T_6278 = _T_6248[29]; // @[Bitwise.scala 50:65:@4225.4]
  assign _T_6279 = _T_6248[30]; // @[Bitwise.scala 50:65:@4226.4]
  assign _T_6280 = _T_6248[31]; // @[Bitwise.scala 50:65:@4227.4]
  assign _T_6281 = _T_6248[32]; // @[Bitwise.scala 50:65:@4228.4]
  assign _T_6282 = _T_6248[33]; // @[Bitwise.scala 50:65:@4229.4]
  assign _T_6283 = _T_6248[34]; // @[Bitwise.scala 50:65:@4230.4]
  assign _T_6284 = _T_6248[35]; // @[Bitwise.scala 50:65:@4231.4]
  assign _T_6285 = _T_6248[36]; // @[Bitwise.scala 50:65:@4232.4]
  assign _T_6286 = _T_6248[37]; // @[Bitwise.scala 50:65:@4233.4]
  assign _T_6287 = _T_6248[38]; // @[Bitwise.scala 50:65:@4234.4]
  assign _T_6288 = _T_6248[39]; // @[Bitwise.scala 50:65:@4235.4]
  assign _T_6289 = _T_6249 + _T_6250; // @[Bitwise.scala 48:55:@4236.4]
  assign _T_6290 = _T_6252 + _T_6253; // @[Bitwise.scala 48:55:@4237.4]
  assign _GEN_733 = {{1'd0}, _T_6251}; // @[Bitwise.scala 48:55:@4238.4]
  assign _T_6291 = _GEN_733 + _T_6290; // @[Bitwise.scala 48:55:@4238.4]
  assign _GEN_734 = {{1'd0}, _T_6289}; // @[Bitwise.scala 48:55:@4239.4]
  assign _T_6292 = _GEN_734 + _T_6291; // @[Bitwise.scala 48:55:@4239.4]
  assign _T_6293 = _T_6254 + _T_6255; // @[Bitwise.scala 48:55:@4240.4]
  assign _T_6294 = _T_6257 + _T_6258; // @[Bitwise.scala 48:55:@4241.4]
  assign _GEN_735 = {{1'd0}, _T_6256}; // @[Bitwise.scala 48:55:@4242.4]
  assign _T_6295 = _GEN_735 + _T_6294; // @[Bitwise.scala 48:55:@4242.4]
  assign _GEN_736 = {{1'd0}, _T_6293}; // @[Bitwise.scala 48:55:@4243.4]
  assign _T_6296 = _GEN_736 + _T_6295; // @[Bitwise.scala 48:55:@4243.4]
  assign _T_6297 = _T_6292 + _T_6296; // @[Bitwise.scala 48:55:@4244.4]
  assign _T_6298 = _T_6259 + _T_6260; // @[Bitwise.scala 48:55:@4245.4]
  assign _T_6299 = _T_6262 + _T_6263; // @[Bitwise.scala 48:55:@4246.4]
  assign _GEN_737 = {{1'd0}, _T_6261}; // @[Bitwise.scala 48:55:@4247.4]
  assign _T_6300 = _GEN_737 + _T_6299; // @[Bitwise.scala 48:55:@4247.4]
  assign _GEN_738 = {{1'd0}, _T_6298}; // @[Bitwise.scala 48:55:@4248.4]
  assign _T_6301 = _GEN_738 + _T_6300; // @[Bitwise.scala 48:55:@4248.4]
  assign _T_6302 = _T_6264 + _T_6265; // @[Bitwise.scala 48:55:@4249.4]
  assign _T_6303 = _T_6267 + _T_6268; // @[Bitwise.scala 48:55:@4250.4]
  assign _GEN_739 = {{1'd0}, _T_6266}; // @[Bitwise.scala 48:55:@4251.4]
  assign _T_6304 = _GEN_739 + _T_6303; // @[Bitwise.scala 48:55:@4251.4]
  assign _GEN_740 = {{1'd0}, _T_6302}; // @[Bitwise.scala 48:55:@4252.4]
  assign _T_6305 = _GEN_740 + _T_6304; // @[Bitwise.scala 48:55:@4252.4]
  assign _T_6306 = _T_6301 + _T_6305; // @[Bitwise.scala 48:55:@4253.4]
  assign _T_6307 = _T_6297 + _T_6306; // @[Bitwise.scala 48:55:@4254.4]
  assign _T_6308 = _T_6269 + _T_6270; // @[Bitwise.scala 48:55:@4255.4]
  assign _T_6309 = _T_6272 + _T_6273; // @[Bitwise.scala 48:55:@4256.4]
  assign _GEN_741 = {{1'd0}, _T_6271}; // @[Bitwise.scala 48:55:@4257.4]
  assign _T_6310 = _GEN_741 + _T_6309; // @[Bitwise.scala 48:55:@4257.4]
  assign _GEN_742 = {{1'd0}, _T_6308}; // @[Bitwise.scala 48:55:@4258.4]
  assign _T_6311 = _GEN_742 + _T_6310; // @[Bitwise.scala 48:55:@4258.4]
  assign _T_6312 = _T_6274 + _T_6275; // @[Bitwise.scala 48:55:@4259.4]
  assign _T_6313 = _T_6277 + _T_6278; // @[Bitwise.scala 48:55:@4260.4]
  assign _GEN_743 = {{1'd0}, _T_6276}; // @[Bitwise.scala 48:55:@4261.4]
  assign _T_6314 = _GEN_743 + _T_6313; // @[Bitwise.scala 48:55:@4261.4]
  assign _GEN_744 = {{1'd0}, _T_6312}; // @[Bitwise.scala 48:55:@4262.4]
  assign _T_6315 = _GEN_744 + _T_6314; // @[Bitwise.scala 48:55:@4262.4]
  assign _T_6316 = _T_6311 + _T_6315; // @[Bitwise.scala 48:55:@4263.4]
  assign _T_6317 = _T_6279 + _T_6280; // @[Bitwise.scala 48:55:@4264.4]
  assign _T_6318 = _T_6282 + _T_6283; // @[Bitwise.scala 48:55:@4265.4]
  assign _GEN_745 = {{1'd0}, _T_6281}; // @[Bitwise.scala 48:55:@4266.4]
  assign _T_6319 = _GEN_745 + _T_6318; // @[Bitwise.scala 48:55:@4266.4]
  assign _GEN_746 = {{1'd0}, _T_6317}; // @[Bitwise.scala 48:55:@4267.4]
  assign _T_6320 = _GEN_746 + _T_6319; // @[Bitwise.scala 48:55:@4267.4]
  assign _T_6321 = _T_6284 + _T_6285; // @[Bitwise.scala 48:55:@4268.4]
  assign _T_6322 = _T_6287 + _T_6288; // @[Bitwise.scala 48:55:@4269.4]
  assign _GEN_747 = {{1'd0}, _T_6286}; // @[Bitwise.scala 48:55:@4270.4]
  assign _T_6323 = _GEN_747 + _T_6322; // @[Bitwise.scala 48:55:@4270.4]
  assign _GEN_748 = {{1'd0}, _T_6321}; // @[Bitwise.scala 48:55:@4271.4]
  assign _T_6324 = _GEN_748 + _T_6323; // @[Bitwise.scala 48:55:@4271.4]
  assign _T_6325 = _T_6320 + _T_6324; // @[Bitwise.scala 48:55:@4272.4]
  assign _T_6326 = _T_6316 + _T_6325; // @[Bitwise.scala 48:55:@4273.4]
  assign _T_6327 = _T_6307 + _T_6326; // @[Bitwise.scala 48:55:@4274.4]
  assign _T_6391 = _T_2230[40:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4339.4]
  assign _T_6392 = _T_6391[0]; // @[Bitwise.scala 50:65:@4340.4]
  assign _T_6393 = _T_6391[1]; // @[Bitwise.scala 50:65:@4341.4]
  assign _T_6394 = _T_6391[2]; // @[Bitwise.scala 50:65:@4342.4]
  assign _T_6395 = _T_6391[3]; // @[Bitwise.scala 50:65:@4343.4]
  assign _T_6396 = _T_6391[4]; // @[Bitwise.scala 50:65:@4344.4]
  assign _T_6397 = _T_6391[5]; // @[Bitwise.scala 50:65:@4345.4]
  assign _T_6398 = _T_6391[6]; // @[Bitwise.scala 50:65:@4346.4]
  assign _T_6399 = _T_6391[7]; // @[Bitwise.scala 50:65:@4347.4]
  assign _T_6400 = _T_6391[8]; // @[Bitwise.scala 50:65:@4348.4]
  assign _T_6401 = _T_6391[9]; // @[Bitwise.scala 50:65:@4349.4]
  assign _T_6402 = _T_6391[10]; // @[Bitwise.scala 50:65:@4350.4]
  assign _T_6403 = _T_6391[11]; // @[Bitwise.scala 50:65:@4351.4]
  assign _T_6404 = _T_6391[12]; // @[Bitwise.scala 50:65:@4352.4]
  assign _T_6405 = _T_6391[13]; // @[Bitwise.scala 50:65:@4353.4]
  assign _T_6406 = _T_6391[14]; // @[Bitwise.scala 50:65:@4354.4]
  assign _T_6407 = _T_6391[15]; // @[Bitwise.scala 50:65:@4355.4]
  assign _T_6408 = _T_6391[16]; // @[Bitwise.scala 50:65:@4356.4]
  assign _T_6409 = _T_6391[17]; // @[Bitwise.scala 50:65:@4357.4]
  assign _T_6410 = _T_6391[18]; // @[Bitwise.scala 50:65:@4358.4]
  assign _T_6411 = _T_6391[19]; // @[Bitwise.scala 50:65:@4359.4]
  assign _T_6412 = _T_6391[20]; // @[Bitwise.scala 50:65:@4360.4]
  assign _T_6413 = _T_6391[21]; // @[Bitwise.scala 50:65:@4361.4]
  assign _T_6414 = _T_6391[22]; // @[Bitwise.scala 50:65:@4362.4]
  assign _T_6415 = _T_6391[23]; // @[Bitwise.scala 50:65:@4363.4]
  assign _T_6416 = _T_6391[24]; // @[Bitwise.scala 50:65:@4364.4]
  assign _T_6417 = _T_6391[25]; // @[Bitwise.scala 50:65:@4365.4]
  assign _T_6418 = _T_6391[26]; // @[Bitwise.scala 50:65:@4366.4]
  assign _T_6419 = _T_6391[27]; // @[Bitwise.scala 50:65:@4367.4]
  assign _T_6420 = _T_6391[28]; // @[Bitwise.scala 50:65:@4368.4]
  assign _T_6421 = _T_6391[29]; // @[Bitwise.scala 50:65:@4369.4]
  assign _T_6422 = _T_6391[30]; // @[Bitwise.scala 50:65:@4370.4]
  assign _T_6423 = _T_6391[31]; // @[Bitwise.scala 50:65:@4371.4]
  assign _T_6424 = _T_6391[32]; // @[Bitwise.scala 50:65:@4372.4]
  assign _T_6425 = _T_6391[33]; // @[Bitwise.scala 50:65:@4373.4]
  assign _T_6426 = _T_6391[34]; // @[Bitwise.scala 50:65:@4374.4]
  assign _T_6427 = _T_6391[35]; // @[Bitwise.scala 50:65:@4375.4]
  assign _T_6428 = _T_6391[36]; // @[Bitwise.scala 50:65:@4376.4]
  assign _T_6429 = _T_6391[37]; // @[Bitwise.scala 50:65:@4377.4]
  assign _T_6430 = _T_6391[38]; // @[Bitwise.scala 50:65:@4378.4]
  assign _T_6431 = _T_6391[39]; // @[Bitwise.scala 50:65:@4379.4]
  assign _T_6432 = _T_6391[40]; // @[Bitwise.scala 50:65:@4380.4]
  assign _T_6433 = _T_6392 + _T_6393; // @[Bitwise.scala 48:55:@4381.4]
  assign _T_6434 = _T_6395 + _T_6396; // @[Bitwise.scala 48:55:@4382.4]
  assign _GEN_749 = {{1'd0}, _T_6394}; // @[Bitwise.scala 48:55:@4383.4]
  assign _T_6435 = _GEN_749 + _T_6434; // @[Bitwise.scala 48:55:@4383.4]
  assign _GEN_750 = {{1'd0}, _T_6433}; // @[Bitwise.scala 48:55:@4384.4]
  assign _T_6436 = _GEN_750 + _T_6435; // @[Bitwise.scala 48:55:@4384.4]
  assign _T_6437 = _T_6397 + _T_6398; // @[Bitwise.scala 48:55:@4385.4]
  assign _T_6438 = _T_6400 + _T_6401; // @[Bitwise.scala 48:55:@4386.4]
  assign _GEN_751 = {{1'd0}, _T_6399}; // @[Bitwise.scala 48:55:@4387.4]
  assign _T_6439 = _GEN_751 + _T_6438; // @[Bitwise.scala 48:55:@4387.4]
  assign _GEN_752 = {{1'd0}, _T_6437}; // @[Bitwise.scala 48:55:@4388.4]
  assign _T_6440 = _GEN_752 + _T_6439; // @[Bitwise.scala 48:55:@4388.4]
  assign _T_6441 = _T_6436 + _T_6440; // @[Bitwise.scala 48:55:@4389.4]
  assign _T_6442 = _T_6402 + _T_6403; // @[Bitwise.scala 48:55:@4390.4]
  assign _T_6443 = _T_6405 + _T_6406; // @[Bitwise.scala 48:55:@4391.4]
  assign _GEN_753 = {{1'd0}, _T_6404}; // @[Bitwise.scala 48:55:@4392.4]
  assign _T_6444 = _GEN_753 + _T_6443; // @[Bitwise.scala 48:55:@4392.4]
  assign _GEN_754 = {{1'd0}, _T_6442}; // @[Bitwise.scala 48:55:@4393.4]
  assign _T_6445 = _GEN_754 + _T_6444; // @[Bitwise.scala 48:55:@4393.4]
  assign _T_6446 = _T_6407 + _T_6408; // @[Bitwise.scala 48:55:@4394.4]
  assign _T_6447 = _T_6410 + _T_6411; // @[Bitwise.scala 48:55:@4395.4]
  assign _GEN_755 = {{1'd0}, _T_6409}; // @[Bitwise.scala 48:55:@4396.4]
  assign _T_6448 = _GEN_755 + _T_6447; // @[Bitwise.scala 48:55:@4396.4]
  assign _GEN_756 = {{1'd0}, _T_6446}; // @[Bitwise.scala 48:55:@4397.4]
  assign _T_6449 = _GEN_756 + _T_6448; // @[Bitwise.scala 48:55:@4397.4]
  assign _T_6450 = _T_6445 + _T_6449; // @[Bitwise.scala 48:55:@4398.4]
  assign _T_6451 = _T_6441 + _T_6450; // @[Bitwise.scala 48:55:@4399.4]
  assign _T_6452 = _T_6412 + _T_6413; // @[Bitwise.scala 48:55:@4400.4]
  assign _T_6453 = _T_6415 + _T_6416; // @[Bitwise.scala 48:55:@4401.4]
  assign _GEN_757 = {{1'd0}, _T_6414}; // @[Bitwise.scala 48:55:@4402.4]
  assign _T_6454 = _GEN_757 + _T_6453; // @[Bitwise.scala 48:55:@4402.4]
  assign _GEN_758 = {{1'd0}, _T_6452}; // @[Bitwise.scala 48:55:@4403.4]
  assign _T_6455 = _GEN_758 + _T_6454; // @[Bitwise.scala 48:55:@4403.4]
  assign _T_6456 = _T_6417 + _T_6418; // @[Bitwise.scala 48:55:@4404.4]
  assign _T_6457 = _T_6420 + _T_6421; // @[Bitwise.scala 48:55:@4405.4]
  assign _GEN_759 = {{1'd0}, _T_6419}; // @[Bitwise.scala 48:55:@4406.4]
  assign _T_6458 = _GEN_759 + _T_6457; // @[Bitwise.scala 48:55:@4406.4]
  assign _GEN_760 = {{1'd0}, _T_6456}; // @[Bitwise.scala 48:55:@4407.4]
  assign _T_6459 = _GEN_760 + _T_6458; // @[Bitwise.scala 48:55:@4407.4]
  assign _T_6460 = _T_6455 + _T_6459; // @[Bitwise.scala 48:55:@4408.4]
  assign _T_6461 = _T_6422 + _T_6423; // @[Bitwise.scala 48:55:@4409.4]
  assign _T_6462 = _T_6425 + _T_6426; // @[Bitwise.scala 48:55:@4410.4]
  assign _GEN_761 = {{1'd0}, _T_6424}; // @[Bitwise.scala 48:55:@4411.4]
  assign _T_6463 = _GEN_761 + _T_6462; // @[Bitwise.scala 48:55:@4411.4]
  assign _GEN_762 = {{1'd0}, _T_6461}; // @[Bitwise.scala 48:55:@4412.4]
  assign _T_6464 = _GEN_762 + _T_6463; // @[Bitwise.scala 48:55:@4412.4]
  assign _T_6465 = _T_6428 + _T_6429; // @[Bitwise.scala 48:55:@4413.4]
  assign _GEN_763 = {{1'd0}, _T_6427}; // @[Bitwise.scala 48:55:@4414.4]
  assign _T_6466 = _GEN_763 + _T_6465; // @[Bitwise.scala 48:55:@4414.4]
  assign _T_6467 = _T_6431 + _T_6432; // @[Bitwise.scala 48:55:@4415.4]
  assign _GEN_764 = {{1'd0}, _T_6430}; // @[Bitwise.scala 48:55:@4416.4]
  assign _T_6468 = _GEN_764 + _T_6467; // @[Bitwise.scala 48:55:@4416.4]
  assign _T_6469 = _T_6466 + _T_6468; // @[Bitwise.scala 48:55:@4417.4]
  assign _T_6470 = _T_6464 + _T_6469; // @[Bitwise.scala 48:55:@4418.4]
  assign _T_6471 = _T_6460 + _T_6470; // @[Bitwise.scala 48:55:@4419.4]
  assign _T_6472 = _T_6451 + _T_6471; // @[Bitwise.scala 48:55:@4420.4]
  assign _T_6536 = _T_2230[41:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4485.4]
  assign _T_6537 = _T_6536[0]; // @[Bitwise.scala 50:65:@4486.4]
  assign _T_6538 = _T_6536[1]; // @[Bitwise.scala 50:65:@4487.4]
  assign _T_6539 = _T_6536[2]; // @[Bitwise.scala 50:65:@4488.4]
  assign _T_6540 = _T_6536[3]; // @[Bitwise.scala 50:65:@4489.4]
  assign _T_6541 = _T_6536[4]; // @[Bitwise.scala 50:65:@4490.4]
  assign _T_6542 = _T_6536[5]; // @[Bitwise.scala 50:65:@4491.4]
  assign _T_6543 = _T_6536[6]; // @[Bitwise.scala 50:65:@4492.4]
  assign _T_6544 = _T_6536[7]; // @[Bitwise.scala 50:65:@4493.4]
  assign _T_6545 = _T_6536[8]; // @[Bitwise.scala 50:65:@4494.4]
  assign _T_6546 = _T_6536[9]; // @[Bitwise.scala 50:65:@4495.4]
  assign _T_6547 = _T_6536[10]; // @[Bitwise.scala 50:65:@4496.4]
  assign _T_6548 = _T_6536[11]; // @[Bitwise.scala 50:65:@4497.4]
  assign _T_6549 = _T_6536[12]; // @[Bitwise.scala 50:65:@4498.4]
  assign _T_6550 = _T_6536[13]; // @[Bitwise.scala 50:65:@4499.4]
  assign _T_6551 = _T_6536[14]; // @[Bitwise.scala 50:65:@4500.4]
  assign _T_6552 = _T_6536[15]; // @[Bitwise.scala 50:65:@4501.4]
  assign _T_6553 = _T_6536[16]; // @[Bitwise.scala 50:65:@4502.4]
  assign _T_6554 = _T_6536[17]; // @[Bitwise.scala 50:65:@4503.4]
  assign _T_6555 = _T_6536[18]; // @[Bitwise.scala 50:65:@4504.4]
  assign _T_6556 = _T_6536[19]; // @[Bitwise.scala 50:65:@4505.4]
  assign _T_6557 = _T_6536[20]; // @[Bitwise.scala 50:65:@4506.4]
  assign _T_6558 = _T_6536[21]; // @[Bitwise.scala 50:65:@4507.4]
  assign _T_6559 = _T_6536[22]; // @[Bitwise.scala 50:65:@4508.4]
  assign _T_6560 = _T_6536[23]; // @[Bitwise.scala 50:65:@4509.4]
  assign _T_6561 = _T_6536[24]; // @[Bitwise.scala 50:65:@4510.4]
  assign _T_6562 = _T_6536[25]; // @[Bitwise.scala 50:65:@4511.4]
  assign _T_6563 = _T_6536[26]; // @[Bitwise.scala 50:65:@4512.4]
  assign _T_6564 = _T_6536[27]; // @[Bitwise.scala 50:65:@4513.4]
  assign _T_6565 = _T_6536[28]; // @[Bitwise.scala 50:65:@4514.4]
  assign _T_6566 = _T_6536[29]; // @[Bitwise.scala 50:65:@4515.4]
  assign _T_6567 = _T_6536[30]; // @[Bitwise.scala 50:65:@4516.4]
  assign _T_6568 = _T_6536[31]; // @[Bitwise.scala 50:65:@4517.4]
  assign _T_6569 = _T_6536[32]; // @[Bitwise.scala 50:65:@4518.4]
  assign _T_6570 = _T_6536[33]; // @[Bitwise.scala 50:65:@4519.4]
  assign _T_6571 = _T_6536[34]; // @[Bitwise.scala 50:65:@4520.4]
  assign _T_6572 = _T_6536[35]; // @[Bitwise.scala 50:65:@4521.4]
  assign _T_6573 = _T_6536[36]; // @[Bitwise.scala 50:65:@4522.4]
  assign _T_6574 = _T_6536[37]; // @[Bitwise.scala 50:65:@4523.4]
  assign _T_6575 = _T_6536[38]; // @[Bitwise.scala 50:65:@4524.4]
  assign _T_6576 = _T_6536[39]; // @[Bitwise.scala 50:65:@4525.4]
  assign _T_6577 = _T_6536[40]; // @[Bitwise.scala 50:65:@4526.4]
  assign _T_6578 = _T_6536[41]; // @[Bitwise.scala 50:65:@4527.4]
  assign _T_6579 = _T_6537 + _T_6538; // @[Bitwise.scala 48:55:@4528.4]
  assign _T_6580 = _T_6540 + _T_6541; // @[Bitwise.scala 48:55:@4529.4]
  assign _GEN_765 = {{1'd0}, _T_6539}; // @[Bitwise.scala 48:55:@4530.4]
  assign _T_6581 = _GEN_765 + _T_6580; // @[Bitwise.scala 48:55:@4530.4]
  assign _GEN_766 = {{1'd0}, _T_6579}; // @[Bitwise.scala 48:55:@4531.4]
  assign _T_6582 = _GEN_766 + _T_6581; // @[Bitwise.scala 48:55:@4531.4]
  assign _T_6583 = _T_6542 + _T_6543; // @[Bitwise.scala 48:55:@4532.4]
  assign _T_6584 = _T_6545 + _T_6546; // @[Bitwise.scala 48:55:@4533.4]
  assign _GEN_767 = {{1'd0}, _T_6544}; // @[Bitwise.scala 48:55:@4534.4]
  assign _T_6585 = _GEN_767 + _T_6584; // @[Bitwise.scala 48:55:@4534.4]
  assign _GEN_768 = {{1'd0}, _T_6583}; // @[Bitwise.scala 48:55:@4535.4]
  assign _T_6586 = _GEN_768 + _T_6585; // @[Bitwise.scala 48:55:@4535.4]
  assign _T_6587 = _T_6582 + _T_6586; // @[Bitwise.scala 48:55:@4536.4]
  assign _T_6588 = _T_6547 + _T_6548; // @[Bitwise.scala 48:55:@4537.4]
  assign _T_6589 = _T_6550 + _T_6551; // @[Bitwise.scala 48:55:@4538.4]
  assign _GEN_769 = {{1'd0}, _T_6549}; // @[Bitwise.scala 48:55:@4539.4]
  assign _T_6590 = _GEN_769 + _T_6589; // @[Bitwise.scala 48:55:@4539.4]
  assign _GEN_770 = {{1'd0}, _T_6588}; // @[Bitwise.scala 48:55:@4540.4]
  assign _T_6591 = _GEN_770 + _T_6590; // @[Bitwise.scala 48:55:@4540.4]
  assign _T_6592 = _T_6553 + _T_6554; // @[Bitwise.scala 48:55:@4541.4]
  assign _GEN_771 = {{1'd0}, _T_6552}; // @[Bitwise.scala 48:55:@4542.4]
  assign _T_6593 = _GEN_771 + _T_6592; // @[Bitwise.scala 48:55:@4542.4]
  assign _T_6594 = _T_6556 + _T_6557; // @[Bitwise.scala 48:55:@4543.4]
  assign _GEN_772 = {{1'd0}, _T_6555}; // @[Bitwise.scala 48:55:@4544.4]
  assign _T_6595 = _GEN_772 + _T_6594; // @[Bitwise.scala 48:55:@4544.4]
  assign _T_6596 = _T_6593 + _T_6595; // @[Bitwise.scala 48:55:@4545.4]
  assign _T_6597 = _T_6591 + _T_6596; // @[Bitwise.scala 48:55:@4546.4]
  assign _T_6598 = _T_6587 + _T_6597; // @[Bitwise.scala 48:55:@4547.4]
  assign _T_6599 = _T_6558 + _T_6559; // @[Bitwise.scala 48:55:@4548.4]
  assign _T_6600 = _T_6561 + _T_6562; // @[Bitwise.scala 48:55:@4549.4]
  assign _GEN_773 = {{1'd0}, _T_6560}; // @[Bitwise.scala 48:55:@4550.4]
  assign _T_6601 = _GEN_773 + _T_6600; // @[Bitwise.scala 48:55:@4550.4]
  assign _GEN_774 = {{1'd0}, _T_6599}; // @[Bitwise.scala 48:55:@4551.4]
  assign _T_6602 = _GEN_774 + _T_6601; // @[Bitwise.scala 48:55:@4551.4]
  assign _T_6603 = _T_6563 + _T_6564; // @[Bitwise.scala 48:55:@4552.4]
  assign _T_6604 = _T_6566 + _T_6567; // @[Bitwise.scala 48:55:@4553.4]
  assign _GEN_775 = {{1'd0}, _T_6565}; // @[Bitwise.scala 48:55:@4554.4]
  assign _T_6605 = _GEN_775 + _T_6604; // @[Bitwise.scala 48:55:@4554.4]
  assign _GEN_776 = {{1'd0}, _T_6603}; // @[Bitwise.scala 48:55:@4555.4]
  assign _T_6606 = _GEN_776 + _T_6605; // @[Bitwise.scala 48:55:@4555.4]
  assign _T_6607 = _T_6602 + _T_6606; // @[Bitwise.scala 48:55:@4556.4]
  assign _T_6608 = _T_6568 + _T_6569; // @[Bitwise.scala 48:55:@4557.4]
  assign _T_6609 = _T_6571 + _T_6572; // @[Bitwise.scala 48:55:@4558.4]
  assign _GEN_777 = {{1'd0}, _T_6570}; // @[Bitwise.scala 48:55:@4559.4]
  assign _T_6610 = _GEN_777 + _T_6609; // @[Bitwise.scala 48:55:@4559.4]
  assign _GEN_778 = {{1'd0}, _T_6608}; // @[Bitwise.scala 48:55:@4560.4]
  assign _T_6611 = _GEN_778 + _T_6610; // @[Bitwise.scala 48:55:@4560.4]
  assign _T_6612 = _T_6574 + _T_6575; // @[Bitwise.scala 48:55:@4561.4]
  assign _GEN_779 = {{1'd0}, _T_6573}; // @[Bitwise.scala 48:55:@4562.4]
  assign _T_6613 = _GEN_779 + _T_6612; // @[Bitwise.scala 48:55:@4562.4]
  assign _T_6614 = _T_6577 + _T_6578; // @[Bitwise.scala 48:55:@4563.4]
  assign _GEN_780 = {{1'd0}, _T_6576}; // @[Bitwise.scala 48:55:@4564.4]
  assign _T_6615 = _GEN_780 + _T_6614; // @[Bitwise.scala 48:55:@4564.4]
  assign _T_6616 = _T_6613 + _T_6615; // @[Bitwise.scala 48:55:@4565.4]
  assign _T_6617 = _T_6611 + _T_6616; // @[Bitwise.scala 48:55:@4566.4]
  assign _T_6618 = _T_6607 + _T_6617; // @[Bitwise.scala 48:55:@4567.4]
  assign _T_6619 = _T_6598 + _T_6618; // @[Bitwise.scala 48:55:@4568.4]
  assign _T_6683 = _T_2230[42:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4633.4]
  assign _T_6684 = _T_6683[0]; // @[Bitwise.scala 50:65:@4634.4]
  assign _T_6685 = _T_6683[1]; // @[Bitwise.scala 50:65:@4635.4]
  assign _T_6686 = _T_6683[2]; // @[Bitwise.scala 50:65:@4636.4]
  assign _T_6687 = _T_6683[3]; // @[Bitwise.scala 50:65:@4637.4]
  assign _T_6688 = _T_6683[4]; // @[Bitwise.scala 50:65:@4638.4]
  assign _T_6689 = _T_6683[5]; // @[Bitwise.scala 50:65:@4639.4]
  assign _T_6690 = _T_6683[6]; // @[Bitwise.scala 50:65:@4640.4]
  assign _T_6691 = _T_6683[7]; // @[Bitwise.scala 50:65:@4641.4]
  assign _T_6692 = _T_6683[8]; // @[Bitwise.scala 50:65:@4642.4]
  assign _T_6693 = _T_6683[9]; // @[Bitwise.scala 50:65:@4643.4]
  assign _T_6694 = _T_6683[10]; // @[Bitwise.scala 50:65:@4644.4]
  assign _T_6695 = _T_6683[11]; // @[Bitwise.scala 50:65:@4645.4]
  assign _T_6696 = _T_6683[12]; // @[Bitwise.scala 50:65:@4646.4]
  assign _T_6697 = _T_6683[13]; // @[Bitwise.scala 50:65:@4647.4]
  assign _T_6698 = _T_6683[14]; // @[Bitwise.scala 50:65:@4648.4]
  assign _T_6699 = _T_6683[15]; // @[Bitwise.scala 50:65:@4649.4]
  assign _T_6700 = _T_6683[16]; // @[Bitwise.scala 50:65:@4650.4]
  assign _T_6701 = _T_6683[17]; // @[Bitwise.scala 50:65:@4651.4]
  assign _T_6702 = _T_6683[18]; // @[Bitwise.scala 50:65:@4652.4]
  assign _T_6703 = _T_6683[19]; // @[Bitwise.scala 50:65:@4653.4]
  assign _T_6704 = _T_6683[20]; // @[Bitwise.scala 50:65:@4654.4]
  assign _T_6705 = _T_6683[21]; // @[Bitwise.scala 50:65:@4655.4]
  assign _T_6706 = _T_6683[22]; // @[Bitwise.scala 50:65:@4656.4]
  assign _T_6707 = _T_6683[23]; // @[Bitwise.scala 50:65:@4657.4]
  assign _T_6708 = _T_6683[24]; // @[Bitwise.scala 50:65:@4658.4]
  assign _T_6709 = _T_6683[25]; // @[Bitwise.scala 50:65:@4659.4]
  assign _T_6710 = _T_6683[26]; // @[Bitwise.scala 50:65:@4660.4]
  assign _T_6711 = _T_6683[27]; // @[Bitwise.scala 50:65:@4661.4]
  assign _T_6712 = _T_6683[28]; // @[Bitwise.scala 50:65:@4662.4]
  assign _T_6713 = _T_6683[29]; // @[Bitwise.scala 50:65:@4663.4]
  assign _T_6714 = _T_6683[30]; // @[Bitwise.scala 50:65:@4664.4]
  assign _T_6715 = _T_6683[31]; // @[Bitwise.scala 50:65:@4665.4]
  assign _T_6716 = _T_6683[32]; // @[Bitwise.scala 50:65:@4666.4]
  assign _T_6717 = _T_6683[33]; // @[Bitwise.scala 50:65:@4667.4]
  assign _T_6718 = _T_6683[34]; // @[Bitwise.scala 50:65:@4668.4]
  assign _T_6719 = _T_6683[35]; // @[Bitwise.scala 50:65:@4669.4]
  assign _T_6720 = _T_6683[36]; // @[Bitwise.scala 50:65:@4670.4]
  assign _T_6721 = _T_6683[37]; // @[Bitwise.scala 50:65:@4671.4]
  assign _T_6722 = _T_6683[38]; // @[Bitwise.scala 50:65:@4672.4]
  assign _T_6723 = _T_6683[39]; // @[Bitwise.scala 50:65:@4673.4]
  assign _T_6724 = _T_6683[40]; // @[Bitwise.scala 50:65:@4674.4]
  assign _T_6725 = _T_6683[41]; // @[Bitwise.scala 50:65:@4675.4]
  assign _T_6726 = _T_6683[42]; // @[Bitwise.scala 50:65:@4676.4]
  assign _T_6727 = _T_6684 + _T_6685; // @[Bitwise.scala 48:55:@4677.4]
  assign _T_6728 = _T_6687 + _T_6688; // @[Bitwise.scala 48:55:@4678.4]
  assign _GEN_781 = {{1'd0}, _T_6686}; // @[Bitwise.scala 48:55:@4679.4]
  assign _T_6729 = _GEN_781 + _T_6728; // @[Bitwise.scala 48:55:@4679.4]
  assign _GEN_782 = {{1'd0}, _T_6727}; // @[Bitwise.scala 48:55:@4680.4]
  assign _T_6730 = _GEN_782 + _T_6729; // @[Bitwise.scala 48:55:@4680.4]
  assign _T_6731 = _T_6689 + _T_6690; // @[Bitwise.scala 48:55:@4681.4]
  assign _T_6732 = _T_6692 + _T_6693; // @[Bitwise.scala 48:55:@4682.4]
  assign _GEN_783 = {{1'd0}, _T_6691}; // @[Bitwise.scala 48:55:@4683.4]
  assign _T_6733 = _GEN_783 + _T_6732; // @[Bitwise.scala 48:55:@4683.4]
  assign _GEN_784 = {{1'd0}, _T_6731}; // @[Bitwise.scala 48:55:@4684.4]
  assign _T_6734 = _GEN_784 + _T_6733; // @[Bitwise.scala 48:55:@4684.4]
  assign _T_6735 = _T_6730 + _T_6734; // @[Bitwise.scala 48:55:@4685.4]
  assign _T_6736 = _T_6694 + _T_6695; // @[Bitwise.scala 48:55:@4686.4]
  assign _T_6737 = _T_6697 + _T_6698; // @[Bitwise.scala 48:55:@4687.4]
  assign _GEN_785 = {{1'd0}, _T_6696}; // @[Bitwise.scala 48:55:@4688.4]
  assign _T_6738 = _GEN_785 + _T_6737; // @[Bitwise.scala 48:55:@4688.4]
  assign _GEN_786 = {{1'd0}, _T_6736}; // @[Bitwise.scala 48:55:@4689.4]
  assign _T_6739 = _GEN_786 + _T_6738; // @[Bitwise.scala 48:55:@4689.4]
  assign _T_6740 = _T_6700 + _T_6701; // @[Bitwise.scala 48:55:@4690.4]
  assign _GEN_787 = {{1'd0}, _T_6699}; // @[Bitwise.scala 48:55:@4691.4]
  assign _T_6741 = _GEN_787 + _T_6740; // @[Bitwise.scala 48:55:@4691.4]
  assign _T_6742 = _T_6703 + _T_6704; // @[Bitwise.scala 48:55:@4692.4]
  assign _GEN_788 = {{1'd0}, _T_6702}; // @[Bitwise.scala 48:55:@4693.4]
  assign _T_6743 = _GEN_788 + _T_6742; // @[Bitwise.scala 48:55:@4693.4]
  assign _T_6744 = _T_6741 + _T_6743; // @[Bitwise.scala 48:55:@4694.4]
  assign _T_6745 = _T_6739 + _T_6744; // @[Bitwise.scala 48:55:@4695.4]
  assign _T_6746 = _T_6735 + _T_6745; // @[Bitwise.scala 48:55:@4696.4]
  assign _T_6747 = _T_6705 + _T_6706; // @[Bitwise.scala 48:55:@4697.4]
  assign _T_6748 = _T_6708 + _T_6709; // @[Bitwise.scala 48:55:@4698.4]
  assign _GEN_789 = {{1'd0}, _T_6707}; // @[Bitwise.scala 48:55:@4699.4]
  assign _T_6749 = _GEN_789 + _T_6748; // @[Bitwise.scala 48:55:@4699.4]
  assign _GEN_790 = {{1'd0}, _T_6747}; // @[Bitwise.scala 48:55:@4700.4]
  assign _T_6750 = _GEN_790 + _T_6749; // @[Bitwise.scala 48:55:@4700.4]
  assign _T_6751 = _T_6711 + _T_6712; // @[Bitwise.scala 48:55:@4701.4]
  assign _GEN_791 = {{1'd0}, _T_6710}; // @[Bitwise.scala 48:55:@4702.4]
  assign _T_6752 = _GEN_791 + _T_6751; // @[Bitwise.scala 48:55:@4702.4]
  assign _T_6753 = _T_6714 + _T_6715; // @[Bitwise.scala 48:55:@4703.4]
  assign _GEN_792 = {{1'd0}, _T_6713}; // @[Bitwise.scala 48:55:@4704.4]
  assign _T_6754 = _GEN_792 + _T_6753; // @[Bitwise.scala 48:55:@4704.4]
  assign _T_6755 = _T_6752 + _T_6754; // @[Bitwise.scala 48:55:@4705.4]
  assign _T_6756 = _T_6750 + _T_6755; // @[Bitwise.scala 48:55:@4706.4]
  assign _T_6757 = _T_6716 + _T_6717; // @[Bitwise.scala 48:55:@4707.4]
  assign _T_6758 = _T_6719 + _T_6720; // @[Bitwise.scala 48:55:@4708.4]
  assign _GEN_793 = {{1'd0}, _T_6718}; // @[Bitwise.scala 48:55:@4709.4]
  assign _T_6759 = _GEN_793 + _T_6758; // @[Bitwise.scala 48:55:@4709.4]
  assign _GEN_794 = {{1'd0}, _T_6757}; // @[Bitwise.scala 48:55:@4710.4]
  assign _T_6760 = _GEN_794 + _T_6759; // @[Bitwise.scala 48:55:@4710.4]
  assign _T_6761 = _T_6722 + _T_6723; // @[Bitwise.scala 48:55:@4711.4]
  assign _GEN_795 = {{1'd0}, _T_6721}; // @[Bitwise.scala 48:55:@4712.4]
  assign _T_6762 = _GEN_795 + _T_6761; // @[Bitwise.scala 48:55:@4712.4]
  assign _T_6763 = _T_6725 + _T_6726; // @[Bitwise.scala 48:55:@4713.4]
  assign _GEN_796 = {{1'd0}, _T_6724}; // @[Bitwise.scala 48:55:@4714.4]
  assign _T_6764 = _GEN_796 + _T_6763; // @[Bitwise.scala 48:55:@4714.4]
  assign _T_6765 = _T_6762 + _T_6764; // @[Bitwise.scala 48:55:@4715.4]
  assign _T_6766 = _T_6760 + _T_6765; // @[Bitwise.scala 48:55:@4716.4]
  assign _T_6767 = _T_6756 + _T_6766; // @[Bitwise.scala 48:55:@4717.4]
  assign _T_6768 = _T_6746 + _T_6767; // @[Bitwise.scala 48:55:@4718.4]
  assign _T_6832 = _T_2230[43:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4783.4]
  assign _T_6833 = _T_6832[0]; // @[Bitwise.scala 50:65:@4784.4]
  assign _T_6834 = _T_6832[1]; // @[Bitwise.scala 50:65:@4785.4]
  assign _T_6835 = _T_6832[2]; // @[Bitwise.scala 50:65:@4786.4]
  assign _T_6836 = _T_6832[3]; // @[Bitwise.scala 50:65:@4787.4]
  assign _T_6837 = _T_6832[4]; // @[Bitwise.scala 50:65:@4788.4]
  assign _T_6838 = _T_6832[5]; // @[Bitwise.scala 50:65:@4789.4]
  assign _T_6839 = _T_6832[6]; // @[Bitwise.scala 50:65:@4790.4]
  assign _T_6840 = _T_6832[7]; // @[Bitwise.scala 50:65:@4791.4]
  assign _T_6841 = _T_6832[8]; // @[Bitwise.scala 50:65:@4792.4]
  assign _T_6842 = _T_6832[9]; // @[Bitwise.scala 50:65:@4793.4]
  assign _T_6843 = _T_6832[10]; // @[Bitwise.scala 50:65:@4794.4]
  assign _T_6844 = _T_6832[11]; // @[Bitwise.scala 50:65:@4795.4]
  assign _T_6845 = _T_6832[12]; // @[Bitwise.scala 50:65:@4796.4]
  assign _T_6846 = _T_6832[13]; // @[Bitwise.scala 50:65:@4797.4]
  assign _T_6847 = _T_6832[14]; // @[Bitwise.scala 50:65:@4798.4]
  assign _T_6848 = _T_6832[15]; // @[Bitwise.scala 50:65:@4799.4]
  assign _T_6849 = _T_6832[16]; // @[Bitwise.scala 50:65:@4800.4]
  assign _T_6850 = _T_6832[17]; // @[Bitwise.scala 50:65:@4801.4]
  assign _T_6851 = _T_6832[18]; // @[Bitwise.scala 50:65:@4802.4]
  assign _T_6852 = _T_6832[19]; // @[Bitwise.scala 50:65:@4803.4]
  assign _T_6853 = _T_6832[20]; // @[Bitwise.scala 50:65:@4804.4]
  assign _T_6854 = _T_6832[21]; // @[Bitwise.scala 50:65:@4805.4]
  assign _T_6855 = _T_6832[22]; // @[Bitwise.scala 50:65:@4806.4]
  assign _T_6856 = _T_6832[23]; // @[Bitwise.scala 50:65:@4807.4]
  assign _T_6857 = _T_6832[24]; // @[Bitwise.scala 50:65:@4808.4]
  assign _T_6858 = _T_6832[25]; // @[Bitwise.scala 50:65:@4809.4]
  assign _T_6859 = _T_6832[26]; // @[Bitwise.scala 50:65:@4810.4]
  assign _T_6860 = _T_6832[27]; // @[Bitwise.scala 50:65:@4811.4]
  assign _T_6861 = _T_6832[28]; // @[Bitwise.scala 50:65:@4812.4]
  assign _T_6862 = _T_6832[29]; // @[Bitwise.scala 50:65:@4813.4]
  assign _T_6863 = _T_6832[30]; // @[Bitwise.scala 50:65:@4814.4]
  assign _T_6864 = _T_6832[31]; // @[Bitwise.scala 50:65:@4815.4]
  assign _T_6865 = _T_6832[32]; // @[Bitwise.scala 50:65:@4816.4]
  assign _T_6866 = _T_6832[33]; // @[Bitwise.scala 50:65:@4817.4]
  assign _T_6867 = _T_6832[34]; // @[Bitwise.scala 50:65:@4818.4]
  assign _T_6868 = _T_6832[35]; // @[Bitwise.scala 50:65:@4819.4]
  assign _T_6869 = _T_6832[36]; // @[Bitwise.scala 50:65:@4820.4]
  assign _T_6870 = _T_6832[37]; // @[Bitwise.scala 50:65:@4821.4]
  assign _T_6871 = _T_6832[38]; // @[Bitwise.scala 50:65:@4822.4]
  assign _T_6872 = _T_6832[39]; // @[Bitwise.scala 50:65:@4823.4]
  assign _T_6873 = _T_6832[40]; // @[Bitwise.scala 50:65:@4824.4]
  assign _T_6874 = _T_6832[41]; // @[Bitwise.scala 50:65:@4825.4]
  assign _T_6875 = _T_6832[42]; // @[Bitwise.scala 50:65:@4826.4]
  assign _T_6876 = _T_6832[43]; // @[Bitwise.scala 50:65:@4827.4]
  assign _T_6877 = _T_6833 + _T_6834; // @[Bitwise.scala 48:55:@4828.4]
  assign _T_6878 = _T_6836 + _T_6837; // @[Bitwise.scala 48:55:@4829.4]
  assign _GEN_797 = {{1'd0}, _T_6835}; // @[Bitwise.scala 48:55:@4830.4]
  assign _T_6879 = _GEN_797 + _T_6878; // @[Bitwise.scala 48:55:@4830.4]
  assign _GEN_798 = {{1'd0}, _T_6877}; // @[Bitwise.scala 48:55:@4831.4]
  assign _T_6880 = _GEN_798 + _T_6879; // @[Bitwise.scala 48:55:@4831.4]
  assign _T_6881 = _T_6839 + _T_6840; // @[Bitwise.scala 48:55:@4832.4]
  assign _GEN_799 = {{1'd0}, _T_6838}; // @[Bitwise.scala 48:55:@4833.4]
  assign _T_6882 = _GEN_799 + _T_6881; // @[Bitwise.scala 48:55:@4833.4]
  assign _T_6883 = _T_6842 + _T_6843; // @[Bitwise.scala 48:55:@4834.4]
  assign _GEN_800 = {{1'd0}, _T_6841}; // @[Bitwise.scala 48:55:@4835.4]
  assign _T_6884 = _GEN_800 + _T_6883; // @[Bitwise.scala 48:55:@4835.4]
  assign _T_6885 = _T_6882 + _T_6884; // @[Bitwise.scala 48:55:@4836.4]
  assign _T_6886 = _T_6880 + _T_6885; // @[Bitwise.scala 48:55:@4837.4]
  assign _T_6887 = _T_6844 + _T_6845; // @[Bitwise.scala 48:55:@4838.4]
  assign _T_6888 = _T_6847 + _T_6848; // @[Bitwise.scala 48:55:@4839.4]
  assign _GEN_801 = {{1'd0}, _T_6846}; // @[Bitwise.scala 48:55:@4840.4]
  assign _T_6889 = _GEN_801 + _T_6888; // @[Bitwise.scala 48:55:@4840.4]
  assign _GEN_802 = {{1'd0}, _T_6887}; // @[Bitwise.scala 48:55:@4841.4]
  assign _T_6890 = _GEN_802 + _T_6889; // @[Bitwise.scala 48:55:@4841.4]
  assign _T_6891 = _T_6850 + _T_6851; // @[Bitwise.scala 48:55:@4842.4]
  assign _GEN_803 = {{1'd0}, _T_6849}; // @[Bitwise.scala 48:55:@4843.4]
  assign _T_6892 = _GEN_803 + _T_6891; // @[Bitwise.scala 48:55:@4843.4]
  assign _T_6893 = _T_6853 + _T_6854; // @[Bitwise.scala 48:55:@4844.4]
  assign _GEN_804 = {{1'd0}, _T_6852}; // @[Bitwise.scala 48:55:@4845.4]
  assign _T_6894 = _GEN_804 + _T_6893; // @[Bitwise.scala 48:55:@4845.4]
  assign _T_6895 = _T_6892 + _T_6894; // @[Bitwise.scala 48:55:@4846.4]
  assign _T_6896 = _T_6890 + _T_6895; // @[Bitwise.scala 48:55:@4847.4]
  assign _T_6897 = _T_6886 + _T_6896; // @[Bitwise.scala 48:55:@4848.4]
  assign _T_6898 = _T_6855 + _T_6856; // @[Bitwise.scala 48:55:@4849.4]
  assign _T_6899 = _T_6858 + _T_6859; // @[Bitwise.scala 48:55:@4850.4]
  assign _GEN_805 = {{1'd0}, _T_6857}; // @[Bitwise.scala 48:55:@4851.4]
  assign _T_6900 = _GEN_805 + _T_6899; // @[Bitwise.scala 48:55:@4851.4]
  assign _GEN_806 = {{1'd0}, _T_6898}; // @[Bitwise.scala 48:55:@4852.4]
  assign _T_6901 = _GEN_806 + _T_6900; // @[Bitwise.scala 48:55:@4852.4]
  assign _T_6902 = _T_6861 + _T_6862; // @[Bitwise.scala 48:55:@4853.4]
  assign _GEN_807 = {{1'd0}, _T_6860}; // @[Bitwise.scala 48:55:@4854.4]
  assign _T_6903 = _GEN_807 + _T_6902; // @[Bitwise.scala 48:55:@4854.4]
  assign _T_6904 = _T_6864 + _T_6865; // @[Bitwise.scala 48:55:@4855.4]
  assign _GEN_808 = {{1'd0}, _T_6863}; // @[Bitwise.scala 48:55:@4856.4]
  assign _T_6905 = _GEN_808 + _T_6904; // @[Bitwise.scala 48:55:@4856.4]
  assign _T_6906 = _T_6903 + _T_6905; // @[Bitwise.scala 48:55:@4857.4]
  assign _T_6907 = _T_6901 + _T_6906; // @[Bitwise.scala 48:55:@4858.4]
  assign _T_6908 = _T_6866 + _T_6867; // @[Bitwise.scala 48:55:@4859.4]
  assign _T_6909 = _T_6869 + _T_6870; // @[Bitwise.scala 48:55:@4860.4]
  assign _GEN_809 = {{1'd0}, _T_6868}; // @[Bitwise.scala 48:55:@4861.4]
  assign _T_6910 = _GEN_809 + _T_6909; // @[Bitwise.scala 48:55:@4861.4]
  assign _GEN_810 = {{1'd0}, _T_6908}; // @[Bitwise.scala 48:55:@4862.4]
  assign _T_6911 = _GEN_810 + _T_6910; // @[Bitwise.scala 48:55:@4862.4]
  assign _T_6912 = _T_6872 + _T_6873; // @[Bitwise.scala 48:55:@4863.4]
  assign _GEN_811 = {{1'd0}, _T_6871}; // @[Bitwise.scala 48:55:@4864.4]
  assign _T_6913 = _GEN_811 + _T_6912; // @[Bitwise.scala 48:55:@4864.4]
  assign _T_6914 = _T_6875 + _T_6876; // @[Bitwise.scala 48:55:@4865.4]
  assign _GEN_812 = {{1'd0}, _T_6874}; // @[Bitwise.scala 48:55:@4866.4]
  assign _T_6915 = _GEN_812 + _T_6914; // @[Bitwise.scala 48:55:@4866.4]
  assign _T_6916 = _T_6913 + _T_6915; // @[Bitwise.scala 48:55:@4867.4]
  assign _T_6917 = _T_6911 + _T_6916; // @[Bitwise.scala 48:55:@4868.4]
  assign _T_6918 = _T_6907 + _T_6917; // @[Bitwise.scala 48:55:@4869.4]
  assign _T_6919 = _T_6897 + _T_6918; // @[Bitwise.scala 48:55:@4870.4]
  assign _T_6983 = _T_2230[44:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@4935.4]
  assign _T_6984 = _T_6983[0]; // @[Bitwise.scala 50:65:@4936.4]
  assign _T_6985 = _T_6983[1]; // @[Bitwise.scala 50:65:@4937.4]
  assign _T_6986 = _T_6983[2]; // @[Bitwise.scala 50:65:@4938.4]
  assign _T_6987 = _T_6983[3]; // @[Bitwise.scala 50:65:@4939.4]
  assign _T_6988 = _T_6983[4]; // @[Bitwise.scala 50:65:@4940.4]
  assign _T_6989 = _T_6983[5]; // @[Bitwise.scala 50:65:@4941.4]
  assign _T_6990 = _T_6983[6]; // @[Bitwise.scala 50:65:@4942.4]
  assign _T_6991 = _T_6983[7]; // @[Bitwise.scala 50:65:@4943.4]
  assign _T_6992 = _T_6983[8]; // @[Bitwise.scala 50:65:@4944.4]
  assign _T_6993 = _T_6983[9]; // @[Bitwise.scala 50:65:@4945.4]
  assign _T_6994 = _T_6983[10]; // @[Bitwise.scala 50:65:@4946.4]
  assign _T_6995 = _T_6983[11]; // @[Bitwise.scala 50:65:@4947.4]
  assign _T_6996 = _T_6983[12]; // @[Bitwise.scala 50:65:@4948.4]
  assign _T_6997 = _T_6983[13]; // @[Bitwise.scala 50:65:@4949.4]
  assign _T_6998 = _T_6983[14]; // @[Bitwise.scala 50:65:@4950.4]
  assign _T_6999 = _T_6983[15]; // @[Bitwise.scala 50:65:@4951.4]
  assign _T_7000 = _T_6983[16]; // @[Bitwise.scala 50:65:@4952.4]
  assign _T_7001 = _T_6983[17]; // @[Bitwise.scala 50:65:@4953.4]
  assign _T_7002 = _T_6983[18]; // @[Bitwise.scala 50:65:@4954.4]
  assign _T_7003 = _T_6983[19]; // @[Bitwise.scala 50:65:@4955.4]
  assign _T_7004 = _T_6983[20]; // @[Bitwise.scala 50:65:@4956.4]
  assign _T_7005 = _T_6983[21]; // @[Bitwise.scala 50:65:@4957.4]
  assign _T_7006 = _T_6983[22]; // @[Bitwise.scala 50:65:@4958.4]
  assign _T_7007 = _T_6983[23]; // @[Bitwise.scala 50:65:@4959.4]
  assign _T_7008 = _T_6983[24]; // @[Bitwise.scala 50:65:@4960.4]
  assign _T_7009 = _T_6983[25]; // @[Bitwise.scala 50:65:@4961.4]
  assign _T_7010 = _T_6983[26]; // @[Bitwise.scala 50:65:@4962.4]
  assign _T_7011 = _T_6983[27]; // @[Bitwise.scala 50:65:@4963.4]
  assign _T_7012 = _T_6983[28]; // @[Bitwise.scala 50:65:@4964.4]
  assign _T_7013 = _T_6983[29]; // @[Bitwise.scala 50:65:@4965.4]
  assign _T_7014 = _T_6983[30]; // @[Bitwise.scala 50:65:@4966.4]
  assign _T_7015 = _T_6983[31]; // @[Bitwise.scala 50:65:@4967.4]
  assign _T_7016 = _T_6983[32]; // @[Bitwise.scala 50:65:@4968.4]
  assign _T_7017 = _T_6983[33]; // @[Bitwise.scala 50:65:@4969.4]
  assign _T_7018 = _T_6983[34]; // @[Bitwise.scala 50:65:@4970.4]
  assign _T_7019 = _T_6983[35]; // @[Bitwise.scala 50:65:@4971.4]
  assign _T_7020 = _T_6983[36]; // @[Bitwise.scala 50:65:@4972.4]
  assign _T_7021 = _T_6983[37]; // @[Bitwise.scala 50:65:@4973.4]
  assign _T_7022 = _T_6983[38]; // @[Bitwise.scala 50:65:@4974.4]
  assign _T_7023 = _T_6983[39]; // @[Bitwise.scala 50:65:@4975.4]
  assign _T_7024 = _T_6983[40]; // @[Bitwise.scala 50:65:@4976.4]
  assign _T_7025 = _T_6983[41]; // @[Bitwise.scala 50:65:@4977.4]
  assign _T_7026 = _T_6983[42]; // @[Bitwise.scala 50:65:@4978.4]
  assign _T_7027 = _T_6983[43]; // @[Bitwise.scala 50:65:@4979.4]
  assign _T_7028 = _T_6983[44]; // @[Bitwise.scala 50:65:@4980.4]
  assign _T_7029 = _T_6984 + _T_6985; // @[Bitwise.scala 48:55:@4981.4]
  assign _T_7030 = _T_6987 + _T_6988; // @[Bitwise.scala 48:55:@4982.4]
  assign _GEN_813 = {{1'd0}, _T_6986}; // @[Bitwise.scala 48:55:@4983.4]
  assign _T_7031 = _GEN_813 + _T_7030; // @[Bitwise.scala 48:55:@4983.4]
  assign _GEN_814 = {{1'd0}, _T_7029}; // @[Bitwise.scala 48:55:@4984.4]
  assign _T_7032 = _GEN_814 + _T_7031; // @[Bitwise.scala 48:55:@4984.4]
  assign _T_7033 = _T_6990 + _T_6991; // @[Bitwise.scala 48:55:@4985.4]
  assign _GEN_815 = {{1'd0}, _T_6989}; // @[Bitwise.scala 48:55:@4986.4]
  assign _T_7034 = _GEN_815 + _T_7033; // @[Bitwise.scala 48:55:@4986.4]
  assign _T_7035 = _T_6993 + _T_6994; // @[Bitwise.scala 48:55:@4987.4]
  assign _GEN_816 = {{1'd0}, _T_6992}; // @[Bitwise.scala 48:55:@4988.4]
  assign _T_7036 = _GEN_816 + _T_7035; // @[Bitwise.scala 48:55:@4988.4]
  assign _T_7037 = _T_7034 + _T_7036; // @[Bitwise.scala 48:55:@4989.4]
  assign _T_7038 = _T_7032 + _T_7037; // @[Bitwise.scala 48:55:@4990.4]
  assign _T_7039 = _T_6995 + _T_6996; // @[Bitwise.scala 48:55:@4991.4]
  assign _T_7040 = _T_6998 + _T_6999; // @[Bitwise.scala 48:55:@4992.4]
  assign _GEN_817 = {{1'd0}, _T_6997}; // @[Bitwise.scala 48:55:@4993.4]
  assign _T_7041 = _GEN_817 + _T_7040; // @[Bitwise.scala 48:55:@4993.4]
  assign _GEN_818 = {{1'd0}, _T_7039}; // @[Bitwise.scala 48:55:@4994.4]
  assign _T_7042 = _GEN_818 + _T_7041; // @[Bitwise.scala 48:55:@4994.4]
  assign _T_7043 = _T_7001 + _T_7002; // @[Bitwise.scala 48:55:@4995.4]
  assign _GEN_819 = {{1'd0}, _T_7000}; // @[Bitwise.scala 48:55:@4996.4]
  assign _T_7044 = _GEN_819 + _T_7043; // @[Bitwise.scala 48:55:@4996.4]
  assign _T_7045 = _T_7004 + _T_7005; // @[Bitwise.scala 48:55:@4997.4]
  assign _GEN_820 = {{1'd0}, _T_7003}; // @[Bitwise.scala 48:55:@4998.4]
  assign _T_7046 = _GEN_820 + _T_7045; // @[Bitwise.scala 48:55:@4998.4]
  assign _T_7047 = _T_7044 + _T_7046; // @[Bitwise.scala 48:55:@4999.4]
  assign _T_7048 = _T_7042 + _T_7047; // @[Bitwise.scala 48:55:@5000.4]
  assign _T_7049 = _T_7038 + _T_7048; // @[Bitwise.scala 48:55:@5001.4]
  assign _T_7050 = _T_7006 + _T_7007; // @[Bitwise.scala 48:55:@5002.4]
  assign _T_7051 = _T_7009 + _T_7010; // @[Bitwise.scala 48:55:@5003.4]
  assign _GEN_821 = {{1'd0}, _T_7008}; // @[Bitwise.scala 48:55:@5004.4]
  assign _T_7052 = _GEN_821 + _T_7051; // @[Bitwise.scala 48:55:@5004.4]
  assign _GEN_822 = {{1'd0}, _T_7050}; // @[Bitwise.scala 48:55:@5005.4]
  assign _T_7053 = _GEN_822 + _T_7052; // @[Bitwise.scala 48:55:@5005.4]
  assign _T_7054 = _T_7012 + _T_7013; // @[Bitwise.scala 48:55:@5006.4]
  assign _GEN_823 = {{1'd0}, _T_7011}; // @[Bitwise.scala 48:55:@5007.4]
  assign _T_7055 = _GEN_823 + _T_7054; // @[Bitwise.scala 48:55:@5007.4]
  assign _T_7056 = _T_7015 + _T_7016; // @[Bitwise.scala 48:55:@5008.4]
  assign _GEN_824 = {{1'd0}, _T_7014}; // @[Bitwise.scala 48:55:@5009.4]
  assign _T_7057 = _GEN_824 + _T_7056; // @[Bitwise.scala 48:55:@5009.4]
  assign _T_7058 = _T_7055 + _T_7057; // @[Bitwise.scala 48:55:@5010.4]
  assign _T_7059 = _T_7053 + _T_7058; // @[Bitwise.scala 48:55:@5011.4]
  assign _T_7060 = _T_7018 + _T_7019; // @[Bitwise.scala 48:55:@5012.4]
  assign _GEN_825 = {{1'd0}, _T_7017}; // @[Bitwise.scala 48:55:@5013.4]
  assign _T_7061 = _GEN_825 + _T_7060; // @[Bitwise.scala 48:55:@5013.4]
  assign _T_7062 = _T_7021 + _T_7022; // @[Bitwise.scala 48:55:@5014.4]
  assign _GEN_826 = {{1'd0}, _T_7020}; // @[Bitwise.scala 48:55:@5015.4]
  assign _T_7063 = _GEN_826 + _T_7062; // @[Bitwise.scala 48:55:@5015.4]
  assign _T_7064 = _T_7061 + _T_7063; // @[Bitwise.scala 48:55:@5016.4]
  assign _T_7065 = _T_7024 + _T_7025; // @[Bitwise.scala 48:55:@5017.4]
  assign _GEN_827 = {{1'd0}, _T_7023}; // @[Bitwise.scala 48:55:@5018.4]
  assign _T_7066 = _GEN_827 + _T_7065; // @[Bitwise.scala 48:55:@5018.4]
  assign _T_7067 = _T_7027 + _T_7028; // @[Bitwise.scala 48:55:@5019.4]
  assign _GEN_828 = {{1'd0}, _T_7026}; // @[Bitwise.scala 48:55:@5020.4]
  assign _T_7068 = _GEN_828 + _T_7067; // @[Bitwise.scala 48:55:@5020.4]
  assign _T_7069 = _T_7066 + _T_7068; // @[Bitwise.scala 48:55:@5021.4]
  assign _T_7070 = _T_7064 + _T_7069; // @[Bitwise.scala 48:55:@5022.4]
  assign _T_7071 = _T_7059 + _T_7070; // @[Bitwise.scala 48:55:@5023.4]
  assign _T_7072 = _T_7049 + _T_7071; // @[Bitwise.scala 48:55:@5024.4]
  assign _T_7136 = _T_2230[45:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5089.4]
  assign _T_7137 = _T_7136[0]; // @[Bitwise.scala 50:65:@5090.4]
  assign _T_7138 = _T_7136[1]; // @[Bitwise.scala 50:65:@5091.4]
  assign _T_7139 = _T_7136[2]; // @[Bitwise.scala 50:65:@5092.4]
  assign _T_7140 = _T_7136[3]; // @[Bitwise.scala 50:65:@5093.4]
  assign _T_7141 = _T_7136[4]; // @[Bitwise.scala 50:65:@5094.4]
  assign _T_7142 = _T_7136[5]; // @[Bitwise.scala 50:65:@5095.4]
  assign _T_7143 = _T_7136[6]; // @[Bitwise.scala 50:65:@5096.4]
  assign _T_7144 = _T_7136[7]; // @[Bitwise.scala 50:65:@5097.4]
  assign _T_7145 = _T_7136[8]; // @[Bitwise.scala 50:65:@5098.4]
  assign _T_7146 = _T_7136[9]; // @[Bitwise.scala 50:65:@5099.4]
  assign _T_7147 = _T_7136[10]; // @[Bitwise.scala 50:65:@5100.4]
  assign _T_7148 = _T_7136[11]; // @[Bitwise.scala 50:65:@5101.4]
  assign _T_7149 = _T_7136[12]; // @[Bitwise.scala 50:65:@5102.4]
  assign _T_7150 = _T_7136[13]; // @[Bitwise.scala 50:65:@5103.4]
  assign _T_7151 = _T_7136[14]; // @[Bitwise.scala 50:65:@5104.4]
  assign _T_7152 = _T_7136[15]; // @[Bitwise.scala 50:65:@5105.4]
  assign _T_7153 = _T_7136[16]; // @[Bitwise.scala 50:65:@5106.4]
  assign _T_7154 = _T_7136[17]; // @[Bitwise.scala 50:65:@5107.4]
  assign _T_7155 = _T_7136[18]; // @[Bitwise.scala 50:65:@5108.4]
  assign _T_7156 = _T_7136[19]; // @[Bitwise.scala 50:65:@5109.4]
  assign _T_7157 = _T_7136[20]; // @[Bitwise.scala 50:65:@5110.4]
  assign _T_7158 = _T_7136[21]; // @[Bitwise.scala 50:65:@5111.4]
  assign _T_7159 = _T_7136[22]; // @[Bitwise.scala 50:65:@5112.4]
  assign _T_7160 = _T_7136[23]; // @[Bitwise.scala 50:65:@5113.4]
  assign _T_7161 = _T_7136[24]; // @[Bitwise.scala 50:65:@5114.4]
  assign _T_7162 = _T_7136[25]; // @[Bitwise.scala 50:65:@5115.4]
  assign _T_7163 = _T_7136[26]; // @[Bitwise.scala 50:65:@5116.4]
  assign _T_7164 = _T_7136[27]; // @[Bitwise.scala 50:65:@5117.4]
  assign _T_7165 = _T_7136[28]; // @[Bitwise.scala 50:65:@5118.4]
  assign _T_7166 = _T_7136[29]; // @[Bitwise.scala 50:65:@5119.4]
  assign _T_7167 = _T_7136[30]; // @[Bitwise.scala 50:65:@5120.4]
  assign _T_7168 = _T_7136[31]; // @[Bitwise.scala 50:65:@5121.4]
  assign _T_7169 = _T_7136[32]; // @[Bitwise.scala 50:65:@5122.4]
  assign _T_7170 = _T_7136[33]; // @[Bitwise.scala 50:65:@5123.4]
  assign _T_7171 = _T_7136[34]; // @[Bitwise.scala 50:65:@5124.4]
  assign _T_7172 = _T_7136[35]; // @[Bitwise.scala 50:65:@5125.4]
  assign _T_7173 = _T_7136[36]; // @[Bitwise.scala 50:65:@5126.4]
  assign _T_7174 = _T_7136[37]; // @[Bitwise.scala 50:65:@5127.4]
  assign _T_7175 = _T_7136[38]; // @[Bitwise.scala 50:65:@5128.4]
  assign _T_7176 = _T_7136[39]; // @[Bitwise.scala 50:65:@5129.4]
  assign _T_7177 = _T_7136[40]; // @[Bitwise.scala 50:65:@5130.4]
  assign _T_7178 = _T_7136[41]; // @[Bitwise.scala 50:65:@5131.4]
  assign _T_7179 = _T_7136[42]; // @[Bitwise.scala 50:65:@5132.4]
  assign _T_7180 = _T_7136[43]; // @[Bitwise.scala 50:65:@5133.4]
  assign _T_7181 = _T_7136[44]; // @[Bitwise.scala 50:65:@5134.4]
  assign _T_7182 = _T_7136[45]; // @[Bitwise.scala 50:65:@5135.4]
  assign _T_7183 = _T_7137 + _T_7138; // @[Bitwise.scala 48:55:@5136.4]
  assign _T_7184 = _T_7140 + _T_7141; // @[Bitwise.scala 48:55:@5137.4]
  assign _GEN_829 = {{1'd0}, _T_7139}; // @[Bitwise.scala 48:55:@5138.4]
  assign _T_7185 = _GEN_829 + _T_7184; // @[Bitwise.scala 48:55:@5138.4]
  assign _GEN_830 = {{1'd0}, _T_7183}; // @[Bitwise.scala 48:55:@5139.4]
  assign _T_7186 = _GEN_830 + _T_7185; // @[Bitwise.scala 48:55:@5139.4]
  assign _T_7187 = _T_7143 + _T_7144; // @[Bitwise.scala 48:55:@5140.4]
  assign _GEN_831 = {{1'd0}, _T_7142}; // @[Bitwise.scala 48:55:@5141.4]
  assign _T_7188 = _GEN_831 + _T_7187; // @[Bitwise.scala 48:55:@5141.4]
  assign _T_7189 = _T_7146 + _T_7147; // @[Bitwise.scala 48:55:@5142.4]
  assign _GEN_832 = {{1'd0}, _T_7145}; // @[Bitwise.scala 48:55:@5143.4]
  assign _T_7190 = _GEN_832 + _T_7189; // @[Bitwise.scala 48:55:@5143.4]
  assign _T_7191 = _T_7188 + _T_7190; // @[Bitwise.scala 48:55:@5144.4]
  assign _T_7192 = _T_7186 + _T_7191; // @[Bitwise.scala 48:55:@5145.4]
  assign _T_7193 = _T_7149 + _T_7150; // @[Bitwise.scala 48:55:@5146.4]
  assign _GEN_833 = {{1'd0}, _T_7148}; // @[Bitwise.scala 48:55:@5147.4]
  assign _T_7194 = _GEN_833 + _T_7193; // @[Bitwise.scala 48:55:@5147.4]
  assign _T_7195 = _T_7152 + _T_7153; // @[Bitwise.scala 48:55:@5148.4]
  assign _GEN_834 = {{1'd0}, _T_7151}; // @[Bitwise.scala 48:55:@5149.4]
  assign _T_7196 = _GEN_834 + _T_7195; // @[Bitwise.scala 48:55:@5149.4]
  assign _T_7197 = _T_7194 + _T_7196; // @[Bitwise.scala 48:55:@5150.4]
  assign _T_7198 = _T_7155 + _T_7156; // @[Bitwise.scala 48:55:@5151.4]
  assign _GEN_835 = {{1'd0}, _T_7154}; // @[Bitwise.scala 48:55:@5152.4]
  assign _T_7199 = _GEN_835 + _T_7198; // @[Bitwise.scala 48:55:@5152.4]
  assign _T_7200 = _T_7158 + _T_7159; // @[Bitwise.scala 48:55:@5153.4]
  assign _GEN_836 = {{1'd0}, _T_7157}; // @[Bitwise.scala 48:55:@5154.4]
  assign _T_7201 = _GEN_836 + _T_7200; // @[Bitwise.scala 48:55:@5154.4]
  assign _T_7202 = _T_7199 + _T_7201; // @[Bitwise.scala 48:55:@5155.4]
  assign _T_7203 = _T_7197 + _T_7202; // @[Bitwise.scala 48:55:@5156.4]
  assign _T_7204 = _T_7192 + _T_7203; // @[Bitwise.scala 48:55:@5157.4]
  assign _T_7205 = _T_7160 + _T_7161; // @[Bitwise.scala 48:55:@5158.4]
  assign _T_7206 = _T_7163 + _T_7164; // @[Bitwise.scala 48:55:@5159.4]
  assign _GEN_837 = {{1'd0}, _T_7162}; // @[Bitwise.scala 48:55:@5160.4]
  assign _T_7207 = _GEN_837 + _T_7206; // @[Bitwise.scala 48:55:@5160.4]
  assign _GEN_838 = {{1'd0}, _T_7205}; // @[Bitwise.scala 48:55:@5161.4]
  assign _T_7208 = _GEN_838 + _T_7207; // @[Bitwise.scala 48:55:@5161.4]
  assign _T_7209 = _T_7166 + _T_7167; // @[Bitwise.scala 48:55:@5162.4]
  assign _GEN_839 = {{1'd0}, _T_7165}; // @[Bitwise.scala 48:55:@5163.4]
  assign _T_7210 = _GEN_839 + _T_7209; // @[Bitwise.scala 48:55:@5163.4]
  assign _T_7211 = _T_7169 + _T_7170; // @[Bitwise.scala 48:55:@5164.4]
  assign _GEN_840 = {{1'd0}, _T_7168}; // @[Bitwise.scala 48:55:@5165.4]
  assign _T_7212 = _GEN_840 + _T_7211; // @[Bitwise.scala 48:55:@5165.4]
  assign _T_7213 = _T_7210 + _T_7212; // @[Bitwise.scala 48:55:@5166.4]
  assign _T_7214 = _T_7208 + _T_7213; // @[Bitwise.scala 48:55:@5167.4]
  assign _T_7215 = _T_7172 + _T_7173; // @[Bitwise.scala 48:55:@5168.4]
  assign _GEN_841 = {{1'd0}, _T_7171}; // @[Bitwise.scala 48:55:@5169.4]
  assign _T_7216 = _GEN_841 + _T_7215; // @[Bitwise.scala 48:55:@5169.4]
  assign _T_7217 = _T_7175 + _T_7176; // @[Bitwise.scala 48:55:@5170.4]
  assign _GEN_842 = {{1'd0}, _T_7174}; // @[Bitwise.scala 48:55:@5171.4]
  assign _T_7218 = _GEN_842 + _T_7217; // @[Bitwise.scala 48:55:@5171.4]
  assign _T_7219 = _T_7216 + _T_7218; // @[Bitwise.scala 48:55:@5172.4]
  assign _T_7220 = _T_7178 + _T_7179; // @[Bitwise.scala 48:55:@5173.4]
  assign _GEN_843 = {{1'd0}, _T_7177}; // @[Bitwise.scala 48:55:@5174.4]
  assign _T_7221 = _GEN_843 + _T_7220; // @[Bitwise.scala 48:55:@5174.4]
  assign _T_7222 = _T_7181 + _T_7182; // @[Bitwise.scala 48:55:@5175.4]
  assign _GEN_844 = {{1'd0}, _T_7180}; // @[Bitwise.scala 48:55:@5176.4]
  assign _T_7223 = _GEN_844 + _T_7222; // @[Bitwise.scala 48:55:@5176.4]
  assign _T_7224 = _T_7221 + _T_7223; // @[Bitwise.scala 48:55:@5177.4]
  assign _T_7225 = _T_7219 + _T_7224; // @[Bitwise.scala 48:55:@5178.4]
  assign _T_7226 = _T_7214 + _T_7225; // @[Bitwise.scala 48:55:@5179.4]
  assign _T_7227 = _T_7204 + _T_7226; // @[Bitwise.scala 48:55:@5180.4]
  assign _T_7291 = _T_2230[46:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5245.4]
  assign _T_7292 = _T_7291[0]; // @[Bitwise.scala 50:65:@5246.4]
  assign _T_7293 = _T_7291[1]; // @[Bitwise.scala 50:65:@5247.4]
  assign _T_7294 = _T_7291[2]; // @[Bitwise.scala 50:65:@5248.4]
  assign _T_7295 = _T_7291[3]; // @[Bitwise.scala 50:65:@5249.4]
  assign _T_7296 = _T_7291[4]; // @[Bitwise.scala 50:65:@5250.4]
  assign _T_7297 = _T_7291[5]; // @[Bitwise.scala 50:65:@5251.4]
  assign _T_7298 = _T_7291[6]; // @[Bitwise.scala 50:65:@5252.4]
  assign _T_7299 = _T_7291[7]; // @[Bitwise.scala 50:65:@5253.4]
  assign _T_7300 = _T_7291[8]; // @[Bitwise.scala 50:65:@5254.4]
  assign _T_7301 = _T_7291[9]; // @[Bitwise.scala 50:65:@5255.4]
  assign _T_7302 = _T_7291[10]; // @[Bitwise.scala 50:65:@5256.4]
  assign _T_7303 = _T_7291[11]; // @[Bitwise.scala 50:65:@5257.4]
  assign _T_7304 = _T_7291[12]; // @[Bitwise.scala 50:65:@5258.4]
  assign _T_7305 = _T_7291[13]; // @[Bitwise.scala 50:65:@5259.4]
  assign _T_7306 = _T_7291[14]; // @[Bitwise.scala 50:65:@5260.4]
  assign _T_7307 = _T_7291[15]; // @[Bitwise.scala 50:65:@5261.4]
  assign _T_7308 = _T_7291[16]; // @[Bitwise.scala 50:65:@5262.4]
  assign _T_7309 = _T_7291[17]; // @[Bitwise.scala 50:65:@5263.4]
  assign _T_7310 = _T_7291[18]; // @[Bitwise.scala 50:65:@5264.4]
  assign _T_7311 = _T_7291[19]; // @[Bitwise.scala 50:65:@5265.4]
  assign _T_7312 = _T_7291[20]; // @[Bitwise.scala 50:65:@5266.4]
  assign _T_7313 = _T_7291[21]; // @[Bitwise.scala 50:65:@5267.4]
  assign _T_7314 = _T_7291[22]; // @[Bitwise.scala 50:65:@5268.4]
  assign _T_7315 = _T_7291[23]; // @[Bitwise.scala 50:65:@5269.4]
  assign _T_7316 = _T_7291[24]; // @[Bitwise.scala 50:65:@5270.4]
  assign _T_7317 = _T_7291[25]; // @[Bitwise.scala 50:65:@5271.4]
  assign _T_7318 = _T_7291[26]; // @[Bitwise.scala 50:65:@5272.4]
  assign _T_7319 = _T_7291[27]; // @[Bitwise.scala 50:65:@5273.4]
  assign _T_7320 = _T_7291[28]; // @[Bitwise.scala 50:65:@5274.4]
  assign _T_7321 = _T_7291[29]; // @[Bitwise.scala 50:65:@5275.4]
  assign _T_7322 = _T_7291[30]; // @[Bitwise.scala 50:65:@5276.4]
  assign _T_7323 = _T_7291[31]; // @[Bitwise.scala 50:65:@5277.4]
  assign _T_7324 = _T_7291[32]; // @[Bitwise.scala 50:65:@5278.4]
  assign _T_7325 = _T_7291[33]; // @[Bitwise.scala 50:65:@5279.4]
  assign _T_7326 = _T_7291[34]; // @[Bitwise.scala 50:65:@5280.4]
  assign _T_7327 = _T_7291[35]; // @[Bitwise.scala 50:65:@5281.4]
  assign _T_7328 = _T_7291[36]; // @[Bitwise.scala 50:65:@5282.4]
  assign _T_7329 = _T_7291[37]; // @[Bitwise.scala 50:65:@5283.4]
  assign _T_7330 = _T_7291[38]; // @[Bitwise.scala 50:65:@5284.4]
  assign _T_7331 = _T_7291[39]; // @[Bitwise.scala 50:65:@5285.4]
  assign _T_7332 = _T_7291[40]; // @[Bitwise.scala 50:65:@5286.4]
  assign _T_7333 = _T_7291[41]; // @[Bitwise.scala 50:65:@5287.4]
  assign _T_7334 = _T_7291[42]; // @[Bitwise.scala 50:65:@5288.4]
  assign _T_7335 = _T_7291[43]; // @[Bitwise.scala 50:65:@5289.4]
  assign _T_7336 = _T_7291[44]; // @[Bitwise.scala 50:65:@5290.4]
  assign _T_7337 = _T_7291[45]; // @[Bitwise.scala 50:65:@5291.4]
  assign _T_7338 = _T_7291[46]; // @[Bitwise.scala 50:65:@5292.4]
  assign _T_7339 = _T_7292 + _T_7293; // @[Bitwise.scala 48:55:@5293.4]
  assign _T_7340 = _T_7295 + _T_7296; // @[Bitwise.scala 48:55:@5294.4]
  assign _GEN_845 = {{1'd0}, _T_7294}; // @[Bitwise.scala 48:55:@5295.4]
  assign _T_7341 = _GEN_845 + _T_7340; // @[Bitwise.scala 48:55:@5295.4]
  assign _GEN_846 = {{1'd0}, _T_7339}; // @[Bitwise.scala 48:55:@5296.4]
  assign _T_7342 = _GEN_846 + _T_7341; // @[Bitwise.scala 48:55:@5296.4]
  assign _T_7343 = _T_7298 + _T_7299; // @[Bitwise.scala 48:55:@5297.4]
  assign _GEN_847 = {{1'd0}, _T_7297}; // @[Bitwise.scala 48:55:@5298.4]
  assign _T_7344 = _GEN_847 + _T_7343; // @[Bitwise.scala 48:55:@5298.4]
  assign _T_7345 = _T_7301 + _T_7302; // @[Bitwise.scala 48:55:@5299.4]
  assign _GEN_848 = {{1'd0}, _T_7300}; // @[Bitwise.scala 48:55:@5300.4]
  assign _T_7346 = _GEN_848 + _T_7345; // @[Bitwise.scala 48:55:@5300.4]
  assign _T_7347 = _T_7344 + _T_7346; // @[Bitwise.scala 48:55:@5301.4]
  assign _T_7348 = _T_7342 + _T_7347; // @[Bitwise.scala 48:55:@5302.4]
  assign _T_7349 = _T_7304 + _T_7305; // @[Bitwise.scala 48:55:@5303.4]
  assign _GEN_849 = {{1'd0}, _T_7303}; // @[Bitwise.scala 48:55:@5304.4]
  assign _T_7350 = _GEN_849 + _T_7349; // @[Bitwise.scala 48:55:@5304.4]
  assign _T_7351 = _T_7307 + _T_7308; // @[Bitwise.scala 48:55:@5305.4]
  assign _GEN_850 = {{1'd0}, _T_7306}; // @[Bitwise.scala 48:55:@5306.4]
  assign _T_7352 = _GEN_850 + _T_7351; // @[Bitwise.scala 48:55:@5306.4]
  assign _T_7353 = _T_7350 + _T_7352; // @[Bitwise.scala 48:55:@5307.4]
  assign _T_7354 = _T_7310 + _T_7311; // @[Bitwise.scala 48:55:@5308.4]
  assign _GEN_851 = {{1'd0}, _T_7309}; // @[Bitwise.scala 48:55:@5309.4]
  assign _T_7355 = _GEN_851 + _T_7354; // @[Bitwise.scala 48:55:@5309.4]
  assign _T_7356 = _T_7313 + _T_7314; // @[Bitwise.scala 48:55:@5310.4]
  assign _GEN_852 = {{1'd0}, _T_7312}; // @[Bitwise.scala 48:55:@5311.4]
  assign _T_7357 = _GEN_852 + _T_7356; // @[Bitwise.scala 48:55:@5311.4]
  assign _T_7358 = _T_7355 + _T_7357; // @[Bitwise.scala 48:55:@5312.4]
  assign _T_7359 = _T_7353 + _T_7358; // @[Bitwise.scala 48:55:@5313.4]
  assign _T_7360 = _T_7348 + _T_7359; // @[Bitwise.scala 48:55:@5314.4]
  assign _T_7361 = _T_7316 + _T_7317; // @[Bitwise.scala 48:55:@5315.4]
  assign _GEN_853 = {{1'd0}, _T_7315}; // @[Bitwise.scala 48:55:@5316.4]
  assign _T_7362 = _GEN_853 + _T_7361; // @[Bitwise.scala 48:55:@5316.4]
  assign _T_7363 = _T_7319 + _T_7320; // @[Bitwise.scala 48:55:@5317.4]
  assign _GEN_854 = {{1'd0}, _T_7318}; // @[Bitwise.scala 48:55:@5318.4]
  assign _T_7364 = _GEN_854 + _T_7363; // @[Bitwise.scala 48:55:@5318.4]
  assign _T_7365 = _T_7362 + _T_7364; // @[Bitwise.scala 48:55:@5319.4]
  assign _T_7366 = _T_7322 + _T_7323; // @[Bitwise.scala 48:55:@5320.4]
  assign _GEN_855 = {{1'd0}, _T_7321}; // @[Bitwise.scala 48:55:@5321.4]
  assign _T_7367 = _GEN_855 + _T_7366; // @[Bitwise.scala 48:55:@5321.4]
  assign _T_7368 = _T_7325 + _T_7326; // @[Bitwise.scala 48:55:@5322.4]
  assign _GEN_856 = {{1'd0}, _T_7324}; // @[Bitwise.scala 48:55:@5323.4]
  assign _T_7369 = _GEN_856 + _T_7368; // @[Bitwise.scala 48:55:@5323.4]
  assign _T_7370 = _T_7367 + _T_7369; // @[Bitwise.scala 48:55:@5324.4]
  assign _T_7371 = _T_7365 + _T_7370; // @[Bitwise.scala 48:55:@5325.4]
  assign _T_7372 = _T_7328 + _T_7329; // @[Bitwise.scala 48:55:@5326.4]
  assign _GEN_857 = {{1'd0}, _T_7327}; // @[Bitwise.scala 48:55:@5327.4]
  assign _T_7373 = _GEN_857 + _T_7372; // @[Bitwise.scala 48:55:@5327.4]
  assign _T_7374 = _T_7331 + _T_7332; // @[Bitwise.scala 48:55:@5328.4]
  assign _GEN_858 = {{1'd0}, _T_7330}; // @[Bitwise.scala 48:55:@5329.4]
  assign _T_7375 = _GEN_858 + _T_7374; // @[Bitwise.scala 48:55:@5329.4]
  assign _T_7376 = _T_7373 + _T_7375; // @[Bitwise.scala 48:55:@5330.4]
  assign _T_7377 = _T_7334 + _T_7335; // @[Bitwise.scala 48:55:@5331.4]
  assign _GEN_859 = {{1'd0}, _T_7333}; // @[Bitwise.scala 48:55:@5332.4]
  assign _T_7378 = _GEN_859 + _T_7377; // @[Bitwise.scala 48:55:@5332.4]
  assign _T_7379 = _T_7337 + _T_7338; // @[Bitwise.scala 48:55:@5333.4]
  assign _GEN_860 = {{1'd0}, _T_7336}; // @[Bitwise.scala 48:55:@5334.4]
  assign _T_7380 = _GEN_860 + _T_7379; // @[Bitwise.scala 48:55:@5334.4]
  assign _T_7381 = _T_7378 + _T_7380; // @[Bitwise.scala 48:55:@5335.4]
  assign _T_7382 = _T_7376 + _T_7381; // @[Bitwise.scala 48:55:@5336.4]
  assign _T_7383 = _T_7371 + _T_7382; // @[Bitwise.scala 48:55:@5337.4]
  assign _T_7384 = _T_7360 + _T_7383; // @[Bitwise.scala 48:55:@5338.4]
  assign _T_7448 = _T_2230[47:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5403.4]
  assign _T_7449 = _T_7448[0]; // @[Bitwise.scala 50:65:@5404.4]
  assign _T_7450 = _T_7448[1]; // @[Bitwise.scala 50:65:@5405.4]
  assign _T_7451 = _T_7448[2]; // @[Bitwise.scala 50:65:@5406.4]
  assign _T_7452 = _T_7448[3]; // @[Bitwise.scala 50:65:@5407.4]
  assign _T_7453 = _T_7448[4]; // @[Bitwise.scala 50:65:@5408.4]
  assign _T_7454 = _T_7448[5]; // @[Bitwise.scala 50:65:@5409.4]
  assign _T_7455 = _T_7448[6]; // @[Bitwise.scala 50:65:@5410.4]
  assign _T_7456 = _T_7448[7]; // @[Bitwise.scala 50:65:@5411.4]
  assign _T_7457 = _T_7448[8]; // @[Bitwise.scala 50:65:@5412.4]
  assign _T_7458 = _T_7448[9]; // @[Bitwise.scala 50:65:@5413.4]
  assign _T_7459 = _T_7448[10]; // @[Bitwise.scala 50:65:@5414.4]
  assign _T_7460 = _T_7448[11]; // @[Bitwise.scala 50:65:@5415.4]
  assign _T_7461 = _T_7448[12]; // @[Bitwise.scala 50:65:@5416.4]
  assign _T_7462 = _T_7448[13]; // @[Bitwise.scala 50:65:@5417.4]
  assign _T_7463 = _T_7448[14]; // @[Bitwise.scala 50:65:@5418.4]
  assign _T_7464 = _T_7448[15]; // @[Bitwise.scala 50:65:@5419.4]
  assign _T_7465 = _T_7448[16]; // @[Bitwise.scala 50:65:@5420.4]
  assign _T_7466 = _T_7448[17]; // @[Bitwise.scala 50:65:@5421.4]
  assign _T_7467 = _T_7448[18]; // @[Bitwise.scala 50:65:@5422.4]
  assign _T_7468 = _T_7448[19]; // @[Bitwise.scala 50:65:@5423.4]
  assign _T_7469 = _T_7448[20]; // @[Bitwise.scala 50:65:@5424.4]
  assign _T_7470 = _T_7448[21]; // @[Bitwise.scala 50:65:@5425.4]
  assign _T_7471 = _T_7448[22]; // @[Bitwise.scala 50:65:@5426.4]
  assign _T_7472 = _T_7448[23]; // @[Bitwise.scala 50:65:@5427.4]
  assign _T_7473 = _T_7448[24]; // @[Bitwise.scala 50:65:@5428.4]
  assign _T_7474 = _T_7448[25]; // @[Bitwise.scala 50:65:@5429.4]
  assign _T_7475 = _T_7448[26]; // @[Bitwise.scala 50:65:@5430.4]
  assign _T_7476 = _T_7448[27]; // @[Bitwise.scala 50:65:@5431.4]
  assign _T_7477 = _T_7448[28]; // @[Bitwise.scala 50:65:@5432.4]
  assign _T_7478 = _T_7448[29]; // @[Bitwise.scala 50:65:@5433.4]
  assign _T_7479 = _T_7448[30]; // @[Bitwise.scala 50:65:@5434.4]
  assign _T_7480 = _T_7448[31]; // @[Bitwise.scala 50:65:@5435.4]
  assign _T_7481 = _T_7448[32]; // @[Bitwise.scala 50:65:@5436.4]
  assign _T_7482 = _T_7448[33]; // @[Bitwise.scala 50:65:@5437.4]
  assign _T_7483 = _T_7448[34]; // @[Bitwise.scala 50:65:@5438.4]
  assign _T_7484 = _T_7448[35]; // @[Bitwise.scala 50:65:@5439.4]
  assign _T_7485 = _T_7448[36]; // @[Bitwise.scala 50:65:@5440.4]
  assign _T_7486 = _T_7448[37]; // @[Bitwise.scala 50:65:@5441.4]
  assign _T_7487 = _T_7448[38]; // @[Bitwise.scala 50:65:@5442.4]
  assign _T_7488 = _T_7448[39]; // @[Bitwise.scala 50:65:@5443.4]
  assign _T_7489 = _T_7448[40]; // @[Bitwise.scala 50:65:@5444.4]
  assign _T_7490 = _T_7448[41]; // @[Bitwise.scala 50:65:@5445.4]
  assign _T_7491 = _T_7448[42]; // @[Bitwise.scala 50:65:@5446.4]
  assign _T_7492 = _T_7448[43]; // @[Bitwise.scala 50:65:@5447.4]
  assign _T_7493 = _T_7448[44]; // @[Bitwise.scala 50:65:@5448.4]
  assign _T_7494 = _T_7448[45]; // @[Bitwise.scala 50:65:@5449.4]
  assign _T_7495 = _T_7448[46]; // @[Bitwise.scala 50:65:@5450.4]
  assign _T_7496 = _T_7448[47]; // @[Bitwise.scala 50:65:@5451.4]
  assign _T_7497 = _T_7450 + _T_7451; // @[Bitwise.scala 48:55:@5452.4]
  assign _GEN_861 = {{1'd0}, _T_7449}; // @[Bitwise.scala 48:55:@5453.4]
  assign _T_7498 = _GEN_861 + _T_7497; // @[Bitwise.scala 48:55:@5453.4]
  assign _T_7499 = _T_7453 + _T_7454; // @[Bitwise.scala 48:55:@5454.4]
  assign _GEN_862 = {{1'd0}, _T_7452}; // @[Bitwise.scala 48:55:@5455.4]
  assign _T_7500 = _GEN_862 + _T_7499; // @[Bitwise.scala 48:55:@5455.4]
  assign _T_7501 = _T_7498 + _T_7500; // @[Bitwise.scala 48:55:@5456.4]
  assign _T_7502 = _T_7456 + _T_7457; // @[Bitwise.scala 48:55:@5457.4]
  assign _GEN_863 = {{1'd0}, _T_7455}; // @[Bitwise.scala 48:55:@5458.4]
  assign _T_7503 = _GEN_863 + _T_7502; // @[Bitwise.scala 48:55:@5458.4]
  assign _T_7504 = _T_7459 + _T_7460; // @[Bitwise.scala 48:55:@5459.4]
  assign _GEN_864 = {{1'd0}, _T_7458}; // @[Bitwise.scala 48:55:@5460.4]
  assign _T_7505 = _GEN_864 + _T_7504; // @[Bitwise.scala 48:55:@5460.4]
  assign _T_7506 = _T_7503 + _T_7505; // @[Bitwise.scala 48:55:@5461.4]
  assign _T_7507 = _T_7501 + _T_7506; // @[Bitwise.scala 48:55:@5462.4]
  assign _T_7508 = _T_7462 + _T_7463; // @[Bitwise.scala 48:55:@5463.4]
  assign _GEN_865 = {{1'd0}, _T_7461}; // @[Bitwise.scala 48:55:@5464.4]
  assign _T_7509 = _GEN_865 + _T_7508; // @[Bitwise.scala 48:55:@5464.4]
  assign _T_7510 = _T_7465 + _T_7466; // @[Bitwise.scala 48:55:@5465.4]
  assign _GEN_866 = {{1'd0}, _T_7464}; // @[Bitwise.scala 48:55:@5466.4]
  assign _T_7511 = _GEN_866 + _T_7510; // @[Bitwise.scala 48:55:@5466.4]
  assign _T_7512 = _T_7509 + _T_7511; // @[Bitwise.scala 48:55:@5467.4]
  assign _T_7513 = _T_7468 + _T_7469; // @[Bitwise.scala 48:55:@5468.4]
  assign _GEN_867 = {{1'd0}, _T_7467}; // @[Bitwise.scala 48:55:@5469.4]
  assign _T_7514 = _GEN_867 + _T_7513; // @[Bitwise.scala 48:55:@5469.4]
  assign _T_7515 = _T_7471 + _T_7472; // @[Bitwise.scala 48:55:@5470.4]
  assign _GEN_868 = {{1'd0}, _T_7470}; // @[Bitwise.scala 48:55:@5471.4]
  assign _T_7516 = _GEN_868 + _T_7515; // @[Bitwise.scala 48:55:@5471.4]
  assign _T_7517 = _T_7514 + _T_7516; // @[Bitwise.scala 48:55:@5472.4]
  assign _T_7518 = _T_7512 + _T_7517; // @[Bitwise.scala 48:55:@5473.4]
  assign _T_7519 = _T_7507 + _T_7518; // @[Bitwise.scala 48:55:@5474.4]
  assign _T_7520 = _T_7474 + _T_7475; // @[Bitwise.scala 48:55:@5475.4]
  assign _GEN_869 = {{1'd0}, _T_7473}; // @[Bitwise.scala 48:55:@5476.4]
  assign _T_7521 = _GEN_869 + _T_7520; // @[Bitwise.scala 48:55:@5476.4]
  assign _T_7522 = _T_7477 + _T_7478; // @[Bitwise.scala 48:55:@5477.4]
  assign _GEN_870 = {{1'd0}, _T_7476}; // @[Bitwise.scala 48:55:@5478.4]
  assign _T_7523 = _GEN_870 + _T_7522; // @[Bitwise.scala 48:55:@5478.4]
  assign _T_7524 = _T_7521 + _T_7523; // @[Bitwise.scala 48:55:@5479.4]
  assign _T_7525 = _T_7480 + _T_7481; // @[Bitwise.scala 48:55:@5480.4]
  assign _GEN_871 = {{1'd0}, _T_7479}; // @[Bitwise.scala 48:55:@5481.4]
  assign _T_7526 = _GEN_871 + _T_7525; // @[Bitwise.scala 48:55:@5481.4]
  assign _T_7527 = _T_7483 + _T_7484; // @[Bitwise.scala 48:55:@5482.4]
  assign _GEN_872 = {{1'd0}, _T_7482}; // @[Bitwise.scala 48:55:@5483.4]
  assign _T_7528 = _GEN_872 + _T_7527; // @[Bitwise.scala 48:55:@5483.4]
  assign _T_7529 = _T_7526 + _T_7528; // @[Bitwise.scala 48:55:@5484.4]
  assign _T_7530 = _T_7524 + _T_7529; // @[Bitwise.scala 48:55:@5485.4]
  assign _T_7531 = _T_7486 + _T_7487; // @[Bitwise.scala 48:55:@5486.4]
  assign _GEN_873 = {{1'd0}, _T_7485}; // @[Bitwise.scala 48:55:@5487.4]
  assign _T_7532 = _GEN_873 + _T_7531; // @[Bitwise.scala 48:55:@5487.4]
  assign _T_7533 = _T_7489 + _T_7490; // @[Bitwise.scala 48:55:@5488.4]
  assign _GEN_874 = {{1'd0}, _T_7488}; // @[Bitwise.scala 48:55:@5489.4]
  assign _T_7534 = _GEN_874 + _T_7533; // @[Bitwise.scala 48:55:@5489.4]
  assign _T_7535 = _T_7532 + _T_7534; // @[Bitwise.scala 48:55:@5490.4]
  assign _T_7536 = _T_7492 + _T_7493; // @[Bitwise.scala 48:55:@5491.4]
  assign _GEN_875 = {{1'd0}, _T_7491}; // @[Bitwise.scala 48:55:@5492.4]
  assign _T_7537 = _GEN_875 + _T_7536; // @[Bitwise.scala 48:55:@5492.4]
  assign _T_7538 = _T_7495 + _T_7496; // @[Bitwise.scala 48:55:@5493.4]
  assign _GEN_876 = {{1'd0}, _T_7494}; // @[Bitwise.scala 48:55:@5494.4]
  assign _T_7539 = _GEN_876 + _T_7538; // @[Bitwise.scala 48:55:@5494.4]
  assign _T_7540 = _T_7537 + _T_7539; // @[Bitwise.scala 48:55:@5495.4]
  assign _T_7541 = _T_7535 + _T_7540; // @[Bitwise.scala 48:55:@5496.4]
  assign _T_7542 = _T_7530 + _T_7541; // @[Bitwise.scala 48:55:@5497.4]
  assign _T_7543 = _T_7519 + _T_7542; // @[Bitwise.scala 48:55:@5498.4]
  assign _T_7607 = _T_2230[48:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5563.4]
  assign _T_7608 = _T_7607[0]; // @[Bitwise.scala 50:65:@5564.4]
  assign _T_7609 = _T_7607[1]; // @[Bitwise.scala 50:65:@5565.4]
  assign _T_7610 = _T_7607[2]; // @[Bitwise.scala 50:65:@5566.4]
  assign _T_7611 = _T_7607[3]; // @[Bitwise.scala 50:65:@5567.4]
  assign _T_7612 = _T_7607[4]; // @[Bitwise.scala 50:65:@5568.4]
  assign _T_7613 = _T_7607[5]; // @[Bitwise.scala 50:65:@5569.4]
  assign _T_7614 = _T_7607[6]; // @[Bitwise.scala 50:65:@5570.4]
  assign _T_7615 = _T_7607[7]; // @[Bitwise.scala 50:65:@5571.4]
  assign _T_7616 = _T_7607[8]; // @[Bitwise.scala 50:65:@5572.4]
  assign _T_7617 = _T_7607[9]; // @[Bitwise.scala 50:65:@5573.4]
  assign _T_7618 = _T_7607[10]; // @[Bitwise.scala 50:65:@5574.4]
  assign _T_7619 = _T_7607[11]; // @[Bitwise.scala 50:65:@5575.4]
  assign _T_7620 = _T_7607[12]; // @[Bitwise.scala 50:65:@5576.4]
  assign _T_7621 = _T_7607[13]; // @[Bitwise.scala 50:65:@5577.4]
  assign _T_7622 = _T_7607[14]; // @[Bitwise.scala 50:65:@5578.4]
  assign _T_7623 = _T_7607[15]; // @[Bitwise.scala 50:65:@5579.4]
  assign _T_7624 = _T_7607[16]; // @[Bitwise.scala 50:65:@5580.4]
  assign _T_7625 = _T_7607[17]; // @[Bitwise.scala 50:65:@5581.4]
  assign _T_7626 = _T_7607[18]; // @[Bitwise.scala 50:65:@5582.4]
  assign _T_7627 = _T_7607[19]; // @[Bitwise.scala 50:65:@5583.4]
  assign _T_7628 = _T_7607[20]; // @[Bitwise.scala 50:65:@5584.4]
  assign _T_7629 = _T_7607[21]; // @[Bitwise.scala 50:65:@5585.4]
  assign _T_7630 = _T_7607[22]; // @[Bitwise.scala 50:65:@5586.4]
  assign _T_7631 = _T_7607[23]; // @[Bitwise.scala 50:65:@5587.4]
  assign _T_7632 = _T_7607[24]; // @[Bitwise.scala 50:65:@5588.4]
  assign _T_7633 = _T_7607[25]; // @[Bitwise.scala 50:65:@5589.4]
  assign _T_7634 = _T_7607[26]; // @[Bitwise.scala 50:65:@5590.4]
  assign _T_7635 = _T_7607[27]; // @[Bitwise.scala 50:65:@5591.4]
  assign _T_7636 = _T_7607[28]; // @[Bitwise.scala 50:65:@5592.4]
  assign _T_7637 = _T_7607[29]; // @[Bitwise.scala 50:65:@5593.4]
  assign _T_7638 = _T_7607[30]; // @[Bitwise.scala 50:65:@5594.4]
  assign _T_7639 = _T_7607[31]; // @[Bitwise.scala 50:65:@5595.4]
  assign _T_7640 = _T_7607[32]; // @[Bitwise.scala 50:65:@5596.4]
  assign _T_7641 = _T_7607[33]; // @[Bitwise.scala 50:65:@5597.4]
  assign _T_7642 = _T_7607[34]; // @[Bitwise.scala 50:65:@5598.4]
  assign _T_7643 = _T_7607[35]; // @[Bitwise.scala 50:65:@5599.4]
  assign _T_7644 = _T_7607[36]; // @[Bitwise.scala 50:65:@5600.4]
  assign _T_7645 = _T_7607[37]; // @[Bitwise.scala 50:65:@5601.4]
  assign _T_7646 = _T_7607[38]; // @[Bitwise.scala 50:65:@5602.4]
  assign _T_7647 = _T_7607[39]; // @[Bitwise.scala 50:65:@5603.4]
  assign _T_7648 = _T_7607[40]; // @[Bitwise.scala 50:65:@5604.4]
  assign _T_7649 = _T_7607[41]; // @[Bitwise.scala 50:65:@5605.4]
  assign _T_7650 = _T_7607[42]; // @[Bitwise.scala 50:65:@5606.4]
  assign _T_7651 = _T_7607[43]; // @[Bitwise.scala 50:65:@5607.4]
  assign _T_7652 = _T_7607[44]; // @[Bitwise.scala 50:65:@5608.4]
  assign _T_7653 = _T_7607[45]; // @[Bitwise.scala 50:65:@5609.4]
  assign _T_7654 = _T_7607[46]; // @[Bitwise.scala 50:65:@5610.4]
  assign _T_7655 = _T_7607[47]; // @[Bitwise.scala 50:65:@5611.4]
  assign _T_7656 = _T_7607[48]; // @[Bitwise.scala 50:65:@5612.4]
  assign _T_7657 = _T_7609 + _T_7610; // @[Bitwise.scala 48:55:@5613.4]
  assign _GEN_877 = {{1'd0}, _T_7608}; // @[Bitwise.scala 48:55:@5614.4]
  assign _T_7658 = _GEN_877 + _T_7657; // @[Bitwise.scala 48:55:@5614.4]
  assign _T_7659 = _T_7612 + _T_7613; // @[Bitwise.scala 48:55:@5615.4]
  assign _GEN_878 = {{1'd0}, _T_7611}; // @[Bitwise.scala 48:55:@5616.4]
  assign _T_7660 = _GEN_878 + _T_7659; // @[Bitwise.scala 48:55:@5616.4]
  assign _T_7661 = _T_7658 + _T_7660; // @[Bitwise.scala 48:55:@5617.4]
  assign _T_7662 = _T_7615 + _T_7616; // @[Bitwise.scala 48:55:@5618.4]
  assign _GEN_879 = {{1'd0}, _T_7614}; // @[Bitwise.scala 48:55:@5619.4]
  assign _T_7663 = _GEN_879 + _T_7662; // @[Bitwise.scala 48:55:@5619.4]
  assign _T_7664 = _T_7618 + _T_7619; // @[Bitwise.scala 48:55:@5620.4]
  assign _GEN_880 = {{1'd0}, _T_7617}; // @[Bitwise.scala 48:55:@5621.4]
  assign _T_7665 = _GEN_880 + _T_7664; // @[Bitwise.scala 48:55:@5621.4]
  assign _T_7666 = _T_7663 + _T_7665; // @[Bitwise.scala 48:55:@5622.4]
  assign _T_7667 = _T_7661 + _T_7666; // @[Bitwise.scala 48:55:@5623.4]
  assign _T_7668 = _T_7621 + _T_7622; // @[Bitwise.scala 48:55:@5624.4]
  assign _GEN_881 = {{1'd0}, _T_7620}; // @[Bitwise.scala 48:55:@5625.4]
  assign _T_7669 = _GEN_881 + _T_7668; // @[Bitwise.scala 48:55:@5625.4]
  assign _T_7670 = _T_7624 + _T_7625; // @[Bitwise.scala 48:55:@5626.4]
  assign _GEN_882 = {{1'd0}, _T_7623}; // @[Bitwise.scala 48:55:@5627.4]
  assign _T_7671 = _GEN_882 + _T_7670; // @[Bitwise.scala 48:55:@5627.4]
  assign _T_7672 = _T_7669 + _T_7671; // @[Bitwise.scala 48:55:@5628.4]
  assign _T_7673 = _T_7627 + _T_7628; // @[Bitwise.scala 48:55:@5629.4]
  assign _GEN_883 = {{1'd0}, _T_7626}; // @[Bitwise.scala 48:55:@5630.4]
  assign _T_7674 = _GEN_883 + _T_7673; // @[Bitwise.scala 48:55:@5630.4]
  assign _T_7675 = _T_7630 + _T_7631; // @[Bitwise.scala 48:55:@5631.4]
  assign _GEN_884 = {{1'd0}, _T_7629}; // @[Bitwise.scala 48:55:@5632.4]
  assign _T_7676 = _GEN_884 + _T_7675; // @[Bitwise.scala 48:55:@5632.4]
  assign _T_7677 = _T_7674 + _T_7676; // @[Bitwise.scala 48:55:@5633.4]
  assign _T_7678 = _T_7672 + _T_7677; // @[Bitwise.scala 48:55:@5634.4]
  assign _T_7679 = _T_7667 + _T_7678; // @[Bitwise.scala 48:55:@5635.4]
  assign _T_7680 = _T_7633 + _T_7634; // @[Bitwise.scala 48:55:@5636.4]
  assign _GEN_885 = {{1'd0}, _T_7632}; // @[Bitwise.scala 48:55:@5637.4]
  assign _T_7681 = _GEN_885 + _T_7680; // @[Bitwise.scala 48:55:@5637.4]
  assign _T_7682 = _T_7636 + _T_7637; // @[Bitwise.scala 48:55:@5638.4]
  assign _GEN_886 = {{1'd0}, _T_7635}; // @[Bitwise.scala 48:55:@5639.4]
  assign _T_7683 = _GEN_886 + _T_7682; // @[Bitwise.scala 48:55:@5639.4]
  assign _T_7684 = _T_7681 + _T_7683; // @[Bitwise.scala 48:55:@5640.4]
  assign _T_7685 = _T_7639 + _T_7640; // @[Bitwise.scala 48:55:@5641.4]
  assign _GEN_887 = {{1'd0}, _T_7638}; // @[Bitwise.scala 48:55:@5642.4]
  assign _T_7686 = _GEN_887 + _T_7685; // @[Bitwise.scala 48:55:@5642.4]
  assign _T_7687 = _T_7642 + _T_7643; // @[Bitwise.scala 48:55:@5643.4]
  assign _GEN_888 = {{1'd0}, _T_7641}; // @[Bitwise.scala 48:55:@5644.4]
  assign _T_7688 = _GEN_888 + _T_7687; // @[Bitwise.scala 48:55:@5644.4]
  assign _T_7689 = _T_7686 + _T_7688; // @[Bitwise.scala 48:55:@5645.4]
  assign _T_7690 = _T_7684 + _T_7689; // @[Bitwise.scala 48:55:@5646.4]
  assign _T_7691 = _T_7645 + _T_7646; // @[Bitwise.scala 48:55:@5647.4]
  assign _GEN_889 = {{1'd0}, _T_7644}; // @[Bitwise.scala 48:55:@5648.4]
  assign _T_7692 = _GEN_889 + _T_7691; // @[Bitwise.scala 48:55:@5648.4]
  assign _T_7693 = _T_7648 + _T_7649; // @[Bitwise.scala 48:55:@5649.4]
  assign _GEN_890 = {{1'd0}, _T_7647}; // @[Bitwise.scala 48:55:@5650.4]
  assign _T_7694 = _GEN_890 + _T_7693; // @[Bitwise.scala 48:55:@5650.4]
  assign _T_7695 = _T_7692 + _T_7694; // @[Bitwise.scala 48:55:@5651.4]
  assign _T_7696 = _T_7651 + _T_7652; // @[Bitwise.scala 48:55:@5652.4]
  assign _GEN_891 = {{1'd0}, _T_7650}; // @[Bitwise.scala 48:55:@5653.4]
  assign _T_7697 = _GEN_891 + _T_7696; // @[Bitwise.scala 48:55:@5653.4]
  assign _T_7698 = _T_7653 + _T_7654; // @[Bitwise.scala 48:55:@5654.4]
  assign _T_7699 = _T_7655 + _T_7656; // @[Bitwise.scala 48:55:@5655.4]
  assign _T_7700 = _T_7698 + _T_7699; // @[Bitwise.scala 48:55:@5656.4]
  assign _T_7701 = _T_7697 + _T_7700; // @[Bitwise.scala 48:55:@5657.4]
  assign _T_7702 = _T_7695 + _T_7701; // @[Bitwise.scala 48:55:@5658.4]
  assign _T_7703 = _T_7690 + _T_7702; // @[Bitwise.scala 48:55:@5659.4]
  assign _T_7704 = _T_7679 + _T_7703; // @[Bitwise.scala 48:55:@5660.4]
  assign _T_7768 = _T_2230[49:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5725.4]
  assign _T_7769 = _T_7768[0]; // @[Bitwise.scala 50:65:@5726.4]
  assign _T_7770 = _T_7768[1]; // @[Bitwise.scala 50:65:@5727.4]
  assign _T_7771 = _T_7768[2]; // @[Bitwise.scala 50:65:@5728.4]
  assign _T_7772 = _T_7768[3]; // @[Bitwise.scala 50:65:@5729.4]
  assign _T_7773 = _T_7768[4]; // @[Bitwise.scala 50:65:@5730.4]
  assign _T_7774 = _T_7768[5]; // @[Bitwise.scala 50:65:@5731.4]
  assign _T_7775 = _T_7768[6]; // @[Bitwise.scala 50:65:@5732.4]
  assign _T_7776 = _T_7768[7]; // @[Bitwise.scala 50:65:@5733.4]
  assign _T_7777 = _T_7768[8]; // @[Bitwise.scala 50:65:@5734.4]
  assign _T_7778 = _T_7768[9]; // @[Bitwise.scala 50:65:@5735.4]
  assign _T_7779 = _T_7768[10]; // @[Bitwise.scala 50:65:@5736.4]
  assign _T_7780 = _T_7768[11]; // @[Bitwise.scala 50:65:@5737.4]
  assign _T_7781 = _T_7768[12]; // @[Bitwise.scala 50:65:@5738.4]
  assign _T_7782 = _T_7768[13]; // @[Bitwise.scala 50:65:@5739.4]
  assign _T_7783 = _T_7768[14]; // @[Bitwise.scala 50:65:@5740.4]
  assign _T_7784 = _T_7768[15]; // @[Bitwise.scala 50:65:@5741.4]
  assign _T_7785 = _T_7768[16]; // @[Bitwise.scala 50:65:@5742.4]
  assign _T_7786 = _T_7768[17]; // @[Bitwise.scala 50:65:@5743.4]
  assign _T_7787 = _T_7768[18]; // @[Bitwise.scala 50:65:@5744.4]
  assign _T_7788 = _T_7768[19]; // @[Bitwise.scala 50:65:@5745.4]
  assign _T_7789 = _T_7768[20]; // @[Bitwise.scala 50:65:@5746.4]
  assign _T_7790 = _T_7768[21]; // @[Bitwise.scala 50:65:@5747.4]
  assign _T_7791 = _T_7768[22]; // @[Bitwise.scala 50:65:@5748.4]
  assign _T_7792 = _T_7768[23]; // @[Bitwise.scala 50:65:@5749.4]
  assign _T_7793 = _T_7768[24]; // @[Bitwise.scala 50:65:@5750.4]
  assign _T_7794 = _T_7768[25]; // @[Bitwise.scala 50:65:@5751.4]
  assign _T_7795 = _T_7768[26]; // @[Bitwise.scala 50:65:@5752.4]
  assign _T_7796 = _T_7768[27]; // @[Bitwise.scala 50:65:@5753.4]
  assign _T_7797 = _T_7768[28]; // @[Bitwise.scala 50:65:@5754.4]
  assign _T_7798 = _T_7768[29]; // @[Bitwise.scala 50:65:@5755.4]
  assign _T_7799 = _T_7768[30]; // @[Bitwise.scala 50:65:@5756.4]
  assign _T_7800 = _T_7768[31]; // @[Bitwise.scala 50:65:@5757.4]
  assign _T_7801 = _T_7768[32]; // @[Bitwise.scala 50:65:@5758.4]
  assign _T_7802 = _T_7768[33]; // @[Bitwise.scala 50:65:@5759.4]
  assign _T_7803 = _T_7768[34]; // @[Bitwise.scala 50:65:@5760.4]
  assign _T_7804 = _T_7768[35]; // @[Bitwise.scala 50:65:@5761.4]
  assign _T_7805 = _T_7768[36]; // @[Bitwise.scala 50:65:@5762.4]
  assign _T_7806 = _T_7768[37]; // @[Bitwise.scala 50:65:@5763.4]
  assign _T_7807 = _T_7768[38]; // @[Bitwise.scala 50:65:@5764.4]
  assign _T_7808 = _T_7768[39]; // @[Bitwise.scala 50:65:@5765.4]
  assign _T_7809 = _T_7768[40]; // @[Bitwise.scala 50:65:@5766.4]
  assign _T_7810 = _T_7768[41]; // @[Bitwise.scala 50:65:@5767.4]
  assign _T_7811 = _T_7768[42]; // @[Bitwise.scala 50:65:@5768.4]
  assign _T_7812 = _T_7768[43]; // @[Bitwise.scala 50:65:@5769.4]
  assign _T_7813 = _T_7768[44]; // @[Bitwise.scala 50:65:@5770.4]
  assign _T_7814 = _T_7768[45]; // @[Bitwise.scala 50:65:@5771.4]
  assign _T_7815 = _T_7768[46]; // @[Bitwise.scala 50:65:@5772.4]
  assign _T_7816 = _T_7768[47]; // @[Bitwise.scala 50:65:@5773.4]
  assign _T_7817 = _T_7768[48]; // @[Bitwise.scala 50:65:@5774.4]
  assign _T_7818 = _T_7768[49]; // @[Bitwise.scala 50:65:@5775.4]
  assign _T_7819 = _T_7770 + _T_7771; // @[Bitwise.scala 48:55:@5776.4]
  assign _GEN_892 = {{1'd0}, _T_7769}; // @[Bitwise.scala 48:55:@5777.4]
  assign _T_7820 = _GEN_892 + _T_7819; // @[Bitwise.scala 48:55:@5777.4]
  assign _T_7821 = _T_7773 + _T_7774; // @[Bitwise.scala 48:55:@5778.4]
  assign _GEN_893 = {{1'd0}, _T_7772}; // @[Bitwise.scala 48:55:@5779.4]
  assign _T_7822 = _GEN_893 + _T_7821; // @[Bitwise.scala 48:55:@5779.4]
  assign _T_7823 = _T_7820 + _T_7822; // @[Bitwise.scala 48:55:@5780.4]
  assign _T_7824 = _T_7776 + _T_7777; // @[Bitwise.scala 48:55:@5781.4]
  assign _GEN_894 = {{1'd0}, _T_7775}; // @[Bitwise.scala 48:55:@5782.4]
  assign _T_7825 = _GEN_894 + _T_7824; // @[Bitwise.scala 48:55:@5782.4]
  assign _T_7826 = _T_7779 + _T_7780; // @[Bitwise.scala 48:55:@5783.4]
  assign _GEN_895 = {{1'd0}, _T_7778}; // @[Bitwise.scala 48:55:@5784.4]
  assign _T_7827 = _GEN_895 + _T_7826; // @[Bitwise.scala 48:55:@5784.4]
  assign _T_7828 = _T_7825 + _T_7827; // @[Bitwise.scala 48:55:@5785.4]
  assign _T_7829 = _T_7823 + _T_7828; // @[Bitwise.scala 48:55:@5786.4]
  assign _T_7830 = _T_7782 + _T_7783; // @[Bitwise.scala 48:55:@5787.4]
  assign _GEN_896 = {{1'd0}, _T_7781}; // @[Bitwise.scala 48:55:@5788.4]
  assign _T_7831 = _GEN_896 + _T_7830; // @[Bitwise.scala 48:55:@5788.4]
  assign _T_7832 = _T_7785 + _T_7786; // @[Bitwise.scala 48:55:@5789.4]
  assign _GEN_897 = {{1'd0}, _T_7784}; // @[Bitwise.scala 48:55:@5790.4]
  assign _T_7833 = _GEN_897 + _T_7832; // @[Bitwise.scala 48:55:@5790.4]
  assign _T_7834 = _T_7831 + _T_7833; // @[Bitwise.scala 48:55:@5791.4]
  assign _T_7835 = _T_7788 + _T_7789; // @[Bitwise.scala 48:55:@5792.4]
  assign _GEN_898 = {{1'd0}, _T_7787}; // @[Bitwise.scala 48:55:@5793.4]
  assign _T_7836 = _GEN_898 + _T_7835; // @[Bitwise.scala 48:55:@5793.4]
  assign _T_7837 = _T_7790 + _T_7791; // @[Bitwise.scala 48:55:@5794.4]
  assign _T_7838 = _T_7792 + _T_7793; // @[Bitwise.scala 48:55:@5795.4]
  assign _T_7839 = _T_7837 + _T_7838; // @[Bitwise.scala 48:55:@5796.4]
  assign _T_7840 = _T_7836 + _T_7839; // @[Bitwise.scala 48:55:@5797.4]
  assign _T_7841 = _T_7834 + _T_7840; // @[Bitwise.scala 48:55:@5798.4]
  assign _T_7842 = _T_7829 + _T_7841; // @[Bitwise.scala 48:55:@5799.4]
  assign _T_7843 = _T_7795 + _T_7796; // @[Bitwise.scala 48:55:@5800.4]
  assign _GEN_899 = {{1'd0}, _T_7794}; // @[Bitwise.scala 48:55:@5801.4]
  assign _T_7844 = _GEN_899 + _T_7843; // @[Bitwise.scala 48:55:@5801.4]
  assign _T_7845 = _T_7798 + _T_7799; // @[Bitwise.scala 48:55:@5802.4]
  assign _GEN_900 = {{1'd0}, _T_7797}; // @[Bitwise.scala 48:55:@5803.4]
  assign _T_7846 = _GEN_900 + _T_7845; // @[Bitwise.scala 48:55:@5803.4]
  assign _T_7847 = _T_7844 + _T_7846; // @[Bitwise.scala 48:55:@5804.4]
  assign _T_7848 = _T_7801 + _T_7802; // @[Bitwise.scala 48:55:@5805.4]
  assign _GEN_901 = {{1'd0}, _T_7800}; // @[Bitwise.scala 48:55:@5806.4]
  assign _T_7849 = _GEN_901 + _T_7848; // @[Bitwise.scala 48:55:@5806.4]
  assign _T_7850 = _T_7804 + _T_7805; // @[Bitwise.scala 48:55:@5807.4]
  assign _GEN_902 = {{1'd0}, _T_7803}; // @[Bitwise.scala 48:55:@5808.4]
  assign _T_7851 = _GEN_902 + _T_7850; // @[Bitwise.scala 48:55:@5808.4]
  assign _T_7852 = _T_7849 + _T_7851; // @[Bitwise.scala 48:55:@5809.4]
  assign _T_7853 = _T_7847 + _T_7852; // @[Bitwise.scala 48:55:@5810.4]
  assign _T_7854 = _T_7807 + _T_7808; // @[Bitwise.scala 48:55:@5811.4]
  assign _GEN_903 = {{1'd0}, _T_7806}; // @[Bitwise.scala 48:55:@5812.4]
  assign _T_7855 = _GEN_903 + _T_7854; // @[Bitwise.scala 48:55:@5812.4]
  assign _T_7856 = _T_7810 + _T_7811; // @[Bitwise.scala 48:55:@5813.4]
  assign _GEN_904 = {{1'd0}, _T_7809}; // @[Bitwise.scala 48:55:@5814.4]
  assign _T_7857 = _GEN_904 + _T_7856; // @[Bitwise.scala 48:55:@5814.4]
  assign _T_7858 = _T_7855 + _T_7857; // @[Bitwise.scala 48:55:@5815.4]
  assign _T_7859 = _T_7813 + _T_7814; // @[Bitwise.scala 48:55:@5816.4]
  assign _GEN_905 = {{1'd0}, _T_7812}; // @[Bitwise.scala 48:55:@5817.4]
  assign _T_7860 = _GEN_905 + _T_7859; // @[Bitwise.scala 48:55:@5817.4]
  assign _T_7861 = _T_7815 + _T_7816; // @[Bitwise.scala 48:55:@5818.4]
  assign _T_7862 = _T_7817 + _T_7818; // @[Bitwise.scala 48:55:@5819.4]
  assign _T_7863 = _T_7861 + _T_7862; // @[Bitwise.scala 48:55:@5820.4]
  assign _T_7864 = _T_7860 + _T_7863; // @[Bitwise.scala 48:55:@5821.4]
  assign _T_7865 = _T_7858 + _T_7864; // @[Bitwise.scala 48:55:@5822.4]
  assign _T_7866 = _T_7853 + _T_7865; // @[Bitwise.scala 48:55:@5823.4]
  assign _T_7867 = _T_7842 + _T_7866; // @[Bitwise.scala 48:55:@5824.4]
  assign _T_7931 = _T_2230[50:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@5889.4]
  assign _T_7932 = _T_7931[0]; // @[Bitwise.scala 50:65:@5890.4]
  assign _T_7933 = _T_7931[1]; // @[Bitwise.scala 50:65:@5891.4]
  assign _T_7934 = _T_7931[2]; // @[Bitwise.scala 50:65:@5892.4]
  assign _T_7935 = _T_7931[3]; // @[Bitwise.scala 50:65:@5893.4]
  assign _T_7936 = _T_7931[4]; // @[Bitwise.scala 50:65:@5894.4]
  assign _T_7937 = _T_7931[5]; // @[Bitwise.scala 50:65:@5895.4]
  assign _T_7938 = _T_7931[6]; // @[Bitwise.scala 50:65:@5896.4]
  assign _T_7939 = _T_7931[7]; // @[Bitwise.scala 50:65:@5897.4]
  assign _T_7940 = _T_7931[8]; // @[Bitwise.scala 50:65:@5898.4]
  assign _T_7941 = _T_7931[9]; // @[Bitwise.scala 50:65:@5899.4]
  assign _T_7942 = _T_7931[10]; // @[Bitwise.scala 50:65:@5900.4]
  assign _T_7943 = _T_7931[11]; // @[Bitwise.scala 50:65:@5901.4]
  assign _T_7944 = _T_7931[12]; // @[Bitwise.scala 50:65:@5902.4]
  assign _T_7945 = _T_7931[13]; // @[Bitwise.scala 50:65:@5903.4]
  assign _T_7946 = _T_7931[14]; // @[Bitwise.scala 50:65:@5904.4]
  assign _T_7947 = _T_7931[15]; // @[Bitwise.scala 50:65:@5905.4]
  assign _T_7948 = _T_7931[16]; // @[Bitwise.scala 50:65:@5906.4]
  assign _T_7949 = _T_7931[17]; // @[Bitwise.scala 50:65:@5907.4]
  assign _T_7950 = _T_7931[18]; // @[Bitwise.scala 50:65:@5908.4]
  assign _T_7951 = _T_7931[19]; // @[Bitwise.scala 50:65:@5909.4]
  assign _T_7952 = _T_7931[20]; // @[Bitwise.scala 50:65:@5910.4]
  assign _T_7953 = _T_7931[21]; // @[Bitwise.scala 50:65:@5911.4]
  assign _T_7954 = _T_7931[22]; // @[Bitwise.scala 50:65:@5912.4]
  assign _T_7955 = _T_7931[23]; // @[Bitwise.scala 50:65:@5913.4]
  assign _T_7956 = _T_7931[24]; // @[Bitwise.scala 50:65:@5914.4]
  assign _T_7957 = _T_7931[25]; // @[Bitwise.scala 50:65:@5915.4]
  assign _T_7958 = _T_7931[26]; // @[Bitwise.scala 50:65:@5916.4]
  assign _T_7959 = _T_7931[27]; // @[Bitwise.scala 50:65:@5917.4]
  assign _T_7960 = _T_7931[28]; // @[Bitwise.scala 50:65:@5918.4]
  assign _T_7961 = _T_7931[29]; // @[Bitwise.scala 50:65:@5919.4]
  assign _T_7962 = _T_7931[30]; // @[Bitwise.scala 50:65:@5920.4]
  assign _T_7963 = _T_7931[31]; // @[Bitwise.scala 50:65:@5921.4]
  assign _T_7964 = _T_7931[32]; // @[Bitwise.scala 50:65:@5922.4]
  assign _T_7965 = _T_7931[33]; // @[Bitwise.scala 50:65:@5923.4]
  assign _T_7966 = _T_7931[34]; // @[Bitwise.scala 50:65:@5924.4]
  assign _T_7967 = _T_7931[35]; // @[Bitwise.scala 50:65:@5925.4]
  assign _T_7968 = _T_7931[36]; // @[Bitwise.scala 50:65:@5926.4]
  assign _T_7969 = _T_7931[37]; // @[Bitwise.scala 50:65:@5927.4]
  assign _T_7970 = _T_7931[38]; // @[Bitwise.scala 50:65:@5928.4]
  assign _T_7971 = _T_7931[39]; // @[Bitwise.scala 50:65:@5929.4]
  assign _T_7972 = _T_7931[40]; // @[Bitwise.scala 50:65:@5930.4]
  assign _T_7973 = _T_7931[41]; // @[Bitwise.scala 50:65:@5931.4]
  assign _T_7974 = _T_7931[42]; // @[Bitwise.scala 50:65:@5932.4]
  assign _T_7975 = _T_7931[43]; // @[Bitwise.scala 50:65:@5933.4]
  assign _T_7976 = _T_7931[44]; // @[Bitwise.scala 50:65:@5934.4]
  assign _T_7977 = _T_7931[45]; // @[Bitwise.scala 50:65:@5935.4]
  assign _T_7978 = _T_7931[46]; // @[Bitwise.scala 50:65:@5936.4]
  assign _T_7979 = _T_7931[47]; // @[Bitwise.scala 50:65:@5937.4]
  assign _T_7980 = _T_7931[48]; // @[Bitwise.scala 50:65:@5938.4]
  assign _T_7981 = _T_7931[49]; // @[Bitwise.scala 50:65:@5939.4]
  assign _T_7982 = _T_7931[50]; // @[Bitwise.scala 50:65:@5940.4]
  assign _T_7983 = _T_7933 + _T_7934; // @[Bitwise.scala 48:55:@5941.4]
  assign _GEN_906 = {{1'd0}, _T_7932}; // @[Bitwise.scala 48:55:@5942.4]
  assign _T_7984 = _GEN_906 + _T_7983; // @[Bitwise.scala 48:55:@5942.4]
  assign _T_7985 = _T_7936 + _T_7937; // @[Bitwise.scala 48:55:@5943.4]
  assign _GEN_907 = {{1'd0}, _T_7935}; // @[Bitwise.scala 48:55:@5944.4]
  assign _T_7986 = _GEN_907 + _T_7985; // @[Bitwise.scala 48:55:@5944.4]
  assign _T_7987 = _T_7984 + _T_7986; // @[Bitwise.scala 48:55:@5945.4]
  assign _T_7988 = _T_7939 + _T_7940; // @[Bitwise.scala 48:55:@5946.4]
  assign _GEN_908 = {{1'd0}, _T_7938}; // @[Bitwise.scala 48:55:@5947.4]
  assign _T_7989 = _GEN_908 + _T_7988; // @[Bitwise.scala 48:55:@5947.4]
  assign _T_7990 = _T_7942 + _T_7943; // @[Bitwise.scala 48:55:@5948.4]
  assign _GEN_909 = {{1'd0}, _T_7941}; // @[Bitwise.scala 48:55:@5949.4]
  assign _T_7991 = _GEN_909 + _T_7990; // @[Bitwise.scala 48:55:@5949.4]
  assign _T_7992 = _T_7989 + _T_7991; // @[Bitwise.scala 48:55:@5950.4]
  assign _T_7993 = _T_7987 + _T_7992; // @[Bitwise.scala 48:55:@5951.4]
  assign _T_7994 = _T_7945 + _T_7946; // @[Bitwise.scala 48:55:@5952.4]
  assign _GEN_910 = {{1'd0}, _T_7944}; // @[Bitwise.scala 48:55:@5953.4]
  assign _T_7995 = _GEN_910 + _T_7994; // @[Bitwise.scala 48:55:@5953.4]
  assign _T_7996 = _T_7948 + _T_7949; // @[Bitwise.scala 48:55:@5954.4]
  assign _GEN_911 = {{1'd0}, _T_7947}; // @[Bitwise.scala 48:55:@5955.4]
  assign _T_7997 = _GEN_911 + _T_7996; // @[Bitwise.scala 48:55:@5955.4]
  assign _T_7998 = _T_7995 + _T_7997; // @[Bitwise.scala 48:55:@5956.4]
  assign _T_7999 = _T_7951 + _T_7952; // @[Bitwise.scala 48:55:@5957.4]
  assign _GEN_912 = {{1'd0}, _T_7950}; // @[Bitwise.scala 48:55:@5958.4]
  assign _T_8000 = _GEN_912 + _T_7999; // @[Bitwise.scala 48:55:@5958.4]
  assign _T_8001 = _T_7953 + _T_7954; // @[Bitwise.scala 48:55:@5959.4]
  assign _T_8002 = _T_7955 + _T_7956; // @[Bitwise.scala 48:55:@5960.4]
  assign _T_8003 = _T_8001 + _T_8002; // @[Bitwise.scala 48:55:@5961.4]
  assign _T_8004 = _T_8000 + _T_8003; // @[Bitwise.scala 48:55:@5962.4]
  assign _T_8005 = _T_7998 + _T_8004; // @[Bitwise.scala 48:55:@5963.4]
  assign _T_8006 = _T_7993 + _T_8005; // @[Bitwise.scala 48:55:@5964.4]
  assign _T_8007 = _T_7958 + _T_7959; // @[Bitwise.scala 48:55:@5965.4]
  assign _GEN_913 = {{1'd0}, _T_7957}; // @[Bitwise.scala 48:55:@5966.4]
  assign _T_8008 = _GEN_913 + _T_8007; // @[Bitwise.scala 48:55:@5966.4]
  assign _T_8009 = _T_7961 + _T_7962; // @[Bitwise.scala 48:55:@5967.4]
  assign _GEN_914 = {{1'd0}, _T_7960}; // @[Bitwise.scala 48:55:@5968.4]
  assign _T_8010 = _GEN_914 + _T_8009; // @[Bitwise.scala 48:55:@5968.4]
  assign _T_8011 = _T_8008 + _T_8010; // @[Bitwise.scala 48:55:@5969.4]
  assign _T_8012 = _T_7964 + _T_7965; // @[Bitwise.scala 48:55:@5970.4]
  assign _GEN_915 = {{1'd0}, _T_7963}; // @[Bitwise.scala 48:55:@5971.4]
  assign _T_8013 = _GEN_915 + _T_8012; // @[Bitwise.scala 48:55:@5971.4]
  assign _T_8014 = _T_7966 + _T_7967; // @[Bitwise.scala 48:55:@5972.4]
  assign _T_8015 = _T_7968 + _T_7969; // @[Bitwise.scala 48:55:@5973.4]
  assign _T_8016 = _T_8014 + _T_8015; // @[Bitwise.scala 48:55:@5974.4]
  assign _T_8017 = _T_8013 + _T_8016; // @[Bitwise.scala 48:55:@5975.4]
  assign _T_8018 = _T_8011 + _T_8017; // @[Bitwise.scala 48:55:@5976.4]
  assign _T_8019 = _T_7971 + _T_7972; // @[Bitwise.scala 48:55:@5977.4]
  assign _GEN_916 = {{1'd0}, _T_7970}; // @[Bitwise.scala 48:55:@5978.4]
  assign _T_8020 = _GEN_916 + _T_8019; // @[Bitwise.scala 48:55:@5978.4]
  assign _T_8021 = _T_7974 + _T_7975; // @[Bitwise.scala 48:55:@5979.4]
  assign _GEN_917 = {{1'd0}, _T_7973}; // @[Bitwise.scala 48:55:@5980.4]
  assign _T_8022 = _GEN_917 + _T_8021; // @[Bitwise.scala 48:55:@5980.4]
  assign _T_8023 = _T_8020 + _T_8022; // @[Bitwise.scala 48:55:@5981.4]
  assign _T_8024 = _T_7977 + _T_7978; // @[Bitwise.scala 48:55:@5982.4]
  assign _GEN_918 = {{1'd0}, _T_7976}; // @[Bitwise.scala 48:55:@5983.4]
  assign _T_8025 = _GEN_918 + _T_8024; // @[Bitwise.scala 48:55:@5983.4]
  assign _T_8026 = _T_7979 + _T_7980; // @[Bitwise.scala 48:55:@5984.4]
  assign _T_8027 = _T_7981 + _T_7982; // @[Bitwise.scala 48:55:@5985.4]
  assign _T_8028 = _T_8026 + _T_8027; // @[Bitwise.scala 48:55:@5986.4]
  assign _T_8029 = _T_8025 + _T_8028; // @[Bitwise.scala 48:55:@5987.4]
  assign _T_8030 = _T_8023 + _T_8029; // @[Bitwise.scala 48:55:@5988.4]
  assign _T_8031 = _T_8018 + _T_8030; // @[Bitwise.scala 48:55:@5989.4]
  assign _T_8032 = _T_8006 + _T_8031; // @[Bitwise.scala 48:55:@5990.4]
  assign _T_8096 = _T_2230[51:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6055.4]
  assign _T_8097 = _T_8096[0]; // @[Bitwise.scala 50:65:@6056.4]
  assign _T_8098 = _T_8096[1]; // @[Bitwise.scala 50:65:@6057.4]
  assign _T_8099 = _T_8096[2]; // @[Bitwise.scala 50:65:@6058.4]
  assign _T_8100 = _T_8096[3]; // @[Bitwise.scala 50:65:@6059.4]
  assign _T_8101 = _T_8096[4]; // @[Bitwise.scala 50:65:@6060.4]
  assign _T_8102 = _T_8096[5]; // @[Bitwise.scala 50:65:@6061.4]
  assign _T_8103 = _T_8096[6]; // @[Bitwise.scala 50:65:@6062.4]
  assign _T_8104 = _T_8096[7]; // @[Bitwise.scala 50:65:@6063.4]
  assign _T_8105 = _T_8096[8]; // @[Bitwise.scala 50:65:@6064.4]
  assign _T_8106 = _T_8096[9]; // @[Bitwise.scala 50:65:@6065.4]
  assign _T_8107 = _T_8096[10]; // @[Bitwise.scala 50:65:@6066.4]
  assign _T_8108 = _T_8096[11]; // @[Bitwise.scala 50:65:@6067.4]
  assign _T_8109 = _T_8096[12]; // @[Bitwise.scala 50:65:@6068.4]
  assign _T_8110 = _T_8096[13]; // @[Bitwise.scala 50:65:@6069.4]
  assign _T_8111 = _T_8096[14]; // @[Bitwise.scala 50:65:@6070.4]
  assign _T_8112 = _T_8096[15]; // @[Bitwise.scala 50:65:@6071.4]
  assign _T_8113 = _T_8096[16]; // @[Bitwise.scala 50:65:@6072.4]
  assign _T_8114 = _T_8096[17]; // @[Bitwise.scala 50:65:@6073.4]
  assign _T_8115 = _T_8096[18]; // @[Bitwise.scala 50:65:@6074.4]
  assign _T_8116 = _T_8096[19]; // @[Bitwise.scala 50:65:@6075.4]
  assign _T_8117 = _T_8096[20]; // @[Bitwise.scala 50:65:@6076.4]
  assign _T_8118 = _T_8096[21]; // @[Bitwise.scala 50:65:@6077.4]
  assign _T_8119 = _T_8096[22]; // @[Bitwise.scala 50:65:@6078.4]
  assign _T_8120 = _T_8096[23]; // @[Bitwise.scala 50:65:@6079.4]
  assign _T_8121 = _T_8096[24]; // @[Bitwise.scala 50:65:@6080.4]
  assign _T_8122 = _T_8096[25]; // @[Bitwise.scala 50:65:@6081.4]
  assign _T_8123 = _T_8096[26]; // @[Bitwise.scala 50:65:@6082.4]
  assign _T_8124 = _T_8096[27]; // @[Bitwise.scala 50:65:@6083.4]
  assign _T_8125 = _T_8096[28]; // @[Bitwise.scala 50:65:@6084.4]
  assign _T_8126 = _T_8096[29]; // @[Bitwise.scala 50:65:@6085.4]
  assign _T_8127 = _T_8096[30]; // @[Bitwise.scala 50:65:@6086.4]
  assign _T_8128 = _T_8096[31]; // @[Bitwise.scala 50:65:@6087.4]
  assign _T_8129 = _T_8096[32]; // @[Bitwise.scala 50:65:@6088.4]
  assign _T_8130 = _T_8096[33]; // @[Bitwise.scala 50:65:@6089.4]
  assign _T_8131 = _T_8096[34]; // @[Bitwise.scala 50:65:@6090.4]
  assign _T_8132 = _T_8096[35]; // @[Bitwise.scala 50:65:@6091.4]
  assign _T_8133 = _T_8096[36]; // @[Bitwise.scala 50:65:@6092.4]
  assign _T_8134 = _T_8096[37]; // @[Bitwise.scala 50:65:@6093.4]
  assign _T_8135 = _T_8096[38]; // @[Bitwise.scala 50:65:@6094.4]
  assign _T_8136 = _T_8096[39]; // @[Bitwise.scala 50:65:@6095.4]
  assign _T_8137 = _T_8096[40]; // @[Bitwise.scala 50:65:@6096.4]
  assign _T_8138 = _T_8096[41]; // @[Bitwise.scala 50:65:@6097.4]
  assign _T_8139 = _T_8096[42]; // @[Bitwise.scala 50:65:@6098.4]
  assign _T_8140 = _T_8096[43]; // @[Bitwise.scala 50:65:@6099.4]
  assign _T_8141 = _T_8096[44]; // @[Bitwise.scala 50:65:@6100.4]
  assign _T_8142 = _T_8096[45]; // @[Bitwise.scala 50:65:@6101.4]
  assign _T_8143 = _T_8096[46]; // @[Bitwise.scala 50:65:@6102.4]
  assign _T_8144 = _T_8096[47]; // @[Bitwise.scala 50:65:@6103.4]
  assign _T_8145 = _T_8096[48]; // @[Bitwise.scala 50:65:@6104.4]
  assign _T_8146 = _T_8096[49]; // @[Bitwise.scala 50:65:@6105.4]
  assign _T_8147 = _T_8096[50]; // @[Bitwise.scala 50:65:@6106.4]
  assign _T_8148 = _T_8096[51]; // @[Bitwise.scala 50:65:@6107.4]
  assign _T_8149 = _T_8098 + _T_8099; // @[Bitwise.scala 48:55:@6108.4]
  assign _GEN_919 = {{1'd0}, _T_8097}; // @[Bitwise.scala 48:55:@6109.4]
  assign _T_8150 = _GEN_919 + _T_8149; // @[Bitwise.scala 48:55:@6109.4]
  assign _T_8151 = _T_8101 + _T_8102; // @[Bitwise.scala 48:55:@6110.4]
  assign _GEN_920 = {{1'd0}, _T_8100}; // @[Bitwise.scala 48:55:@6111.4]
  assign _T_8152 = _GEN_920 + _T_8151; // @[Bitwise.scala 48:55:@6111.4]
  assign _T_8153 = _T_8150 + _T_8152; // @[Bitwise.scala 48:55:@6112.4]
  assign _T_8154 = _T_8104 + _T_8105; // @[Bitwise.scala 48:55:@6113.4]
  assign _GEN_921 = {{1'd0}, _T_8103}; // @[Bitwise.scala 48:55:@6114.4]
  assign _T_8155 = _GEN_921 + _T_8154; // @[Bitwise.scala 48:55:@6114.4]
  assign _T_8156 = _T_8106 + _T_8107; // @[Bitwise.scala 48:55:@6115.4]
  assign _T_8157 = _T_8108 + _T_8109; // @[Bitwise.scala 48:55:@6116.4]
  assign _T_8158 = _T_8156 + _T_8157; // @[Bitwise.scala 48:55:@6117.4]
  assign _T_8159 = _T_8155 + _T_8158; // @[Bitwise.scala 48:55:@6118.4]
  assign _T_8160 = _T_8153 + _T_8159; // @[Bitwise.scala 48:55:@6119.4]
  assign _T_8161 = _T_8111 + _T_8112; // @[Bitwise.scala 48:55:@6120.4]
  assign _GEN_922 = {{1'd0}, _T_8110}; // @[Bitwise.scala 48:55:@6121.4]
  assign _T_8162 = _GEN_922 + _T_8161; // @[Bitwise.scala 48:55:@6121.4]
  assign _T_8163 = _T_8114 + _T_8115; // @[Bitwise.scala 48:55:@6122.4]
  assign _GEN_923 = {{1'd0}, _T_8113}; // @[Bitwise.scala 48:55:@6123.4]
  assign _T_8164 = _GEN_923 + _T_8163; // @[Bitwise.scala 48:55:@6123.4]
  assign _T_8165 = _T_8162 + _T_8164; // @[Bitwise.scala 48:55:@6124.4]
  assign _T_8166 = _T_8117 + _T_8118; // @[Bitwise.scala 48:55:@6125.4]
  assign _GEN_924 = {{1'd0}, _T_8116}; // @[Bitwise.scala 48:55:@6126.4]
  assign _T_8167 = _GEN_924 + _T_8166; // @[Bitwise.scala 48:55:@6126.4]
  assign _T_8168 = _T_8119 + _T_8120; // @[Bitwise.scala 48:55:@6127.4]
  assign _T_8169 = _T_8121 + _T_8122; // @[Bitwise.scala 48:55:@6128.4]
  assign _T_8170 = _T_8168 + _T_8169; // @[Bitwise.scala 48:55:@6129.4]
  assign _T_8171 = _T_8167 + _T_8170; // @[Bitwise.scala 48:55:@6130.4]
  assign _T_8172 = _T_8165 + _T_8171; // @[Bitwise.scala 48:55:@6131.4]
  assign _T_8173 = _T_8160 + _T_8172; // @[Bitwise.scala 48:55:@6132.4]
  assign _T_8174 = _T_8124 + _T_8125; // @[Bitwise.scala 48:55:@6133.4]
  assign _GEN_925 = {{1'd0}, _T_8123}; // @[Bitwise.scala 48:55:@6134.4]
  assign _T_8175 = _GEN_925 + _T_8174; // @[Bitwise.scala 48:55:@6134.4]
  assign _T_8176 = _T_8127 + _T_8128; // @[Bitwise.scala 48:55:@6135.4]
  assign _GEN_926 = {{1'd0}, _T_8126}; // @[Bitwise.scala 48:55:@6136.4]
  assign _T_8177 = _GEN_926 + _T_8176; // @[Bitwise.scala 48:55:@6136.4]
  assign _T_8178 = _T_8175 + _T_8177; // @[Bitwise.scala 48:55:@6137.4]
  assign _T_8179 = _T_8130 + _T_8131; // @[Bitwise.scala 48:55:@6138.4]
  assign _GEN_927 = {{1'd0}, _T_8129}; // @[Bitwise.scala 48:55:@6139.4]
  assign _T_8180 = _GEN_927 + _T_8179; // @[Bitwise.scala 48:55:@6139.4]
  assign _T_8181 = _T_8132 + _T_8133; // @[Bitwise.scala 48:55:@6140.4]
  assign _T_8182 = _T_8134 + _T_8135; // @[Bitwise.scala 48:55:@6141.4]
  assign _T_8183 = _T_8181 + _T_8182; // @[Bitwise.scala 48:55:@6142.4]
  assign _T_8184 = _T_8180 + _T_8183; // @[Bitwise.scala 48:55:@6143.4]
  assign _T_8185 = _T_8178 + _T_8184; // @[Bitwise.scala 48:55:@6144.4]
  assign _T_8186 = _T_8137 + _T_8138; // @[Bitwise.scala 48:55:@6145.4]
  assign _GEN_928 = {{1'd0}, _T_8136}; // @[Bitwise.scala 48:55:@6146.4]
  assign _T_8187 = _GEN_928 + _T_8186; // @[Bitwise.scala 48:55:@6146.4]
  assign _T_8188 = _T_8140 + _T_8141; // @[Bitwise.scala 48:55:@6147.4]
  assign _GEN_929 = {{1'd0}, _T_8139}; // @[Bitwise.scala 48:55:@6148.4]
  assign _T_8189 = _GEN_929 + _T_8188; // @[Bitwise.scala 48:55:@6148.4]
  assign _T_8190 = _T_8187 + _T_8189; // @[Bitwise.scala 48:55:@6149.4]
  assign _T_8191 = _T_8143 + _T_8144; // @[Bitwise.scala 48:55:@6150.4]
  assign _GEN_930 = {{1'd0}, _T_8142}; // @[Bitwise.scala 48:55:@6151.4]
  assign _T_8192 = _GEN_930 + _T_8191; // @[Bitwise.scala 48:55:@6151.4]
  assign _T_8193 = _T_8145 + _T_8146; // @[Bitwise.scala 48:55:@6152.4]
  assign _T_8194 = _T_8147 + _T_8148; // @[Bitwise.scala 48:55:@6153.4]
  assign _T_8195 = _T_8193 + _T_8194; // @[Bitwise.scala 48:55:@6154.4]
  assign _T_8196 = _T_8192 + _T_8195; // @[Bitwise.scala 48:55:@6155.4]
  assign _T_8197 = _T_8190 + _T_8196; // @[Bitwise.scala 48:55:@6156.4]
  assign _T_8198 = _T_8185 + _T_8197; // @[Bitwise.scala 48:55:@6157.4]
  assign _T_8199 = _T_8173 + _T_8198; // @[Bitwise.scala 48:55:@6158.4]
  assign _T_8263 = _T_2230[52:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6223.4]
  assign _T_8264 = _T_8263[0]; // @[Bitwise.scala 50:65:@6224.4]
  assign _T_8265 = _T_8263[1]; // @[Bitwise.scala 50:65:@6225.4]
  assign _T_8266 = _T_8263[2]; // @[Bitwise.scala 50:65:@6226.4]
  assign _T_8267 = _T_8263[3]; // @[Bitwise.scala 50:65:@6227.4]
  assign _T_8268 = _T_8263[4]; // @[Bitwise.scala 50:65:@6228.4]
  assign _T_8269 = _T_8263[5]; // @[Bitwise.scala 50:65:@6229.4]
  assign _T_8270 = _T_8263[6]; // @[Bitwise.scala 50:65:@6230.4]
  assign _T_8271 = _T_8263[7]; // @[Bitwise.scala 50:65:@6231.4]
  assign _T_8272 = _T_8263[8]; // @[Bitwise.scala 50:65:@6232.4]
  assign _T_8273 = _T_8263[9]; // @[Bitwise.scala 50:65:@6233.4]
  assign _T_8274 = _T_8263[10]; // @[Bitwise.scala 50:65:@6234.4]
  assign _T_8275 = _T_8263[11]; // @[Bitwise.scala 50:65:@6235.4]
  assign _T_8276 = _T_8263[12]; // @[Bitwise.scala 50:65:@6236.4]
  assign _T_8277 = _T_8263[13]; // @[Bitwise.scala 50:65:@6237.4]
  assign _T_8278 = _T_8263[14]; // @[Bitwise.scala 50:65:@6238.4]
  assign _T_8279 = _T_8263[15]; // @[Bitwise.scala 50:65:@6239.4]
  assign _T_8280 = _T_8263[16]; // @[Bitwise.scala 50:65:@6240.4]
  assign _T_8281 = _T_8263[17]; // @[Bitwise.scala 50:65:@6241.4]
  assign _T_8282 = _T_8263[18]; // @[Bitwise.scala 50:65:@6242.4]
  assign _T_8283 = _T_8263[19]; // @[Bitwise.scala 50:65:@6243.4]
  assign _T_8284 = _T_8263[20]; // @[Bitwise.scala 50:65:@6244.4]
  assign _T_8285 = _T_8263[21]; // @[Bitwise.scala 50:65:@6245.4]
  assign _T_8286 = _T_8263[22]; // @[Bitwise.scala 50:65:@6246.4]
  assign _T_8287 = _T_8263[23]; // @[Bitwise.scala 50:65:@6247.4]
  assign _T_8288 = _T_8263[24]; // @[Bitwise.scala 50:65:@6248.4]
  assign _T_8289 = _T_8263[25]; // @[Bitwise.scala 50:65:@6249.4]
  assign _T_8290 = _T_8263[26]; // @[Bitwise.scala 50:65:@6250.4]
  assign _T_8291 = _T_8263[27]; // @[Bitwise.scala 50:65:@6251.4]
  assign _T_8292 = _T_8263[28]; // @[Bitwise.scala 50:65:@6252.4]
  assign _T_8293 = _T_8263[29]; // @[Bitwise.scala 50:65:@6253.4]
  assign _T_8294 = _T_8263[30]; // @[Bitwise.scala 50:65:@6254.4]
  assign _T_8295 = _T_8263[31]; // @[Bitwise.scala 50:65:@6255.4]
  assign _T_8296 = _T_8263[32]; // @[Bitwise.scala 50:65:@6256.4]
  assign _T_8297 = _T_8263[33]; // @[Bitwise.scala 50:65:@6257.4]
  assign _T_8298 = _T_8263[34]; // @[Bitwise.scala 50:65:@6258.4]
  assign _T_8299 = _T_8263[35]; // @[Bitwise.scala 50:65:@6259.4]
  assign _T_8300 = _T_8263[36]; // @[Bitwise.scala 50:65:@6260.4]
  assign _T_8301 = _T_8263[37]; // @[Bitwise.scala 50:65:@6261.4]
  assign _T_8302 = _T_8263[38]; // @[Bitwise.scala 50:65:@6262.4]
  assign _T_8303 = _T_8263[39]; // @[Bitwise.scala 50:65:@6263.4]
  assign _T_8304 = _T_8263[40]; // @[Bitwise.scala 50:65:@6264.4]
  assign _T_8305 = _T_8263[41]; // @[Bitwise.scala 50:65:@6265.4]
  assign _T_8306 = _T_8263[42]; // @[Bitwise.scala 50:65:@6266.4]
  assign _T_8307 = _T_8263[43]; // @[Bitwise.scala 50:65:@6267.4]
  assign _T_8308 = _T_8263[44]; // @[Bitwise.scala 50:65:@6268.4]
  assign _T_8309 = _T_8263[45]; // @[Bitwise.scala 50:65:@6269.4]
  assign _T_8310 = _T_8263[46]; // @[Bitwise.scala 50:65:@6270.4]
  assign _T_8311 = _T_8263[47]; // @[Bitwise.scala 50:65:@6271.4]
  assign _T_8312 = _T_8263[48]; // @[Bitwise.scala 50:65:@6272.4]
  assign _T_8313 = _T_8263[49]; // @[Bitwise.scala 50:65:@6273.4]
  assign _T_8314 = _T_8263[50]; // @[Bitwise.scala 50:65:@6274.4]
  assign _T_8315 = _T_8263[51]; // @[Bitwise.scala 50:65:@6275.4]
  assign _T_8316 = _T_8263[52]; // @[Bitwise.scala 50:65:@6276.4]
  assign _T_8317 = _T_8265 + _T_8266; // @[Bitwise.scala 48:55:@6277.4]
  assign _GEN_931 = {{1'd0}, _T_8264}; // @[Bitwise.scala 48:55:@6278.4]
  assign _T_8318 = _GEN_931 + _T_8317; // @[Bitwise.scala 48:55:@6278.4]
  assign _T_8319 = _T_8268 + _T_8269; // @[Bitwise.scala 48:55:@6279.4]
  assign _GEN_932 = {{1'd0}, _T_8267}; // @[Bitwise.scala 48:55:@6280.4]
  assign _T_8320 = _GEN_932 + _T_8319; // @[Bitwise.scala 48:55:@6280.4]
  assign _T_8321 = _T_8318 + _T_8320; // @[Bitwise.scala 48:55:@6281.4]
  assign _T_8322 = _T_8271 + _T_8272; // @[Bitwise.scala 48:55:@6282.4]
  assign _GEN_933 = {{1'd0}, _T_8270}; // @[Bitwise.scala 48:55:@6283.4]
  assign _T_8323 = _GEN_933 + _T_8322; // @[Bitwise.scala 48:55:@6283.4]
  assign _T_8324 = _T_8273 + _T_8274; // @[Bitwise.scala 48:55:@6284.4]
  assign _T_8325 = _T_8275 + _T_8276; // @[Bitwise.scala 48:55:@6285.4]
  assign _T_8326 = _T_8324 + _T_8325; // @[Bitwise.scala 48:55:@6286.4]
  assign _T_8327 = _T_8323 + _T_8326; // @[Bitwise.scala 48:55:@6287.4]
  assign _T_8328 = _T_8321 + _T_8327; // @[Bitwise.scala 48:55:@6288.4]
  assign _T_8329 = _T_8278 + _T_8279; // @[Bitwise.scala 48:55:@6289.4]
  assign _GEN_934 = {{1'd0}, _T_8277}; // @[Bitwise.scala 48:55:@6290.4]
  assign _T_8330 = _GEN_934 + _T_8329; // @[Bitwise.scala 48:55:@6290.4]
  assign _T_8331 = _T_8281 + _T_8282; // @[Bitwise.scala 48:55:@6291.4]
  assign _GEN_935 = {{1'd0}, _T_8280}; // @[Bitwise.scala 48:55:@6292.4]
  assign _T_8332 = _GEN_935 + _T_8331; // @[Bitwise.scala 48:55:@6292.4]
  assign _T_8333 = _T_8330 + _T_8332; // @[Bitwise.scala 48:55:@6293.4]
  assign _T_8334 = _T_8284 + _T_8285; // @[Bitwise.scala 48:55:@6294.4]
  assign _GEN_936 = {{1'd0}, _T_8283}; // @[Bitwise.scala 48:55:@6295.4]
  assign _T_8335 = _GEN_936 + _T_8334; // @[Bitwise.scala 48:55:@6295.4]
  assign _T_8336 = _T_8286 + _T_8287; // @[Bitwise.scala 48:55:@6296.4]
  assign _T_8337 = _T_8288 + _T_8289; // @[Bitwise.scala 48:55:@6297.4]
  assign _T_8338 = _T_8336 + _T_8337; // @[Bitwise.scala 48:55:@6298.4]
  assign _T_8339 = _T_8335 + _T_8338; // @[Bitwise.scala 48:55:@6299.4]
  assign _T_8340 = _T_8333 + _T_8339; // @[Bitwise.scala 48:55:@6300.4]
  assign _T_8341 = _T_8328 + _T_8340; // @[Bitwise.scala 48:55:@6301.4]
  assign _T_8342 = _T_8291 + _T_8292; // @[Bitwise.scala 48:55:@6302.4]
  assign _GEN_937 = {{1'd0}, _T_8290}; // @[Bitwise.scala 48:55:@6303.4]
  assign _T_8343 = _GEN_937 + _T_8342; // @[Bitwise.scala 48:55:@6303.4]
  assign _T_8344 = _T_8294 + _T_8295; // @[Bitwise.scala 48:55:@6304.4]
  assign _GEN_938 = {{1'd0}, _T_8293}; // @[Bitwise.scala 48:55:@6305.4]
  assign _T_8345 = _GEN_938 + _T_8344; // @[Bitwise.scala 48:55:@6305.4]
  assign _T_8346 = _T_8343 + _T_8345; // @[Bitwise.scala 48:55:@6306.4]
  assign _T_8347 = _T_8297 + _T_8298; // @[Bitwise.scala 48:55:@6307.4]
  assign _GEN_939 = {{1'd0}, _T_8296}; // @[Bitwise.scala 48:55:@6308.4]
  assign _T_8348 = _GEN_939 + _T_8347; // @[Bitwise.scala 48:55:@6308.4]
  assign _T_8349 = _T_8299 + _T_8300; // @[Bitwise.scala 48:55:@6309.4]
  assign _T_8350 = _T_8301 + _T_8302; // @[Bitwise.scala 48:55:@6310.4]
  assign _T_8351 = _T_8349 + _T_8350; // @[Bitwise.scala 48:55:@6311.4]
  assign _T_8352 = _T_8348 + _T_8351; // @[Bitwise.scala 48:55:@6312.4]
  assign _T_8353 = _T_8346 + _T_8352; // @[Bitwise.scala 48:55:@6313.4]
  assign _T_8354 = _T_8304 + _T_8305; // @[Bitwise.scala 48:55:@6314.4]
  assign _GEN_940 = {{1'd0}, _T_8303}; // @[Bitwise.scala 48:55:@6315.4]
  assign _T_8355 = _GEN_940 + _T_8354; // @[Bitwise.scala 48:55:@6315.4]
  assign _T_8356 = _T_8306 + _T_8307; // @[Bitwise.scala 48:55:@6316.4]
  assign _T_8357 = _T_8308 + _T_8309; // @[Bitwise.scala 48:55:@6317.4]
  assign _T_8358 = _T_8356 + _T_8357; // @[Bitwise.scala 48:55:@6318.4]
  assign _T_8359 = _T_8355 + _T_8358; // @[Bitwise.scala 48:55:@6319.4]
  assign _T_8360 = _T_8311 + _T_8312; // @[Bitwise.scala 48:55:@6320.4]
  assign _GEN_941 = {{1'd0}, _T_8310}; // @[Bitwise.scala 48:55:@6321.4]
  assign _T_8361 = _GEN_941 + _T_8360; // @[Bitwise.scala 48:55:@6321.4]
  assign _T_8362 = _T_8313 + _T_8314; // @[Bitwise.scala 48:55:@6322.4]
  assign _T_8363 = _T_8315 + _T_8316; // @[Bitwise.scala 48:55:@6323.4]
  assign _T_8364 = _T_8362 + _T_8363; // @[Bitwise.scala 48:55:@6324.4]
  assign _T_8365 = _T_8361 + _T_8364; // @[Bitwise.scala 48:55:@6325.4]
  assign _T_8366 = _T_8359 + _T_8365; // @[Bitwise.scala 48:55:@6326.4]
  assign _T_8367 = _T_8353 + _T_8366; // @[Bitwise.scala 48:55:@6327.4]
  assign _T_8368 = _T_8341 + _T_8367; // @[Bitwise.scala 48:55:@6328.4]
  assign _T_8432 = _T_2230[53:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6393.4]
  assign _T_8433 = _T_8432[0]; // @[Bitwise.scala 50:65:@6394.4]
  assign _T_8434 = _T_8432[1]; // @[Bitwise.scala 50:65:@6395.4]
  assign _T_8435 = _T_8432[2]; // @[Bitwise.scala 50:65:@6396.4]
  assign _T_8436 = _T_8432[3]; // @[Bitwise.scala 50:65:@6397.4]
  assign _T_8437 = _T_8432[4]; // @[Bitwise.scala 50:65:@6398.4]
  assign _T_8438 = _T_8432[5]; // @[Bitwise.scala 50:65:@6399.4]
  assign _T_8439 = _T_8432[6]; // @[Bitwise.scala 50:65:@6400.4]
  assign _T_8440 = _T_8432[7]; // @[Bitwise.scala 50:65:@6401.4]
  assign _T_8441 = _T_8432[8]; // @[Bitwise.scala 50:65:@6402.4]
  assign _T_8442 = _T_8432[9]; // @[Bitwise.scala 50:65:@6403.4]
  assign _T_8443 = _T_8432[10]; // @[Bitwise.scala 50:65:@6404.4]
  assign _T_8444 = _T_8432[11]; // @[Bitwise.scala 50:65:@6405.4]
  assign _T_8445 = _T_8432[12]; // @[Bitwise.scala 50:65:@6406.4]
  assign _T_8446 = _T_8432[13]; // @[Bitwise.scala 50:65:@6407.4]
  assign _T_8447 = _T_8432[14]; // @[Bitwise.scala 50:65:@6408.4]
  assign _T_8448 = _T_8432[15]; // @[Bitwise.scala 50:65:@6409.4]
  assign _T_8449 = _T_8432[16]; // @[Bitwise.scala 50:65:@6410.4]
  assign _T_8450 = _T_8432[17]; // @[Bitwise.scala 50:65:@6411.4]
  assign _T_8451 = _T_8432[18]; // @[Bitwise.scala 50:65:@6412.4]
  assign _T_8452 = _T_8432[19]; // @[Bitwise.scala 50:65:@6413.4]
  assign _T_8453 = _T_8432[20]; // @[Bitwise.scala 50:65:@6414.4]
  assign _T_8454 = _T_8432[21]; // @[Bitwise.scala 50:65:@6415.4]
  assign _T_8455 = _T_8432[22]; // @[Bitwise.scala 50:65:@6416.4]
  assign _T_8456 = _T_8432[23]; // @[Bitwise.scala 50:65:@6417.4]
  assign _T_8457 = _T_8432[24]; // @[Bitwise.scala 50:65:@6418.4]
  assign _T_8458 = _T_8432[25]; // @[Bitwise.scala 50:65:@6419.4]
  assign _T_8459 = _T_8432[26]; // @[Bitwise.scala 50:65:@6420.4]
  assign _T_8460 = _T_8432[27]; // @[Bitwise.scala 50:65:@6421.4]
  assign _T_8461 = _T_8432[28]; // @[Bitwise.scala 50:65:@6422.4]
  assign _T_8462 = _T_8432[29]; // @[Bitwise.scala 50:65:@6423.4]
  assign _T_8463 = _T_8432[30]; // @[Bitwise.scala 50:65:@6424.4]
  assign _T_8464 = _T_8432[31]; // @[Bitwise.scala 50:65:@6425.4]
  assign _T_8465 = _T_8432[32]; // @[Bitwise.scala 50:65:@6426.4]
  assign _T_8466 = _T_8432[33]; // @[Bitwise.scala 50:65:@6427.4]
  assign _T_8467 = _T_8432[34]; // @[Bitwise.scala 50:65:@6428.4]
  assign _T_8468 = _T_8432[35]; // @[Bitwise.scala 50:65:@6429.4]
  assign _T_8469 = _T_8432[36]; // @[Bitwise.scala 50:65:@6430.4]
  assign _T_8470 = _T_8432[37]; // @[Bitwise.scala 50:65:@6431.4]
  assign _T_8471 = _T_8432[38]; // @[Bitwise.scala 50:65:@6432.4]
  assign _T_8472 = _T_8432[39]; // @[Bitwise.scala 50:65:@6433.4]
  assign _T_8473 = _T_8432[40]; // @[Bitwise.scala 50:65:@6434.4]
  assign _T_8474 = _T_8432[41]; // @[Bitwise.scala 50:65:@6435.4]
  assign _T_8475 = _T_8432[42]; // @[Bitwise.scala 50:65:@6436.4]
  assign _T_8476 = _T_8432[43]; // @[Bitwise.scala 50:65:@6437.4]
  assign _T_8477 = _T_8432[44]; // @[Bitwise.scala 50:65:@6438.4]
  assign _T_8478 = _T_8432[45]; // @[Bitwise.scala 50:65:@6439.4]
  assign _T_8479 = _T_8432[46]; // @[Bitwise.scala 50:65:@6440.4]
  assign _T_8480 = _T_8432[47]; // @[Bitwise.scala 50:65:@6441.4]
  assign _T_8481 = _T_8432[48]; // @[Bitwise.scala 50:65:@6442.4]
  assign _T_8482 = _T_8432[49]; // @[Bitwise.scala 50:65:@6443.4]
  assign _T_8483 = _T_8432[50]; // @[Bitwise.scala 50:65:@6444.4]
  assign _T_8484 = _T_8432[51]; // @[Bitwise.scala 50:65:@6445.4]
  assign _T_8485 = _T_8432[52]; // @[Bitwise.scala 50:65:@6446.4]
  assign _T_8486 = _T_8432[53]; // @[Bitwise.scala 50:65:@6447.4]
  assign _T_8487 = _T_8434 + _T_8435; // @[Bitwise.scala 48:55:@6448.4]
  assign _GEN_942 = {{1'd0}, _T_8433}; // @[Bitwise.scala 48:55:@6449.4]
  assign _T_8488 = _GEN_942 + _T_8487; // @[Bitwise.scala 48:55:@6449.4]
  assign _T_8489 = _T_8437 + _T_8438; // @[Bitwise.scala 48:55:@6450.4]
  assign _GEN_943 = {{1'd0}, _T_8436}; // @[Bitwise.scala 48:55:@6451.4]
  assign _T_8490 = _GEN_943 + _T_8489; // @[Bitwise.scala 48:55:@6451.4]
  assign _T_8491 = _T_8488 + _T_8490; // @[Bitwise.scala 48:55:@6452.4]
  assign _T_8492 = _T_8440 + _T_8441; // @[Bitwise.scala 48:55:@6453.4]
  assign _GEN_944 = {{1'd0}, _T_8439}; // @[Bitwise.scala 48:55:@6454.4]
  assign _T_8493 = _GEN_944 + _T_8492; // @[Bitwise.scala 48:55:@6454.4]
  assign _T_8494 = _T_8442 + _T_8443; // @[Bitwise.scala 48:55:@6455.4]
  assign _T_8495 = _T_8444 + _T_8445; // @[Bitwise.scala 48:55:@6456.4]
  assign _T_8496 = _T_8494 + _T_8495; // @[Bitwise.scala 48:55:@6457.4]
  assign _T_8497 = _T_8493 + _T_8496; // @[Bitwise.scala 48:55:@6458.4]
  assign _T_8498 = _T_8491 + _T_8497; // @[Bitwise.scala 48:55:@6459.4]
  assign _T_8499 = _T_8447 + _T_8448; // @[Bitwise.scala 48:55:@6460.4]
  assign _GEN_945 = {{1'd0}, _T_8446}; // @[Bitwise.scala 48:55:@6461.4]
  assign _T_8500 = _GEN_945 + _T_8499; // @[Bitwise.scala 48:55:@6461.4]
  assign _T_8501 = _T_8449 + _T_8450; // @[Bitwise.scala 48:55:@6462.4]
  assign _T_8502 = _T_8451 + _T_8452; // @[Bitwise.scala 48:55:@6463.4]
  assign _T_8503 = _T_8501 + _T_8502; // @[Bitwise.scala 48:55:@6464.4]
  assign _T_8504 = _T_8500 + _T_8503; // @[Bitwise.scala 48:55:@6465.4]
  assign _T_8505 = _T_8454 + _T_8455; // @[Bitwise.scala 48:55:@6466.4]
  assign _GEN_946 = {{1'd0}, _T_8453}; // @[Bitwise.scala 48:55:@6467.4]
  assign _T_8506 = _GEN_946 + _T_8505; // @[Bitwise.scala 48:55:@6467.4]
  assign _T_8507 = _T_8456 + _T_8457; // @[Bitwise.scala 48:55:@6468.4]
  assign _T_8508 = _T_8458 + _T_8459; // @[Bitwise.scala 48:55:@6469.4]
  assign _T_8509 = _T_8507 + _T_8508; // @[Bitwise.scala 48:55:@6470.4]
  assign _T_8510 = _T_8506 + _T_8509; // @[Bitwise.scala 48:55:@6471.4]
  assign _T_8511 = _T_8504 + _T_8510; // @[Bitwise.scala 48:55:@6472.4]
  assign _T_8512 = _T_8498 + _T_8511; // @[Bitwise.scala 48:55:@6473.4]
  assign _T_8513 = _T_8461 + _T_8462; // @[Bitwise.scala 48:55:@6474.4]
  assign _GEN_947 = {{1'd0}, _T_8460}; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_8514 = _GEN_947 + _T_8513; // @[Bitwise.scala 48:55:@6475.4]
  assign _T_8515 = _T_8464 + _T_8465; // @[Bitwise.scala 48:55:@6476.4]
  assign _GEN_948 = {{1'd0}, _T_8463}; // @[Bitwise.scala 48:55:@6477.4]
  assign _T_8516 = _GEN_948 + _T_8515; // @[Bitwise.scala 48:55:@6477.4]
  assign _T_8517 = _T_8514 + _T_8516; // @[Bitwise.scala 48:55:@6478.4]
  assign _T_8518 = _T_8467 + _T_8468; // @[Bitwise.scala 48:55:@6479.4]
  assign _GEN_949 = {{1'd0}, _T_8466}; // @[Bitwise.scala 48:55:@6480.4]
  assign _T_8519 = _GEN_949 + _T_8518; // @[Bitwise.scala 48:55:@6480.4]
  assign _T_8520 = _T_8469 + _T_8470; // @[Bitwise.scala 48:55:@6481.4]
  assign _T_8521 = _T_8471 + _T_8472; // @[Bitwise.scala 48:55:@6482.4]
  assign _T_8522 = _T_8520 + _T_8521; // @[Bitwise.scala 48:55:@6483.4]
  assign _T_8523 = _T_8519 + _T_8522; // @[Bitwise.scala 48:55:@6484.4]
  assign _T_8524 = _T_8517 + _T_8523; // @[Bitwise.scala 48:55:@6485.4]
  assign _T_8525 = _T_8474 + _T_8475; // @[Bitwise.scala 48:55:@6486.4]
  assign _GEN_950 = {{1'd0}, _T_8473}; // @[Bitwise.scala 48:55:@6487.4]
  assign _T_8526 = _GEN_950 + _T_8525; // @[Bitwise.scala 48:55:@6487.4]
  assign _T_8527 = _T_8476 + _T_8477; // @[Bitwise.scala 48:55:@6488.4]
  assign _T_8528 = _T_8478 + _T_8479; // @[Bitwise.scala 48:55:@6489.4]
  assign _T_8529 = _T_8527 + _T_8528; // @[Bitwise.scala 48:55:@6490.4]
  assign _T_8530 = _T_8526 + _T_8529; // @[Bitwise.scala 48:55:@6491.4]
  assign _T_8531 = _T_8481 + _T_8482; // @[Bitwise.scala 48:55:@6492.4]
  assign _GEN_951 = {{1'd0}, _T_8480}; // @[Bitwise.scala 48:55:@6493.4]
  assign _T_8532 = _GEN_951 + _T_8531; // @[Bitwise.scala 48:55:@6493.4]
  assign _T_8533 = _T_8483 + _T_8484; // @[Bitwise.scala 48:55:@6494.4]
  assign _T_8534 = _T_8485 + _T_8486; // @[Bitwise.scala 48:55:@6495.4]
  assign _T_8535 = _T_8533 + _T_8534; // @[Bitwise.scala 48:55:@6496.4]
  assign _T_8536 = _T_8532 + _T_8535; // @[Bitwise.scala 48:55:@6497.4]
  assign _T_8537 = _T_8530 + _T_8536; // @[Bitwise.scala 48:55:@6498.4]
  assign _T_8538 = _T_8524 + _T_8537; // @[Bitwise.scala 48:55:@6499.4]
  assign _T_8539 = _T_8512 + _T_8538; // @[Bitwise.scala 48:55:@6500.4]
  assign _T_8603 = _T_2230[54:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6565.4]
  assign _T_8604 = _T_8603[0]; // @[Bitwise.scala 50:65:@6566.4]
  assign _T_8605 = _T_8603[1]; // @[Bitwise.scala 50:65:@6567.4]
  assign _T_8606 = _T_8603[2]; // @[Bitwise.scala 50:65:@6568.4]
  assign _T_8607 = _T_8603[3]; // @[Bitwise.scala 50:65:@6569.4]
  assign _T_8608 = _T_8603[4]; // @[Bitwise.scala 50:65:@6570.4]
  assign _T_8609 = _T_8603[5]; // @[Bitwise.scala 50:65:@6571.4]
  assign _T_8610 = _T_8603[6]; // @[Bitwise.scala 50:65:@6572.4]
  assign _T_8611 = _T_8603[7]; // @[Bitwise.scala 50:65:@6573.4]
  assign _T_8612 = _T_8603[8]; // @[Bitwise.scala 50:65:@6574.4]
  assign _T_8613 = _T_8603[9]; // @[Bitwise.scala 50:65:@6575.4]
  assign _T_8614 = _T_8603[10]; // @[Bitwise.scala 50:65:@6576.4]
  assign _T_8615 = _T_8603[11]; // @[Bitwise.scala 50:65:@6577.4]
  assign _T_8616 = _T_8603[12]; // @[Bitwise.scala 50:65:@6578.4]
  assign _T_8617 = _T_8603[13]; // @[Bitwise.scala 50:65:@6579.4]
  assign _T_8618 = _T_8603[14]; // @[Bitwise.scala 50:65:@6580.4]
  assign _T_8619 = _T_8603[15]; // @[Bitwise.scala 50:65:@6581.4]
  assign _T_8620 = _T_8603[16]; // @[Bitwise.scala 50:65:@6582.4]
  assign _T_8621 = _T_8603[17]; // @[Bitwise.scala 50:65:@6583.4]
  assign _T_8622 = _T_8603[18]; // @[Bitwise.scala 50:65:@6584.4]
  assign _T_8623 = _T_8603[19]; // @[Bitwise.scala 50:65:@6585.4]
  assign _T_8624 = _T_8603[20]; // @[Bitwise.scala 50:65:@6586.4]
  assign _T_8625 = _T_8603[21]; // @[Bitwise.scala 50:65:@6587.4]
  assign _T_8626 = _T_8603[22]; // @[Bitwise.scala 50:65:@6588.4]
  assign _T_8627 = _T_8603[23]; // @[Bitwise.scala 50:65:@6589.4]
  assign _T_8628 = _T_8603[24]; // @[Bitwise.scala 50:65:@6590.4]
  assign _T_8629 = _T_8603[25]; // @[Bitwise.scala 50:65:@6591.4]
  assign _T_8630 = _T_8603[26]; // @[Bitwise.scala 50:65:@6592.4]
  assign _T_8631 = _T_8603[27]; // @[Bitwise.scala 50:65:@6593.4]
  assign _T_8632 = _T_8603[28]; // @[Bitwise.scala 50:65:@6594.4]
  assign _T_8633 = _T_8603[29]; // @[Bitwise.scala 50:65:@6595.4]
  assign _T_8634 = _T_8603[30]; // @[Bitwise.scala 50:65:@6596.4]
  assign _T_8635 = _T_8603[31]; // @[Bitwise.scala 50:65:@6597.4]
  assign _T_8636 = _T_8603[32]; // @[Bitwise.scala 50:65:@6598.4]
  assign _T_8637 = _T_8603[33]; // @[Bitwise.scala 50:65:@6599.4]
  assign _T_8638 = _T_8603[34]; // @[Bitwise.scala 50:65:@6600.4]
  assign _T_8639 = _T_8603[35]; // @[Bitwise.scala 50:65:@6601.4]
  assign _T_8640 = _T_8603[36]; // @[Bitwise.scala 50:65:@6602.4]
  assign _T_8641 = _T_8603[37]; // @[Bitwise.scala 50:65:@6603.4]
  assign _T_8642 = _T_8603[38]; // @[Bitwise.scala 50:65:@6604.4]
  assign _T_8643 = _T_8603[39]; // @[Bitwise.scala 50:65:@6605.4]
  assign _T_8644 = _T_8603[40]; // @[Bitwise.scala 50:65:@6606.4]
  assign _T_8645 = _T_8603[41]; // @[Bitwise.scala 50:65:@6607.4]
  assign _T_8646 = _T_8603[42]; // @[Bitwise.scala 50:65:@6608.4]
  assign _T_8647 = _T_8603[43]; // @[Bitwise.scala 50:65:@6609.4]
  assign _T_8648 = _T_8603[44]; // @[Bitwise.scala 50:65:@6610.4]
  assign _T_8649 = _T_8603[45]; // @[Bitwise.scala 50:65:@6611.4]
  assign _T_8650 = _T_8603[46]; // @[Bitwise.scala 50:65:@6612.4]
  assign _T_8651 = _T_8603[47]; // @[Bitwise.scala 50:65:@6613.4]
  assign _T_8652 = _T_8603[48]; // @[Bitwise.scala 50:65:@6614.4]
  assign _T_8653 = _T_8603[49]; // @[Bitwise.scala 50:65:@6615.4]
  assign _T_8654 = _T_8603[50]; // @[Bitwise.scala 50:65:@6616.4]
  assign _T_8655 = _T_8603[51]; // @[Bitwise.scala 50:65:@6617.4]
  assign _T_8656 = _T_8603[52]; // @[Bitwise.scala 50:65:@6618.4]
  assign _T_8657 = _T_8603[53]; // @[Bitwise.scala 50:65:@6619.4]
  assign _T_8658 = _T_8603[54]; // @[Bitwise.scala 50:65:@6620.4]
  assign _T_8659 = _T_8605 + _T_8606; // @[Bitwise.scala 48:55:@6621.4]
  assign _GEN_952 = {{1'd0}, _T_8604}; // @[Bitwise.scala 48:55:@6622.4]
  assign _T_8660 = _GEN_952 + _T_8659; // @[Bitwise.scala 48:55:@6622.4]
  assign _T_8661 = _T_8608 + _T_8609; // @[Bitwise.scala 48:55:@6623.4]
  assign _GEN_953 = {{1'd0}, _T_8607}; // @[Bitwise.scala 48:55:@6624.4]
  assign _T_8662 = _GEN_953 + _T_8661; // @[Bitwise.scala 48:55:@6624.4]
  assign _T_8663 = _T_8660 + _T_8662; // @[Bitwise.scala 48:55:@6625.4]
  assign _T_8664 = _T_8611 + _T_8612; // @[Bitwise.scala 48:55:@6626.4]
  assign _GEN_954 = {{1'd0}, _T_8610}; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_8665 = _GEN_954 + _T_8664; // @[Bitwise.scala 48:55:@6627.4]
  assign _T_8666 = _T_8613 + _T_8614; // @[Bitwise.scala 48:55:@6628.4]
  assign _T_8667 = _T_8615 + _T_8616; // @[Bitwise.scala 48:55:@6629.4]
  assign _T_8668 = _T_8666 + _T_8667; // @[Bitwise.scala 48:55:@6630.4]
  assign _T_8669 = _T_8665 + _T_8668; // @[Bitwise.scala 48:55:@6631.4]
  assign _T_8670 = _T_8663 + _T_8669; // @[Bitwise.scala 48:55:@6632.4]
  assign _T_8671 = _T_8618 + _T_8619; // @[Bitwise.scala 48:55:@6633.4]
  assign _GEN_955 = {{1'd0}, _T_8617}; // @[Bitwise.scala 48:55:@6634.4]
  assign _T_8672 = _GEN_955 + _T_8671; // @[Bitwise.scala 48:55:@6634.4]
  assign _T_8673 = _T_8620 + _T_8621; // @[Bitwise.scala 48:55:@6635.4]
  assign _T_8674 = _T_8622 + _T_8623; // @[Bitwise.scala 48:55:@6636.4]
  assign _T_8675 = _T_8673 + _T_8674; // @[Bitwise.scala 48:55:@6637.4]
  assign _T_8676 = _T_8672 + _T_8675; // @[Bitwise.scala 48:55:@6638.4]
  assign _T_8677 = _T_8625 + _T_8626; // @[Bitwise.scala 48:55:@6639.4]
  assign _GEN_956 = {{1'd0}, _T_8624}; // @[Bitwise.scala 48:55:@6640.4]
  assign _T_8678 = _GEN_956 + _T_8677; // @[Bitwise.scala 48:55:@6640.4]
  assign _T_8679 = _T_8627 + _T_8628; // @[Bitwise.scala 48:55:@6641.4]
  assign _T_8680 = _T_8629 + _T_8630; // @[Bitwise.scala 48:55:@6642.4]
  assign _T_8681 = _T_8679 + _T_8680; // @[Bitwise.scala 48:55:@6643.4]
  assign _T_8682 = _T_8678 + _T_8681; // @[Bitwise.scala 48:55:@6644.4]
  assign _T_8683 = _T_8676 + _T_8682; // @[Bitwise.scala 48:55:@6645.4]
  assign _T_8684 = _T_8670 + _T_8683; // @[Bitwise.scala 48:55:@6646.4]
  assign _T_8685 = _T_8632 + _T_8633; // @[Bitwise.scala 48:55:@6647.4]
  assign _GEN_957 = {{1'd0}, _T_8631}; // @[Bitwise.scala 48:55:@6648.4]
  assign _T_8686 = _GEN_957 + _T_8685; // @[Bitwise.scala 48:55:@6648.4]
  assign _T_8687 = _T_8634 + _T_8635; // @[Bitwise.scala 48:55:@6649.4]
  assign _T_8688 = _T_8636 + _T_8637; // @[Bitwise.scala 48:55:@6650.4]
  assign _T_8689 = _T_8687 + _T_8688; // @[Bitwise.scala 48:55:@6651.4]
  assign _T_8690 = _T_8686 + _T_8689; // @[Bitwise.scala 48:55:@6652.4]
  assign _T_8691 = _T_8639 + _T_8640; // @[Bitwise.scala 48:55:@6653.4]
  assign _GEN_958 = {{1'd0}, _T_8638}; // @[Bitwise.scala 48:55:@6654.4]
  assign _T_8692 = _GEN_958 + _T_8691; // @[Bitwise.scala 48:55:@6654.4]
  assign _T_8693 = _T_8641 + _T_8642; // @[Bitwise.scala 48:55:@6655.4]
  assign _T_8694 = _T_8643 + _T_8644; // @[Bitwise.scala 48:55:@6656.4]
  assign _T_8695 = _T_8693 + _T_8694; // @[Bitwise.scala 48:55:@6657.4]
  assign _T_8696 = _T_8692 + _T_8695; // @[Bitwise.scala 48:55:@6658.4]
  assign _T_8697 = _T_8690 + _T_8696; // @[Bitwise.scala 48:55:@6659.4]
  assign _T_8698 = _T_8646 + _T_8647; // @[Bitwise.scala 48:55:@6660.4]
  assign _GEN_959 = {{1'd0}, _T_8645}; // @[Bitwise.scala 48:55:@6661.4]
  assign _T_8699 = _GEN_959 + _T_8698; // @[Bitwise.scala 48:55:@6661.4]
  assign _T_8700 = _T_8648 + _T_8649; // @[Bitwise.scala 48:55:@6662.4]
  assign _T_8701 = _T_8650 + _T_8651; // @[Bitwise.scala 48:55:@6663.4]
  assign _T_8702 = _T_8700 + _T_8701; // @[Bitwise.scala 48:55:@6664.4]
  assign _T_8703 = _T_8699 + _T_8702; // @[Bitwise.scala 48:55:@6665.4]
  assign _T_8704 = _T_8653 + _T_8654; // @[Bitwise.scala 48:55:@6666.4]
  assign _GEN_960 = {{1'd0}, _T_8652}; // @[Bitwise.scala 48:55:@6667.4]
  assign _T_8705 = _GEN_960 + _T_8704; // @[Bitwise.scala 48:55:@6667.4]
  assign _T_8706 = _T_8655 + _T_8656; // @[Bitwise.scala 48:55:@6668.4]
  assign _T_8707 = _T_8657 + _T_8658; // @[Bitwise.scala 48:55:@6669.4]
  assign _T_8708 = _T_8706 + _T_8707; // @[Bitwise.scala 48:55:@6670.4]
  assign _T_8709 = _T_8705 + _T_8708; // @[Bitwise.scala 48:55:@6671.4]
  assign _T_8710 = _T_8703 + _T_8709; // @[Bitwise.scala 48:55:@6672.4]
  assign _T_8711 = _T_8697 + _T_8710; // @[Bitwise.scala 48:55:@6673.4]
  assign _T_8712 = _T_8684 + _T_8711; // @[Bitwise.scala 48:55:@6674.4]
  assign _T_8776 = _T_2230[55:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6739.4]
  assign _T_8777 = _T_8776[0]; // @[Bitwise.scala 50:65:@6740.4]
  assign _T_8778 = _T_8776[1]; // @[Bitwise.scala 50:65:@6741.4]
  assign _T_8779 = _T_8776[2]; // @[Bitwise.scala 50:65:@6742.4]
  assign _T_8780 = _T_8776[3]; // @[Bitwise.scala 50:65:@6743.4]
  assign _T_8781 = _T_8776[4]; // @[Bitwise.scala 50:65:@6744.4]
  assign _T_8782 = _T_8776[5]; // @[Bitwise.scala 50:65:@6745.4]
  assign _T_8783 = _T_8776[6]; // @[Bitwise.scala 50:65:@6746.4]
  assign _T_8784 = _T_8776[7]; // @[Bitwise.scala 50:65:@6747.4]
  assign _T_8785 = _T_8776[8]; // @[Bitwise.scala 50:65:@6748.4]
  assign _T_8786 = _T_8776[9]; // @[Bitwise.scala 50:65:@6749.4]
  assign _T_8787 = _T_8776[10]; // @[Bitwise.scala 50:65:@6750.4]
  assign _T_8788 = _T_8776[11]; // @[Bitwise.scala 50:65:@6751.4]
  assign _T_8789 = _T_8776[12]; // @[Bitwise.scala 50:65:@6752.4]
  assign _T_8790 = _T_8776[13]; // @[Bitwise.scala 50:65:@6753.4]
  assign _T_8791 = _T_8776[14]; // @[Bitwise.scala 50:65:@6754.4]
  assign _T_8792 = _T_8776[15]; // @[Bitwise.scala 50:65:@6755.4]
  assign _T_8793 = _T_8776[16]; // @[Bitwise.scala 50:65:@6756.4]
  assign _T_8794 = _T_8776[17]; // @[Bitwise.scala 50:65:@6757.4]
  assign _T_8795 = _T_8776[18]; // @[Bitwise.scala 50:65:@6758.4]
  assign _T_8796 = _T_8776[19]; // @[Bitwise.scala 50:65:@6759.4]
  assign _T_8797 = _T_8776[20]; // @[Bitwise.scala 50:65:@6760.4]
  assign _T_8798 = _T_8776[21]; // @[Bitwise.scala 50:65:@6761.4]
  assign _T_8799 = _T_8776[22]; // @[Bitwise.scala 50:65:@6762.4]
  assign _T_8800 = _T_8776[23]; // @[Bitwise.scala 50:65:@6763.4]
  assign _T_8801 = _T_8776[24]; // @[Bitwise.scala 50:65:@6764.4]
  assign _T_8802 = _T_8776[25]; // @[Bitwise.scala 50:65:@6765.4]
  assign _T_8803 = _T_8776[26]; // @[Bitwise.scala 50:65:@6766.4]
  assign _T_8804 = _T_8776[27]; // @[Bitwise.scala 50:65:@6767.4]
  assign _T_8805 = _T_8776[28]; // @[Bitwise.scala 50:65:@6768.4]
  assign _T_8806 = _T_8776[29]; // @[Bitwise.scala 50:65:@6769.4]
  assign _T_8807 = _T_8776[30]; // @[Bitwise.scala 50:65:@6770.4]
  assign _T_8808 = _T_8776[31]; // @[Bitwise.scala 50:65:@6771.4]
  assign _T_8809 = _T_8776[32]; // @[Bitwise.scala 50:65:@6772.4]
  assign _T_8810 = _T_8776[33]; // @[Bitwise.scala 50:65:@6773.4]
  assign _T_8811 = _T_8776[34]; // @[Bitwise.scala 50:65:@6774.4]
  assign _T_8812 = _T_8776[35]; // @[Bitwise.scala 50:65:@6775.4]
  assign _T_8813 = _T_8776[36]; // @[Bitwise.scala 50:65:@6776.4]
  assign _T_8814 = _T_8776[37]; // @[Bitwise.scala 50:65:@6777.4]
  assign _T_8815 = _T_8776[38]; // @[Bitwise.scala 50:65:@6778.4]
  assign _T_8816 = _T_8776[39]; // @[Bitwise.scala 50:65:@6779.4]
  assign _T_8817 = _T_8776[40]; // @[Bitwise.scala 50:65:@6780.4]
  assign _T_8818 = _T_8776[41]; // @[Bitwise.scala 50:65:@6781.4]
  assign _T_8819 = _T_8776[42]; // @[Bitwise.scala 50:65:@6782.4]
  assign _T_8820 = _T_8776[43]; // @[Bitwise.scala 50:65:@6783.4]
  assign _T_8821 = _T_8776[44]; // @[Bitwise.scala 50:65:@6784.4]
  assign _T_8822 = _T_8776[45]; // @[Bitwise.scala 50:65:@6785.4]
  assign _T_8823 = _T_8776[46]; // @[Bitwise.scala 50:65:@6786.4]
  assign _T_8824 = _T_8776[47]; // @[Bitwise.scala 50:65:@6787.4]
  assign _T_8825 = _T_8776[48]; // @[Bitwise.scala 50:65:@6788.4]
  assign _T_8826 = _T_8776[49]; // @[Bitwise.scala 50:65:@6789.4]
  assign _T_8827 = _T_8776[50]; // @[Bitwise.scala 50:65:@6790.4]
  assign _T_8828 = _T_8776[51]; // @[Bitwise.scala 50:65:@6791.4]
  assign _T_8829 = _T_8776[52]; // @[Bitwise.scala 50:65:@6792.4]
  assign _T_8830 = _T_8776[53]; // @[Bitwise.scala 50:65:@6793.4]
  assign _T_8831 = _T_8776[54]; // @[Bitwise.scala 50:65:@6794.4]
  assign _T_8832 = _T_8776[55]; // @[Bitwise.scala 50:65:@6795.4]
  assign _T_8833 = _T_8778 + _T_8779; // @[Bitwise.scala 48:55:@6796.4]
  assign _GEN_961 = {{1'd0}, _T_8777}; // @[Bitwise.scala 48:55:@6797.4]
  assign _T_8834 = _GEN_961 + _T_8833; // @[Bitwise.scala 48:55:@6797.4]
  assign _T_8835 = _T_8780 + _T_8781; // @[Bitwise.scala 48:55:@6798.4]
  assign _T_8836 = _T_8782 + _T_8783; // @[Bitwise.scala 48:55:@6799.4]
  assign _T_8837 = _T_8835 + _T_8836; // @[Bitwise.scala 48:55:@6800.4]
  assign _T_8838 = _T_8834 + _T_8837; // @[Bitwise.scala 48:55:@6801.4]
  assign _T_8839 = _T_8785 + _T_8786; // @[Bitwise.scala 48:55:@6802.4]
  assign _GEN_962 = {{1'd0}, _T_8784}; // @[Bitwise.scala 48:55:@6803.4]
  assign _T_8840 = _GEN_962 + _T_8839; // @[Bitwise.scala 48:55:@6803.4]
  assign _T_8841 = _T_8787 + _T_8788; // @[Bitwise.scala 48:55:@6804.4]
  assign _T_8842 = _T_8789 + _T_8790; // @[Bitwise.scala 48:55:@6805.4]
  assign _T_8843 = _T_8841 + _T_8842; // @[Bitwise.scala 48:55:@6806.4]
  assign _T_8844 = _T_8840 + _T_8843; // @[Bitwise.scala 48:55:@6807.4]
  assign _T_8845 = _T_8838 + _T_8844; // @[Bitwise.scala 48:55:@6808.4]
  assign _T_8846 = _T_8792 + _T_8793; // @[Bitwise.scala 48:55:@6809.4]
  assign _GEN_963 = {{1'd0}, _T_8791}; // @[Bitwise.scala 48:55:@6810.4]
  assign _T_8847 = _GEN_963 + _T_8846; // @[Bitwise.scala 48:55:@6810.4]
  assign _T_8848 = _T_8794 + _T_8795; // @[Bitwise.scala 48:55:@6811.4]
  assign _T_8849 = _T_8796 + _T_8797; // @[Bitwise.scala 48:55:@6812.4]
  assign _T_8850 = _T_8848 + _T_8849; // @[Bitwise.scala 48:55:@6813.4]
  assign _T_8851 = _T_8847 + _T_8850; // @[Bitwise.scala 48:55:@6814.4]
  assign _T_8852 = _T_8799 + _T_8800; // @[Bitwise.scala 48:55:@6815.4]
  assign _GEN_964 = {{1'd0}, _T_8798}; // @[Bitwise.scala 48:55:@6816.4]
  assign _T_8853 = _GEN_964 + _T_8852; // @[Bitwise.scala 48:55:@6816.4]
  assign _T_8854 = _T_8801 + _T_8802; // @[Bitwise.scala 48:55:@6817.4]
  assign _T_8855 = _T_8803 + _T_8804; // @[Bitwise.scala 48:55:@6818.4]
  assign _T_8856 = _T_8854 + _T_8855; // @[Bitwise.scala 48:55:@6819.4]
  assign _T_8857 = _T_8853 + _T_8856; // @[Bitwise.scala 48:55:@6820.4]
  assign _T_8858 = _T_8851 + _T_8857; // @[Bitwise.scala 48:55:@6821.4]
  assign _T_8859 = _T_8845 + _T_8858; // @[Bitwise.scala 48:55:@6822.4]
  assign _T_8860 = _T_8806 + _T_8807; // @[Bitwise.scala 48:55:@6823.4]
  assign _GEN_965 = {{1'd0}, _T_8805}; // @[Bitwise.scala 48:55:@6824.4]
  assign _T_8861 = _GEN_965 + _T_8860; // @[Bitwise.scala 48:55:@6824.4]
  assign _T_8862 = _T_8808 + _T_8809; // @[Bitwise.scala 48:55:@6825.4]
  assign _T_8863 = _T_8810 + _T_8811; // @[Bitwise.scala 48:55:@6826.4]
  assign _T_8864 = _T_8862 + _T_8863; // @[Bitwise.scala 48:55:@6827.4]
  assign _T_8865 = _T_8861 + _T_8864; // @[Bitwise.scala 48:55:@6828.4]
  assign _T_8866 = _T_8813 + _T_8814; // @[Bitwise.scala 48:55:@6829.4]
  assign _GEN_966 = {{1'd0}, _T_8812}; // @[Bitwise.scala 48:55:@6830.4]
  assign _T_8867 = _GEN_966 + _T_8866; // @[Bitwise.scala 48:55:@6830.4]
  assign _T_8868 = _T_8815 + _T_8816; // @[Bitwise.scala 48:55:@6831.4]
  assign _T_8869 = _T_8817 + _T_8818; // @[Bitwise.scala 48:55:@6832.4]
  assign _T_8870 = _T_8868 + _T_8869; // @[Bitwise.scala 48:55:@6833.4]
  assign _T_8871 = _T_8867 + _T_8870; // @[Bitwise.scala 48:55:@6834.4]
  assign _T_8872 = _T_8865 + _T_8871; // @[Bitwise.scala 48:55:@6835.4]
  assign _T_8873 = _T_8820 + _T_8821; // @[Bitwise.scala 48:55:@6836.4]
  assign _GEN_967 = {{1'd0}, _T_8819}; // @[Bitwise.scala 48:55:@6837.4]
  assign _T_8874 = _GEN_967 + _T_8873; // @[Bitwise.scala 48:55:@6837.4]
  assign _T_8875 = _T_8822 + _T_8823; // @[Bitwise.scala 48:55:@6838.4]
  assign _T_8876 = _T_8824 + _T_8825; // @[Bitwise.scala 48:55:@6839.4]
  assign _T_8877 = _T_8875 + _T_8876; // @[Bitwise.scala 48:55:@6840.4]
  assign _T_8878 = _T_8874 + _T_8877; // @[Bitwise.scala 48:55:@6841.4]
  assign _T_8879 = _T_8827 + _T_8828; // @[Bitwise.scala 48:55:@6842.4]
  assign _GEN_968 = {{1'd0}, _T_8826}; // @[Bitwise.scala 48:55:@6843.4]
  assign _T_8880 = _GEN_968 + _T_8879; // @[Bitwise.scala 48:55:@6843.4]
  assign _T_8881 = _T_8829 + _T_8830; // @[Bitwise.scala 48:55:@6844.4]
  assign _T_8882 = _T_8831 + _T_8832; // @[Bitwise.scala 48:55:@6845.4]
  assign _T_8883 = _T_8881 + _T_8882; // @[Bitwise.scala 48:55:@6846.4]
  assign _T_8884 = _T_8880 + _T_8883; // @[Bitwise.scala 48:55:@6847.4]
  assign _T_8885 = _T_8878 + _T_8884; // @[Bitwise.scala 48:55:@6848.4]
  assign _T_8886 = _T_8872 + _T_8885; // @[Bitwise.scala 48:55:@6849.4]
  assign _T_8887 = _T_8859 + _T_8886; // @[Bitwise.scala 48:55:@6850.4]
  assign _T_8951 = _T_2230[56:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@6915.4]
  assign _T_8952 = _T_8951[0]; // @[Bitwise.scala 50:65:@6916.4]
  assign _T_8953 = _T_8951[1]; // @[Bitwise.scala 50:65:@6917.4]
  assign _T_8954 = _T_8951[2]; // @[Bitwise.scala 50:65:@6918.4]
  assign _T_8955 = _T_8951[3]; // @[Bitwise.scala 50:65:@6919.4]
  assign _T_8956 = _T_8951[4]; // @[Bitwise.scala 50:65:@6920.4]
  assign _T_8957 = _T_8951[5]; // @[Bitwise.scala 50:65:@6921.4]
  assign _T_8958 = _T_8951[6]; // @[Bitwise.scala 50:65:@6922.4]
  assign _T_8959 = _T_8951[7]; // @[Bitwise.scala 50:65:@6923.4]
  assign _T_8960 = _T_8951[8]; // @[Bitwise.scala 50:65:@6924.4]
  assign _T_8961 = _T_8951[9]; // @[Bitwise.scala 50:65:@6925.4]
  assign _T_8962 = _T_8951[10]; // @[Bitwise.scala 50:65:@6926.4]
  assign _T_8963 = _T_8951[11]; // @[Bitwise.scala 50:65:@6927.4]
  assign _T_8964 = _T_8951[12]; // @[Bitwise.scala 50:65:@6928.4]
  assign _T_8965 = _T_8951[13]; // @[Bitwise.scala 50:65:@6929.4]
  assign _T_8966 = _T_8951[14]; // @[Bitwise.scala 50:65:@6930.4]
  assign _T_8967 = _T_8951[15]; // @[Bitwise.scala 50:65:@6931.4]
  assign _T_8968 = _T_8951[16]; // @[Bitwise.scala 50:65:@6932.4]
  assign _T_8969 = _T_8951[17]; // @[Bitwise.scala 50:65:@6933.4]
  assign _T_8970 = _T_8951[18]; // @[Bitwise.scala 50:65:@6934.4]
  assign _T_8971 = _T_8951[19]; // @[Bitwise.scala 50:65:@6935.4]
  assign _T_8972 = _T_8951[20]; // @[Bitwise.scala 50:65:@6936.4]
  assign _T_8973 = _T_8951[21]; // @[Bitwise.scala 50:65:@6937.4]
  assign _T_8974 = _T_8951[22]; // @[Bitwise.scala 50:65:@6938.4]
  assign _T_8975 = _T_8951[23]; // @[Bitwise.scala 50:65:@6939.4]
  assign _T_8976 = _T_8951[24]; // @[Bitwise.scala 50:65:@6940.4]
  assign _T_8977 = _T_8951[25]; // @[Bitwise.scala 50:65:@6941.4]
  assign _T_8978 = _T_8951[26]; // @[Bitwise.scala 50:65:@6942.4]
  assign _T_8979 = _T_8951[27]; // @[Bitwise.scala 50:65:@6943.4]
  assign _T_8980 = _T_8951[28]; // @[Bitwise.scala 50:65:@6944.4]
  assign _T_8981 = _T_8951[29]; // @[Bitwise.scala 50:65:@6945.4]
  assign _T_8982 = _T_8951[30]; // @[Bitwise.scala 50:65:@6946.4]
  assign _T_8983 = _T_8951[31]; // @[Bitwise.scala 50:65:@6947.4]
  assign _T_8984 = _T_8951[32]; // @[Bitwise.scala 50:65:@6948.4]
  assign _T_8985 = _T_8951[33]; // @[Bitwise.scala 50:65:@6949.4]
  assign _T_8986 = _T_8951[34]; // @[Bitwise.scala 50:65:@6950.4]
  assign _T_8987 = _T_8951[35]; // @[Bitwise.scala 50:65:@6951.4]
  assign _T_8988 = _T_8951[36]; // @[Bitwise.scala 50:65:@6952.4]
  assign _T_8989 = _T_8951[37]; // @[Bitwise.scala 50:65:@6953.4]
  assign _T_8990 = _T_8951[38]; // @[Bitwise.scala 50:65:@6954.4]
  assign _T_8991 = _T_8951[39]; // @[Bitwise.scala 50:65:@6955.4]
  assign _T_8992 = _T_8951[40]; // @[Bitwise.scala 50:65:@6956.4]
  assign _T_8993 = _T_8951[41]; // @[Bitwise.scala 50:65:@6957.4]
  assign _T_8994 = _T_8951[42]; // @[Bitwise.scala 50:65:@6958.4]
  assign _T_8995 = _T_8951[43]; // @[Bitwise.scala 50:65:@6959.4]
  assign _T_8996 = _T_8951[44]; // @[Bitwise.scala 50:65:@6960.4]
  assign _T_8997 = _T_8951[45]; // @[Bitwise.scala 50:65:@6961.4]
  assign _T_8998 = _T_8951[46]; // @[Bitwise.scala 50:65:@6962.4]
  assign _T_8999 = _T_8951[47]; // @[Bitwise.scala 50:65:@6963.4]
  assign _T_9000 = _T_8951[48]; // @[Bitwise.scala 50:65:@6964.4]
  assign _T_9001 = _T_8951[49]; // @[Bitwise.scala 50:65:@6965.4]
  assign _T_9002 = _T_8951[50]; // @[Bitwise.scala 50:65:@6966.4]
  assign _T_9003 = _T_8951[51]; // @[Bitwise.scala 50:65:@6967.4]
  assign _T_9004 = _T_8951[52]; // @[Bitwise.scala 50:65:@6968.4]
  assign _T_9005 = _T_8951[53]; // @[Bitwise.scala 50:65:@6969.4]
  assign _T_9006 = _T_8951[54]; // @[Bitwise.scala 50:65:@6970.4]
  assign _T_9007 = _T_8951[55]; // @[Bitwise.scala 50:65:@6971.4]
  assign _T_9008 = _T_8951[56]; // @[Bitwise.scala 50:65:@6972.4]
  assign _T_9009 = _T_8953 + _T_8954; // @[Bitwise.scala 48:55:@6973.4]
  assign _GEN_969 = {{1'd0}, _T_8952}; // @[Bitwise.scala 48:55:@6974.4]
  assign _T_9010 = _GEN_969 + _T_9009; // @[Bitwise.scala 48:55:@6974.4]
  assign _T_9011 = _T_8955 + _T_8956; // @[Bitwise.scala 48:55:@6975.4]
  assign _T_9012 = _T_8957 + _T_8958; // @[Bitwise.scala 48:55:@6976.4]
  assign _T_9013 = _T_9011 + _T_9012; // @[Bitwise.scala 48:55:@6977.4]
  assign _T_9014 = _T_9010 + _T_9013; // @[Bitwise.scala 48:55:@6978.4]
  assign _T_9015 = _T_8960 + _T_8961; // @[Bitwise.scala 48:55:@6979.4]
  assign _GEN_970 = {{1'd0}, _T_8959}; // @[Bitwise.scala 48:55:@6980.4]
  assign _T_9016 = _GEN_970 + _T_9015; // @[Bitwise.scala 48:55:@6980.4]
  assign _T_9017 = _T_8962 + _T_8963; // @[Bitwise.scala 48:55:@6981.4]
  assign _T_9018 = _T_8964 + _T_8965; // @[Bitwise.scala 48:55:@6982.4]
  assign _T_9019 = _T_9017 + _T_9018; // @[Bitwise.scala 48:55:@6983.4]
  assign _T_9020 = _T_9016 + _T_9019; // @[Bitwise.scala 48:55:@6984.4]
  assign _T_9021 = _T_9014 + _T_9020; // @[Bitwise.scala 48:55:@6985.4]
  assign _T_9022 = _T_8967 + _T_8968; // @[Bitwise.scala 48:55:@6986.4]
  assign _GEN_971 = {{1'd0}, _T_8966}; // @[Bitwise.scala 48:55:@6987.4]
  assign _T_9023 = _GEN_971 + _T_9022; // @[Bitwise.scala 48:55:@6987.4]
  assign _T_9024 = _T_8969 + _T_8970; // @[Bitwise.scala 48:55:@6988.4]
  assign _T_9025 = _T_8971 + _T_8972; // @[Bitwise.scala 48:55:@6989.4]
  assign _T_9026 = _T_9024 + _T_9025; // @[Bitwise.scala 48:55:@6990.4]
  assign _T_9027 = _T_9023 + _T_9026; // @[Bitwise.scala 48:55:@6991.4]
  assign _T_9028 = _T_8974 + _T_8975; // @[Bitwise.scala 48:55:@6992.4]
  assign _GEN_972 = {{1'd0}, _T_8973}; // @[Bitwise.scala 48:55:@6993.4]
  assign _T_9029 = _GEN_972 + _T_9028; // @[Bitwise.scala 48:55:@6993.4]
  assign _T_9030 = _T_8976 + _T_8977; // @[Bitwise.scala 48:55:@6994.4]
  assign _T_9031 = _T_8978 + _T_8979; // @[Bitwise.scala 48:55:@6995.4]
  assign _T_9032 = _T_9030 + _T_9031; // @[Bitwise.scala 48:55:@6996.4]
  assign _T_9033 = _T_9029 + _T_9032; // @[Bitwise.scala 48:55:@6997.4]
  assign _T_9034 = _T_9027 + _T_9033; // @[Bitwise.scala 48:55:@6998.4]
  assign _T_9035 = _T_9021 + _T_9034; // @[Bitwise.scala 48:55:@6999.4]
  assign _T_9036 = _T_8981 + _T_8982; // @[Bitwise.scala 48:55:@7000.4]
  assign _GEN_973 = {{1'd0}, _T_8980}; // @[Bitwise.scala 48:55:@7001.4]
  assign _T_9037 = _GEN_973 + _T_9036; // @[Bitwise.scala 48:55:@7001.4]
  assign _T_9038 = _T_8983 + _T_8984; // @[Bitwise.scala 48:55:@7002.4]
  assign _T_9039 = _T_8985 + _T_8986; // @[Bitwise.scala 48:55:@7003.4]
  assign _T_9040 = _T_9038 + _T_9039; // @[Bitwise.scala 48:55:@7004.4]
  assign _T_9041 = _T_9037 + _T_9040; // @[Bitwise.scala 48:55:@7005.4]
  assign _T_9042 = _T_8988 + _T_8989; // @[Bitwise.scala 48:55:@7006.4]
  assign _GEN_974 = {{1'd0}, _T_8987}; // @[Bitwise.scala 48:55:@7007.4]
  assign _T_9043 = _GEN_974 + _T_9042; // @[Bitwise.scala 48:55:@7007.4]
  assign _T_9044 = _T_8990 + _T_8991; // @[Bitwise.scala 48:55:@7008.4]
  assign _T_9045 = _T_8992 + _T_8993; // @[Bitwise.scala 48:55:@7009.4]
  assign _T_9046 = _T_9044 + _T_9045; // @[Bitwise.scala 48:55:@7010.4]
  assign _T_9047 = _T_9043 + _T_9046; // @[Bitwise.scala 48:55:@7011.4]
  assign _T_9048 = _T_9041 + _T_9047; // @[Bitwise.scala 48:55:@7012.4]
  assign _T_9049 = _T_8995 + _T_8996; // @[Bitwise.scala 48:55:@7013.4]
  assign _GEN_975 = {{1'd0}, _T_8994}; // @[Bitwise.scala 48:55:@7014.4]
  assign _T_9050 = _GEN_975 + _T_9049; // @[Bitwise.scala 48:55:@7014.4]
  assign _T_9051 = _T_8997 + _T_8998; // @[Bitwise.scala 48:55:@7015.4]
  assign _T_9052 = _T_8999 + _T_9000; // @[Bitwise.scala 48:55:@7016.4]
  assign _T_9053 = _T_9051 + _T_9052; // @[Bitwise.scala 48:55:@7017.4]
  assign _T_9054 = _T_9050 + _T_9053; // @[Bitwise.scala 48:55:@7018.4]
  assign _T_9055 = _T_9001 + _T_9002; // @[Bitwise.scala 48:55:@7019.4]
  assign _T_9056 = _T_9003 + _T_9004; // @[Bitwise.scala 48:55:@7020.4]
  assign _T_9057 = _T_9055 + _T_9056; // @[Bitwise.scala 48:55:@7021.4]
  assign _T_9058 = _T_9005 + _T_9006; // @[Bitwise.scala 48:55:@7022.4]
  assign _T_9059 = _T_9007 + _T_9008; // @[Bitwise.scala 48:55:@7023.4]
  assign _T_9060 = _T_9058 + _T_9059; // @[Bitwise.scala 48:55:@7024.4]
  assign _T_9061 = _T_9057 + _T_9060; // @[Bitwise.scala 48:55:@7025.4]
  assign _T_9062 = _T_9054 + _T_9061; // @[Bitwise.scala 48:55:@7026.4]
  assign _T_9063 = _T_9048 + _T_9062; // @[Bitwise.scala 48:55:@7027.4]
  assign _T_9064 = _T_9035 + _T_9063; // @[Bitwise.scala 48:55:@7028.4]
  assign _T_9128 = _T_2230[57:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7093.4]
  assign _T_9129 = _T_9128[0]; // @[Bitwise.scala 50:65:@7094.4]
  assign _T_9130 = _T_9128[1]; // @[Bitwise.scala 50:65:@7095.4]
  assign _T_9131 = _T_9128[2]; // @[Bitwise.scala 50:65:@7096.4]
  assign _T_9132 = _T_9128[3]; // @[Bitwise.scala 50:65:@7097.4]
  assign _T_9133 = _T_9128[4]; // @[Bitwise.scala 50:65:@7098.4]
  assign _T_9134 = _T_9128[5]; // @[Bitwise.scala 50:65:@7099.4]
  assign _T_9135 = _T_9128[6]; // @[Bitwise.scala 50:65:@7100.4]
  assign _T_9136 = _T_9128[7]; // @[Bitwise.scala 50:65:@7101.4]
  assign _T_9137 = _T_9128[8]; // @[Bitwise.scala 50:65:@7102.4]
  assign _T_9138 = _T_9128[9]; // @[Bitwise.scala 50:65:@7103.4]
  assign _T_9139 = _T_9128[10]; // @[Bitwise.scala 50:65:@7104.4]
  assign _T_9140 = _T_9128[11]; // @[Bitwise.scala 50:65:@7105.4]
  assign _T_9141 = _T_9128[12]; // @[Bitwise.scala 50:65:@7106.4]
  assign _T_9142 = _T_9128[13]; // @[Bitwise.scala 50:65:@7107.4]
  assign _T_9143 = _T_9128[14]; // @[Bitwise.scala 50:65:@7108.4]
  assign _T_9144 = _T_9128[15]; // @[Bitwise.scala 50:65:@7109.4]
  assign _T_9145 = _T_9128[16]; // @[Bitwise.scala 50:65:@7110.4]
  assign _T_9146 = _T_9128[17]; // @[Bitwise.scala 50:65:@7111.4]
  assign _T_9147 = _T_9128[18]; // @[Bitwise.scala 50:65:@7112.4]
  assign _T_9148 = _T_9128[19]; // @[Bitwise.scala 50:65:@7113.4]
  assign _T_9149 = _T_9128[20]; // @[Bitwise.scala 50:65:@7114.4]
  assign _T_9150 = _T_9128[21]; // @[Bitwise.scala 50:65:@7115.4]
  assign _T_9151 = _T_9128[22]; // @[Bitwise.scala 50:65:@7116.4]
  assign _T_9152 = _T_9128[23]; // @[Bitwise.scala 50:65:@7117.4]
  assign _T_9153 = _T_9128[24]; // @[Bitwise.scala 50:65:@7118.4]
  assign _T_9154 = _T_9128[25]; // @[Bitwise.scala 50:65:@7119.4]
  assign _T_9155 = _T_9128[26]; // @[Bitwise.scala 50:65:@7120.4]
  assign _T_9156 = _T_9128[27]; // @[Bitwise.scala 50:65:@7121.4]
  assign _T_9157 = _T_9128[28]; // @[Bitwise.scala 50:65:@7122.4]
  assign _T_9158 = _T_9128[29]; // @[Bitwise.scala 50:65:@7123.4]
  assign _T_9159 = _T_9128[30]; // @[Bitwise.scala 50:65:@7124.4]
  assign _T_9160 = _T_9128[31]; // @[Bitwise.scala 50:65:@7125.4]
  assign _T_9161 = _T_9128[32]; // @[Bitwise.scala 50:65:@7126.4]
  assign _T_9162 = _T_9128[33]; // @[Bitwise.scala 50:65:@7127.4]
  assign _T_9163 = _T_9128[34]; // @[Bitwise.scala 50:65:@7128.4]
  assign _T_9164 = _T_9128[35]; // @[Bitwise.scala 50:65:@7129.4]
  assign _T_9165 = _T_9128[36]; // @[Bitwise.scala 50:65:@7130.4]
  assign _T_9166 = _T_9128[37]; // @[Bitwise.scala 50:65:@7131.4]
  assign _T_9167 = _T_9128[38]; // @[Bitwise.scala 50:65:@7132.4]
  assign _T_9168 = _T_9128[39]; // @[Bitwise.scala 50:65:@7133.4]
  assign _T_9169 = _T_9128[40]; // @[Bitwise.scala 50:65:@7134.4]
  assign _T_9170 = _T_9128[41]; // @[Bitwise.scala 50:65:@7135.4]
  assign _T_9171 = _T_9128[42]; // @[Bitwise.scala 50:65:@7136.4]
  assign _T_9172 = _T_9128[43]; // @[Bitwise.scala 50:65:@7137.4]
  assign _T_9173 = _T_9128[44]; // @[Bitwise.scala 50:65:@7138.4]
  assign _T_9174 = _T_9128[45]; // @[Bitwise.scala 50:65:@7139.4]
  assign _T_9175 = _T_9128[46]; // @[Bitwise.scala 50:65:@7140.4]
  assign _T_9176 = _T_9128[47]; // @[Bitwise.scala 50:65:@7141.4]
  assign _T_9177 = _T_9128[48]; // @[Bitwise.scala 50:65:@7142.4]
  assign _T_9178 = _T_9128[49]; // @[Bitwise.scala 50:65:@7143.4]
  assign _T_9179 = _T_9128[50]; // @[Bitwise.scala 50:65:@7144.4]
  assign _T_9180 = _T_9128[51]; // @[Bitwise.scala 50:65:@7145.4]
  assign _T_9181 = _T_9128[52]; // @[Bitwise.scala 50:65:@7146.4]
  assign _T_9182 = _T_9128[53]; // @[Bitwise.scala 50:65:@7147.4]
  assign _T_9183 = _T_9128[54]; // @[Bitwise.scala 50:65:@7148.4]
  assign _T_9184 = _T_9128[55]; // @[Bitwise.scala 50:65:@7149.4]
  assign _T_9185 = _T_9128[56]; // @[Bitwise.scala 50:65:@7150.4]
  assign _T_9186 = _T_9128[57]; // @[Bitwise.scala 50:65:@7151.4]
  assign _T_9187 = _T_9130 + _T_9131; // @[Bitwise.scala 48:55:@7152.4]
  assign _GEN_976 = {{1'd0}, _T_9129}; // @[Bitwise.scala 48:55:@7153.4]
  assign _T_9188 = _GEN_976 + _T_9187; // @[Bitwise.scala 48:55:@7153.4]
  assign _T_9189 = _T_9132 + _T_9133; // @[Bitwise.scala 48:55:@7154.4]
  assign _T_9190 = _T_9134 + _T_9135; // @[Bitwise.scala 48:55:@7155.4]
  assign _T_9191 = _T_9189 + _T_9190; // @[Bitwise.scala 48:55:@7156.4]
  assign _T_9192 = _T_9188 + _T_9191; // @[Bitwise.scala 48:55:@7157.4]
  assign _T_9193 = _T_9137 + _T_9138; // @[Bitwise.scala 48:55:@7158.4]
  assign _GEN_977 = {{1'd0}, _T_9136}; // @[Bitwise.scala 48:55:@7159.4]
  assign _T_9194 = _GEN_977 + _T_9193; // @[Bitwise.scala 48:55:@7159.4]
  assign _T_9195 = _T_9139 + _T_9140; // @[Bitwise.scala 48:55:@7160.4]
  assign _T_9196 = _T_9141 + _T_9142; // @[Bitwise.scala 48:55:@7161.4]
  assign _T_9197 = _T_9195 + _T_9196; // @[Bitwise.scala 48:55:@7162.4]
  assign _T_9198 = _T_9194 + _T_9197; // @[Bitwise.scala 48:55:@7163.4]
  assign _T_9199 = _T_9192 + _T_9198; // @[Bitwise.scala 48:55:@7164.4]
  assign _T_9200 = _T_9144 + _T_9145; // @[Bitwise.scala 48:55:@7165.4]
  assign _GEN_978 = {{1'd0}, _T_9143}; // @[Bitwise.scala 48:55:@7166.4]
  assign _T_9201 = _GEN_978 + _T_9200; // @[Bitwise.scala 48:55:@7166.4]
  assign _T_9202 = _T_9146 + _T_9147; // @[Bitwise.scala 48:55:@7167.4]
  assign _T_9203 = _T_9148 + _T_9149; // @[Bitwise.scala 48:55:@7168.4]
  assign _T_9204 = _T_9202 + _T_9203; // @[Bitwise.scala 48:55:@7169.4]
  assign _T_9205 = _T_9201 + _T_9204; // @[Bitwise.scala 48:55:@7170.4]
  assign _T_9206 = _T_9150 + _T_9151; // @[Bitwise.scala 48:55:@7171.4]
  assign _T_9207 = _T_9152 + _T_9153; // @[Bitwise.scala 48:55:@7172.4]
  assign _T_9208 = _T_9206 + _T_9207; // @[Bitwise.scala 48:55:@7173.4]
  assign _T_9209 = _T_9154 + _T_9155; // @[Bitwise.scala 48:55:@7174.4]
  assign _T_9210 = _T_9156 + _T_9157; // @[Bitwise.scala 48:55:@7175.4]
  assign _T_9211 = _T_9209 + _T_9210; // @[Bitwise.scala 48:55:@7176.4]
  assign _T_9212 = _T_9208 + _T_9211; // @[Bitwise.scala 48:55:@7177.4]
  assign _T_9213 = _T_9205 + _T_9212; // @[Bitwise.scala 48:55:@7178.4]
  assign _T_9214 = _T_9199 + _T_9213; // @[Bitwise.scala 48:55:@7179.4]
  assign _T_9215 = _T_9159 + _T_9160; // @[Bitwise.scala 48:55:@7180.4]
  assign _GEN_979 = {{1'd0}, _T_9158}; // @[Bitwise.scala 48:55:@7181.4]
  assign _T_9216 = _GEN_979 + _T_9215; // @[Bitwise.scala 48:55:@7181.4]
  assign _T_9217 = _T_9161 + _T_9162; // @[Bitwise.scala 48:55:@7182.4]
  assign _T_9218 = _T_9163 + _T_9164; // @[Bitwise.scala 48:55:@7183.4]
  assign _T_9219 = _T_9217 + _T_9218; // @[Bitwise.scala 48:55:@7184.4]
  assign _T_9220 = _T_9216 + _T_9219; // @[Bitwise.scala 48:55:@7185.4]
  assign _T_9221 = _T_9166 + _T_9167; // @[Bitwise.scala 48:55:@7186.4]
  assign _GEN_980 = {{1'd0}, _T_9165}; // @[Bitwise.scala 48:55:@7187.4]
  assign _T_9222 = _GEN_980 + _T_9221; // @[Bitwise.scala 48:55:@7187.4]
  assign _T_9223 = _T_9168 + _T_9169; // @[Bitwise.scala 48:55:@7188.4]
  assign _T_9224 = _T_9170 + _T_9171; // @[Bitwise.scala 48:55:@7189.4]
  assign _T_9225 = _T_9223 + _T_9224; // @[Bitwise.scala 48:55:@7190.4]
  assign _T_9226 = _T_9222 + _T_9225; // @[Bitwise.scala 48:55:@7191.4]
  assign _T_9227 = _T_9220 + _T_9226; // @[Bitwise.scala 48:55:@7192.4]
  assign _T_9228 = _T_9173 + _T_9174; // @[Bitwise.scala 48:55:@7193.4]
  assign _GEN_981 = {{1'd0}, _T_9172}; // @[Bitwise.scala 48:55:@7194.4]
  assign _T_9229 = _GEN_981 + _T_9228; // @[Bitwise.scala 48:55:@7194.4]
  assign _T_9230 = _T_9175 + _T_9176; // @[Bitwise.scala 48:55:@7195.4]
  assign _T_9231 = _T_9177 + _T_9178; // @[Bitwise.scala 48:55:@7196.4]
  assign _T_9232 = _T_9230 + _T_9231; // @[Bitwise.scala 48:55:@7197.4]
  assign _T_9233 = _T_9229 + _T_9232; // @[Bitwise.scala 48:55:@7198.4]
  assign _T_9234 = _T_9179 + _T_9180; // @[Bitwise.scala 48:55:@7199.4]
  assign _T_9235 = _T_9181 + _T_9182; // @[Bitwise.scala 48:55:@7200.4]
  assign _T_9236 = _T_9234 + _T_9235; // @[Bitwise.scala 48:55:@7201.4]
  assign _T_9237 = _T_9183 + _T_9184; // @[Bitwise.scala 48:55:@7202.4]
  assign _T_9238 = _T_9185 + _T_9186; // @[Bitwise.scala 48:55:@7203.4]
  assign _T_9239 = _T_9237 + _T_9238; // @[Bitwise.scala 48:55:@7204.4]
  assign _T_9240 = _T_9236 + _T_9239; // @[Bitwise.scala 48:55:@7205.4]
  assign _T_9241 = _T_9233 + _T_9240; // @[Bitwise.scala 48:55:@7206.4]
  assign _T_9242 = _T_9227 + _T_9241; // @[Bitwise.scala 48:55:@7207.4]
  assign _T_9243 = _T_9214 + _T_9242; // @[Bitwise.scala 48:55:@7208.4]
  assign _T_9307 = _T_2230[58:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7273.4]
  assign _T_9308 = _T_9307[0]; // @[Bitwise.scala 50:65:@7274.4]
  assign _T_9309 = _T_9307[1]; // @[Bitwise.scala 50:65:@7275.4]
  assign _T_9310 = _T_9307[2]; // @[Bitwise.scala 50:65:@7276.4]
  assign _T_9311 = _T_9307[3]; // @[Bitwise.scala 50:65:@7277.4]
  assign _T_9312 = _T_9307[4]; // @[Bitwise.scala 50:65:@7278.4]
  assign _T_9313 = _T_9307[5]; // @[Bitwise.scala 50:65:@7279.4]
  assign _T_9314 = _T_9307[6]; // @[Bitwise.scala 50:65:@7280.4]
  assign _T_9315 = _T_9307[7]; // @[Bitwise.scala 50:65:@7281.4]
  assign _T_9316 = _T_9307[8]; // @[Bitwise.scala 50:65:@7282.4]
  assign _T_9317 = _T_9307[9]; // @[Bitwise.scala 50:65:@7283.4]
  assign _T_9318 = _T_9307[10]; // @[Bitwise.scala 50:65:@7284.4]
  assign _T_9319 = _T_9307[11]; // @[Bitwise.scala 50:65:@7285.4]
  assign _T_9320 = _T_9307[12]; // @[Bitwise.scala 50:65:@7286.4]
  assign _T_9321 = _T_9307[13]; // @[Bitwise.scala 50:65:@7287.4]
  assign _T_9322 = _T_9307[14]; // @[Bitwise.scala 50:65:@7288.4]
  assign _T_9323 = _T_9307[15]; // @[Bitwise.scala 50:65:@7289.4]
  assign _T_9324 = _T_9307[16]; // @[Bitwise.scala 50:65:@7290.4]
  assign _T_9325 = _T_9307[17]; // @[Bitwise.scala 50:65:@7291.4]
  assign _T_9326 = _T_9307[18]; // @[Bitwise.scala 50:65:@7292.4]
  assign _T_9327 = _T_9307[19]; // @[Bitwise.scala 50:65:@7293.4]
  assign _T_9328 = _T_9307[20]; // @[Bitwise.scala 50:65:@7294.4]
  assign _T_9329 = _T_9307[21]; // @[Bitwise.scala 50:65:@7295.4]
  assign _T_9330 = _T_9307[22]; // @[Bitwise.scala 50:65:@7296.4]
  assign _T_9331 = _T_9307[23]; // @[Bitwise.scala 50:65:@7297.4]
  assign _T_9332 = _T_9307[24]; // @[Bitwise.scala 50:65:@7298.4]
  assign _T_9333 = _T_9307[25]; // @[Bitwise.scala 50:65:@7299.4]
  assign _T_9334 = _T_9307[26]; // @[Bitwise.scala 50:65:@7300.4]
  assign _T_9335 = _T_9307[27]; // @[Bitwise.scala 50:65:@7301.4]
  assign _T_9336 = _T_9307[28]; // @[Bitwise.scala 50:65:@7302.4]
  assign _T_9337 = _T_9307[29]; // @[Bitwise.scala 50:65:@7303.4]
  assign _T_9338 = _T_9307[30]; // @[Bitwise.scala 50:65:@7304.4]
  assign _T_9339 = _T_9307[31]; // @[Bitwise.scala 50:65:@7305.4]
  assign _T_9340 = _T_9307[32]; // @[Bitwise.scala 50:65:@7306.4]
  assign _T_9341 = _T_9307[33]; // @[Bitwise.scala 50:65:@7307.4]
  assign _T_9342 = _T_9307[34]; // @[Bitwise.scala 50:65:@7308.4]
  assign _T_9343 = _T_9307[35]; // @[Bitwise.scala 50:65:@7309.4]
  assign _T_9344 = _T_9307[36]; // @[Bitwise.scala 50:65:@7310.4]
  assign _T_9345 = _T_9307[37]; // @[Bitwise.scala 50:65:@7311.4]
  assign _T_9346 = _T_9307[38]; // @[Bitwise.scala 50:65:@7312.4]
  assign _T_9347 = _T_9307[39]; // @[Bitwise.scala 50:65:@7313.4]
  assign _T_9348 = _T_9307[40]; // @[Bitwise.scala 50:65:@7314.4]
  assign _T_9349 = _T_9307[41]; // @[Bitwise.scala 50:65:@7315.4]
  assign _T_9350 = _T_9307[42]; // @[Bitwise.scala 50:65:@7316.4]
  assign _T_9351 = _T_9307[43]; // @[Bitwise.scala 50:65:@7317.4]
  assign _T_9352 = _T_9307[44]; // @[Bitwise.scala 50:65:@7318.4]
  assign _T_9353 = _T_9307[45]; // @[Bitwise.scala 50:65:@7319.4]
  assign _T_9354 = _T_9307[46]; // @[Bitwise.scala 50:65:@7320.4]
  assign _T_9355 = _T_9307[47]; // @[Bitwise.scala 50:65:@7321.4]
  assign _T_9356 = _T_9307[48]; // @[Bitwise.scala 50:65:@7322.4]
  assign _T_9357 = _T_9307[49]; // @[Bitwise.scala 50:65:@7323.4]
  assign _T_9358 = _T_9307[50]; // @[Bitwise.scala 50:65:@7324.4]
  assign _T_9359 = _T_9307[51]; // @[Bitwise.scala 50:65:@7325.4]
  assign _T_9360 = _T_9307[52]; // @[Bitwise.scala 50:65:@7326.4]
  assign _T_9361 = _T_9307[53]; // @[Bitwise.scala 50:65:@7327.4]
  assign _T_9362 = _T_9307[54]; // @[Bitwise.scala 50:65:@7328.4]
  assign _T_9363 = _T_9307[55]; // @[Bitwise.scala 50:65:@7329.4]
  assign _T_9364 = _T_9307[56]; // @[Bitwise.scala 50:65:@7330.4]
  assign _T_9365 = _T_9307[57]; // @[Bitwise.scala 50:65:@7331.4]
  assign _T_9366 = _T_9307[58]; // @[Bitwise.scala 50:65:@7332.4]
  assign _T_9367 = _T_9309 + _T_9310; // @[Bitwise.scala 48:55:@7333.4]
  assign _GEN_982 = {{1'd0}, _T_9308}; // @[Bitwise.scala 48:55:@7334.4]
  assign _T_9368 = _GEN_982 + _T_9367; // @[Bitwise.scala 48:55:@7334.4]
  assign _T_9369 = _T_9311 + _T_9312; // @[Bitwise.scala 48:55:@7335.4]
  assign _T_9370 = _T_9313 + _T_9314; // @[Bitwise.scala 48:55:@7336.4]
  assign _T_9371 = _T_9369 + _T_9370; // @[Bitwise.scala 48:55:@7337.4]
  assign _T_9372 = _T_9368 + _T_9371; // @[Bitwise.scala 48:55:@7338.4]
  assign _T_9373 = _T_9316 + _T_9317; // @[Bitwise.scala 48:55:@7339.4]
  assign _GEN_983 = {{1'd0}, _T_9315}; // @[Bitwise.scala 48:55:@7340.4]
  assign _T_9374 = _GEN_983 + _T_9373; // @[Bitwise.scala 48:55:@7340.4]
  assign _T_9375 = _T_9318 + _T_9319; // @[Bitwise.scala 48:55:@7341.4]
  assign _T_9376 = _T_9320 + _T_9321; // @[Bitwise.scala 48:55:@7342.4]
  assign _T_9377 = _T_9375 + _T_9376; // @[Bitwise.scala 48:55:@7343.4]
  assign _T_9378 = _T_9374 + _T_9377; // @[Bitwise.scala 48:55:@7344.4]
  assign _T_9379 = _T_9372 + _T_9378; // @[Bitwise.scala 48:55:@7345.4]
  assign _T_9380 = _T_9323 + _T_9324; // @[Bitwise.scala 48:55:@7346.4]
  assign _GEN_984 = {{1'd0}, _T_9322}; // @[Bitwise.scala 48:55:@7347.4]
  assign _T_9381 = _GEN_984 + _T_9380; // @[Bitwise.scala 48:55:@7347.4]
  assign _T_9382 = _T_9325 + _T_9326; // @[Bitwise.scala 48:55:@7348.4]
  assign _T_9383 = _T_9327 + _T_9328; // @[Bitwise.scala 48:55:@7349.4]
  assign _T_9384 = _T_9382 + _T_9383; // @[Bitwise.scala 48:55:@7350.4]
  assign _T_9385 = _T_9381 + _T_9384; // @[Bitwise.scala 48:55:@7351.4]
  assign _T_9386 = _T_9329 + _T_9330; // @[Bitwise.scala 48:55:@7352.4]
  assign _T_9387 = _T_9331 + _T_9332; // @[Bitwise.scala 48:55:@7353.4]
  assign _T_9388 = _T_9386 + _T_9387; // @[Bitwise.scala 48:55:@7354.4]
  assign _T_9389 = _T_9333 + _T_9334; // @[Bitwise.scala 48:55:@7355.4]
  assign _T_9390 = _T_9335 + _T_9336; // @[Bitwise.scala 48:55:@7356.4]
  assign _T_9391 = _T_9389 + _T_9390; // @[Bitwise.scala 48:55:@7357.4]
  assign _T_9392 = _T_9388 + _T_9391; // @[Bitwise.scala 48:55:@7358.4]
  assign _T_9393 = _T_9385 + _T_9392; // @[Bitwise.scala 48:55:@7359.4]
  assign _T_9394 = _T_9379 + _T_9393; // @[Bitwise.scala 48:55:@7360.4]
  assign _T_9395 = _T_9338 + _T_9339; // @[Bitwise.scala 48:55:@7361.4]
  assign _GEN_985 = {{1'd0}, _T_9337}; // @[Bitwise.scala 48:55:@7362.4]
  assign _T_9396 = _GEN_985 + _T_9395; // @[Bitwise.scala 48:55:@7362.4]
  assign _T_9397 = _T_9340 + _T_9341; // @[Bitwise.scala 48:55:@7363.4]
  assign _T_9398 = _T_9342 + _T_9343; // @[Bitwise.scala 48:55:@7364.4]
  assign _T_9399 = _T_9397 + _T_9398; // @[Bitwise.scala 48:55:@7365.4]
  assign _T_9400 = _T_9396 + _T_9399; // @[Bitwise.scala 48:55:@7366.4]
  assign _T_9401 = _T_9344 + _T_9345; // @[Bitwise.scala 48:55:@7367.4]
  assign _T_9402 = _T_9346 + _T_9347; // @[Bitwise.scala 48:55:@7368.4]
  assign _T_9403 = _T_9401 + _T_9402; // @[Bitwise.scala 48:55:@7369.4]
  assign _T_9404 = _T_9348 + _T_9349; // @[Bitwise.scala 48:55:@7370.4]
  assign _T_9405 = _T_9350 + _T_9351; // @[Bitwise.scala 48:55:@7371.4]
  assign _T_9406 = _T_9404 + _T_9405; // @[Bitwise.scala 48:55:@7372.4]
  assign _T_9407 = _T_9403 + _T_9406; // @[Bitwise.scala 48:55:@7373.4]
  assign _T_9408 = _T_9400 + _T_9407; // @[Bitwise.scala 48:55:@7374.4]
  assign _T_9409 = _T_9353 + _T_9354; // @[Bitwise.scala 48:55:@7375.4]
  assign _GEN_986 = {{1'd0}, _T_9352}; // @[Bitwise.scala 48:55:@7376.4]
  assign _T_9410 = _GEN_986 + _T_9409; // @[Bitwise.scala 48:55:@7376.4]
  assign _T_9411 = _T_9355 + _T_9356; // @[Bitwise.scala 48:55:@7377.4]
  assign _T_9412 = _T_9357 + _T_9358; // @[Bitwise.scala 48:55:@7378.4]
  assign _T_9413 = _T_9411 + _T_9412; // @[Bitwise.scala 48:55:@7379.4]
  assign _T_9414 = _T_9410 + _T_9413; // @[Bitwise.scala 48:55:@7380.4]
  assign _T_9415 = _T_9359 + _T_9360; // @[Bitwise.scala 48:55:@7381.4]
  assign _T_9416 = _T_9361 + _T_9362; // @[Bitwise.scala 48:55:@7382.4]
  assign _T_9417 = _T_9415 + _T_9416; // @[Bitwise.scala 48:55:@7383.4]
  assign _T_9418 = _T_9363 + _T_9364; // @[Bitwise.scala 48:55:@7384.4]
  assign _T_9419 = _T_9365 + _T_9366; // @[Bitwise.scala 48:55:@7385.4]
  assign _T_9420 = _T_9418 + _T_9419; // @[Bitwise.scala 48:55:@7386.4]
  assign _T_9421 = _T_9417 + _T_9420; // @[Bitwise.scala 48:55:@7387.4]
  assign _T_9422 = _T_9414 + _T_9421; // @[Bitwise.scala 48:55:@7388.4]
  assign _T_9423 = _T_9408 + _T_9422; // @[Bitwise.scala 48:55:@7389.4]
  assign _T_9424 = _T_9394 + _T_9423; // @[Bitwise.scala 48:55:@7390.4]
  assign _T_9488 = _T_2230[59:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7455.4]
  assign _T_9489 = _T_9488[0]; // @[Bitwise.scala 50:65:@7456.4]
  assign _T_9490 = _T_9488[1]; // @[Bitwise.scala 50:65:@7457.4]
  assign _T_9491 = _T_9488[2]; // @[Bitwise.scala 50:65:@7458.4]
  assign _T_9492 = _T_9488[3]; // @[Bitwise.scala 50:65:@7459.4]
  assign _T_9493 = _T_9488[4]; // @[Bitwise.scala 50:65:@7460.4]
  assign _T_9494 = _T_9488[5]; // @[Bitwise.scala 50:65:@7461.4]
  assign _T_9495 = _T_9488[6]; // @[Bitwise.scala 50:65:@7462.4]
  assign _T_9496 = _T_9488[7]; // @[Bitwise.scala 50:65:@7463.4]
  assign _T_9497 = _T_9488[8]; // @[Bitwise.scala 50:65:@7464.4]
  assign _T_9498 = _T_9488[9]; // @[Bitwise.scala 50:65:@7465.4]
  assign _T_9499 = _T_9488[10]; // @[Bitwise.scala 50:65:@7466.4]
  assign _T_9500 = _T_9488[11]; // @[Bitwise.scala 50:65:@7467.4]
  assign _T_9501 = _T_9488[12]; // @[Bitwise.scala 50:65:@7468.4]
  assign _T_9502 = _T_9488[13]; // @[Bitwise.scala 50:65:@7469.4]
  assign _T_9503 = _T_9488[14]; // @[Bitwise.scala 50:65:@7470.4]
  assign _T_9504 = _T_9488[15]; // @[Bitwise.scala 50:65:@7471.4]
  assign _T_9505 = _T_9488[16]; // @[Bitwise.scala 50:65:@7472.4]
  assign _T_9506 = _T_9488[17]; // @[Bitwise.scala 50:65:@7473.4]
  assign _T_9507 = _T_9488[18]; // @[Bitwise.scala 50:65:@7474.4]
  assign _T_9508 = _T_9488[19]; // @[Bitwise.scala 50:65:@7475.4]
  assign _T_9509 = _T_9488[20]; // @[Bitwise.scala 50:65:@7476.4]
  assign _T_9510 = _T_9488[21]; // @[Bitwise.scala 50:65:@7477.4]
  assign _T_9511 = _T_9488[22]; // @[Bitwise.scala 50:65:@7478.4]
  assign _T_9512 = _T_9488[23]; // @[Bitwise.scala 50:65:@7479.4]
  assign _T_9513 = _T_9488[24]; // @[Bitwise.scala 50:65:@7480.4]
  assign _T_9514 = _T_9488[25]; // @[Bitwise.scala 50:65:@7481.4]
  assign _T_9515 = _T_9488[26]; // @[Bitwise.scala 50:65:@7482.4]
  assign _T_9516 = _T_9488[27]; // @[Bitwise.scala 50:65:@7483.4]
  assign _T_9517 = _T_9488[28]; // @[Bitwise.scala 50:65:@7484.4]
  assign _T_9518 = _T_9488[29]; // @[Bitwise.scala 50:65:@7485.4]
  assign _T_9519 = _T_9488[30]; // @[Bitwise.scala 50:65:@7486.4]
  assign _T_9520 = _T_9488[31]; // @[Bitwise.scala 50:65:@7487.4]
  assign _T_9521 = _T_9488[32]; // @[Bitwise.scala 50:65:@7488.4]
  assign _T_9522 = _T_9488[33]; // @[Bitwise.scala 50:65:@7489.4]
  assign _T_9523 = _T_9488[34]; // @[Bitwise.scala 50:65:@7490.4]
  assign _T_9524 = _T_9488[35]; // @[Bitwise.scala 50:65:@7491.4]
  assign _T_9525 = _T_9488[36]; // @[Bitwise.scala 50:65:@7492.4]
  assign _T_9526 = _T_9488[37]; // @[Bitwise.scala 50:65:@7493.4]
  assign _T_9527 = _T_9488[38]; // @[Bitwise.scala 50:65:@7494.4]
  assign _T_9528 = _T_9488[39]; // @[Bitwise.scala 50:65:@7495.4]
  assign _T_9529 = _T_9488[40]; // @[Bitwise.scala 50:65:@7496.4]
  assign _T_9530 = _T_9488[41]; // @[Bitwise.scala 50:65:@7497.4]
  assign _T_9531 = _T_9488[42]; // @[Bitwise.scala 50:65:@7498.4]
  assign _T_9532 = _T_9488[43]; // @[Bitwise.scala 50:65:@7499.4]
  assign _T_9533 = _T_9488[44]; // @[Bitwise.scala 50:65:@7500.4]
  assign _T_9534 = _T_9488[45]; // @[Bitwise.scala 50:65:@7501.4]
  assign _T_9535 = _T_9488[46]; // @[Bitwise.scala 50:65:@7502.4]
  assign _T_9536 = _T_9488[47]; // @[Bitwise.scala 50:65:@7503.4]
  assign _T_9537 = _T_9488[48]; // @[Bitwise.scala 50:65:@7504.4]
  assign _T_9538 = _T_9488[49]; // @[Bitwise.scala 50:65:@7505.4]
  assign _T_9539 = _T_9488[50]; // @[Bitwise.scala 50:65:@7506.4]
  assign _T_9540 = _T_9488[51]; // @[Bitwise.scala 50:65:@7507.4]
  assign _T_9541 = _T_9488[52]; // @[Bitwise.scala 50:65:@7508.4]
  assign _T_9542 = _T_9488[53]; // @[Bitwise.scala 50:65:@7509.4]
  assign _T_9543 = _T_9488[54]; // @[Bitwise.scala 50:65:@7510.4]
  assign _T_9544 = _T_9488[55]; // @[Bitwise.scala 50:65:@7511.4]
  assign _T_9545 = _T_9488[56]; // @[Bitwise.scala 50:65:@7512.4]
  assign _T_9546 = _T_9488[57]; // @[Bitwise.scala 50:65:@7513.4]
  assign _T_9547 = _T_9488[58]; // @[Bitwise.scala 50:65:@7514.4]
  assign _T_9548 = _T_9488[59]; // @[Bitwise.scala 50:65:@7515.4]
  assign _T_9549 = _T_9490 + _T_9491; // @[Bitwise.scala 48:55:@7516.4]
  assign _GEN_987 = {{1'd0}, _T_9489}; // @[Bitwise.scala 48:55:@7517.4]
  assign _T_9550 = _GEN_987 + _T_9549; // @[Bitwise.scala 48:55:@7517.4]
  assign _T_9551 = _T_9492 + _T_9493; // @[Bitwise.scala 48:55:@7518.4]
  assign _T_9552 = _T_9494 + _T_9495; // @[Bitwise.scala 48:55:@7519.4]
  assign _T_9553 = _T_9551 + _T_9552; // @[Bitwise.scala 48:55:@7520.4]
  assign _T_9554 = _T_9550 + _T_9553; // @[Bitwise.scala 48:55:@7521.4]
  assign _T_9555 = _T_9496 + _T_9497; // @[Bitwise.scala 48:55:@7522.4]
  assign _T_9556 = _T_9498 + _T_9499; // @[Bitwise.scala 48:55:@7523.4]
  assign _T_9557 = _T_9555 + _T_9556; // @[Bitwise.scala 48:55:@7524.4]
  assign _T_9558 = _T_9500 + _T_9501; // @[Bitwise.scala 48:55:@7525.4]
  assign _T_9559 = _T_9502 + _T_9503; // @[Bitwise.scala 48:55:@7526.4]
  assign _T_9560 = _T_9558 + _T_9559; // @[Bitwise.scala 48:55:@7527.4]
  assign _T_9561 = _T_9557 + _T_9560; // @[Bitwise.scala 48:55:@7528.4]
  assign _T_9562 = _T_9554 + _T_9561; // @[Bitwise.scala 48:55:@7529.4]
  assign _T_9563 = _T_9505 + _T_9506; // @[Bitwise.scala 48:55:@7530.4]
  assign _GEN_988 = {{1'd0}, _T_9504}; // @[Bitwise.scala 48:55:@7531.4]
  assign _T_9564 = _GEN_988 + _T_9563; // @[Bitwise.scala 48:55:@7531.4]
  assign _T_9565 = _T_9507 + _T_9508; // @[Bitwise.scala 48:55:@7532.4]
  assign _T_9566 = _T_9509 + _T_9510; // @[Bitwise.scala 48:55:@7533.4]
  assign _T_9567 = _T_9565 + _T_9566; // @[Bitwise.scala 48:55:@7534.4]
  assign _T_9568 = _T_9564 + _T_9567; // @[Bitwise.scala 48:55:@7535.4]
  assign _T_9569 = _T_9511 + _T_9512; // @[Bitwise.scala 48:55:@7536.4]
  assign _T_9570 = _T_9513 + _T_9514; // @[Bitwise.scala 48:55:@7537.4]
  assign _T_9571 = _T_9569 + _T_9570; // @[Bitwise.scala 48:55:@7538.4]
  assign _T_9572 = _T_9515 + _T_9516; // @[Bitwise.scala 48:55:@7539.4]
  assign _T_9573 = _T_9517 + _T_9518; // @[Bitwise.scala 48:55:@7540.4]
  assign _T_9574 = _T_9572 + _T_9573; // @[Bitwise.scala 48:55:@7541.4]
  assign _T_9575 = _T_9571 + _T_9574; // @[Bitwise.scala 48:55:@7542.4]
  assign _T_9576 = _T_9568 + _T_9575; // @[Bitwise.scala 48:55:@7543.4]
  assign _T_9577 = _T_9562 + _T_9576; // @[Bitwise.scala 48:55:@7544.4]
  assign _T_9578 = _T_9520 + _T_9521; // @[Bitwise.scala 48:55:@7545.4]
  assign _GEN_989 = {{1'd0}, _T_9519}; // @[Bitwise.scala 48:55:@7546.4]
  assign _T_9579 = _GEN_989 + _T_9578; // @[Bitwise.scala 48:55:@7546.4]
  assign _T_9580 = _T_9522 + _T_9523; // @[Bitwise.scala 48:55:@7547.4]
  assign _T_9581 = _T_9524 + _T_9525; // @[Bitwise.scala 48:55:@7548.4]
  assign _T_9582 = _T_9580 + _T_9581; // @[Bitwise.scala 48:55:@7549.4]
  assign _T_9583 = _T_9579 + _T_9582; // @[Bitwise.scala 48:55:@7550.4]
  assign _T_9584 = _T_9526 + _T_9527; // @[Bitwise.scala 48:55:@7551.4]
  assign _T_9585 = _T_9528 + _T_9529; // @[Bitwise.scala 48:55:@7552.4]
  assign _T_9586 = _T_9584 + _T_9585; // @[Bitwise.scala 48:55:@7553.4]
  assign _T_9587 = _T_9530 + _T_9531; // @[Bitwise.scala 48:55:@7554.4]
  assign _T_9588 = _T_9532 + _T_9533; // @[Bitwise.scala 48:55:@7555.4]
  assign _T_9589 = _T_9587 + _T_9588; // @[Bitwise.scala 48:55:@7556.4]
  assign _T_9590 = _T_9586 + _T_9589; // @[Bitwise.scala 48:55:@7557.4]
  assign _T_9591 = _T_9583 + _T_9590; // @[Bitwise.scala 48:55:@7558.4]
  assign _T_9592 = _T_9535 + _T_9536; // @[Bitwise.scala 48:55:@7559.4]
  assign _GEN_990 = {{1'd0}, _T_9534}; // @[Bitwise.scala 48:55:@7560.4]
  assign _T_9593 = _GEN_990 + _T_9592; // @[Bitwise.scala 48:55:@7560.4]
  assign _T_9594 = _T_9537 + _T_9538; // @[Bitwise.scala 48:55:@7561.4]
  assign _T_9595 = _T_9539 + _T_9540; // @[Bitwise.scala 48:55:@7562.4]
  assign _T_9596 = _T_9594 + _T_9595; // @[Bitwise.scala 48:55:@7563.4]
  assign _T_9597 = _T_9593 + _T_9596; // @[Bitwise.scala 48:55:@7564.4]
  assign _T_9598 = _T_9541 + _T_9542; // @[Bitwise.scala 48:55:@7565.4]
  assign _T_9599 = _T_9543 + _T_9544; // @[Bitwise.scala 48:55:@7566.4]
  assign _T_9600 = _T_9598 + _T_9599; // @[Bitwise.scala 48:55:@7567.4]
  assign _T_9601 = _T_9545 + _T_9546; // @[Bitwise.scala 48:55:@7568.4]
  assign _T_9602 = _T_9547 + _T_9548; // @[Bitwise.scala 48:55:@7569.4]
  assign _T_9603 = _T_9601 + _T_9602; // @[Bitwise.scala 48:55:@7570.4]
  assign _T_9604 = _T_9600 + _T_9603; // @[Bitwise.scala 48:55:@7571.4]
  assign _T_9605 = _T_9597 + _T_9604; // @[Bitwise.scala 48:55:@7572.4]
  assign _T_9606 = _T_9591 + _T_9605; // @[Bitwise.scala 48:55:@7573.4]
  assign _T_9607 = _T_9577 + _T_9606; // @[Bitwise.scala 48:55:@7574.4]
  assign _T_9671 = _T_2230[60:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7639.4]
  assign _T_9672 = _T_9671[0]; // @[Bitwise.scala 50:65:@7640.4]
  assign _T_9673 = _T_9671[1]; // @[Bitwise.scala 50:65:@7641.4]
  assign _T_9674 = _T_9671[2]; // @[Bitwise.scala 50:65:@7642.4]
  assign _T_9675 = _T_9671[3]; // @[Bitwise.scala 50:65:@7643.4]
  assign _T_9676 = _T_9671[4]; // @[Bitwise.scala 50:65:@7644.4]
  assign _T_9677 = _T_9671[5]; // @[Bitwise.scala 50:65:@7645.4]
  assign _T_9678 = _T_9671[6]; // @[Bitwise.scala 50:65:@7646.4]
  assign _T_9679 = _T_9671[7]; // @[Bitwise.scala 50:65:@7647.4]
  assign _T_9680 = _T_9671[8]; // @[Bitwise.scala 50:65:@7648.4]
  assign _T_9681 = _T_9671[9]; // @[Bitwise.scala 50:65:@7649.4]
  assign _T_9682 = _T_9671[10]; // @[Bitwise.scala 50:65:@7650.4]
  assign _T_9683 = _T_9671[11]; // @[Bitwise.scala 50:65:@7651.4]
  assign _T_9684 = _T_9671[12]; // @[Bitwise.scala 50:65:@7652.4]
  assign _T_9685 = _T_9671[13]; // @[Bitwise.scala 50:65:@7653.4]
  assign _T_9686 = _T_9671[14]; // @[Bitwise.scala 50:65:@7654.4]
  assign _T_9687 = _T_9671[15]; // @[Bitwise.scala 50:65:@7655.4]
  assign _T_9688 = _T_9671[16]; // @[Bitwise.scala 50:65:@7656.4]
  assign _T_9689 = _T_9671[17]; // @[Bitwise.scala 50:65:@7657.4]
  assign _T_9690 = _T_9671[18]; // @[Bitwise.scala 50:65:@7658.4]
  assign _T_9691 = _T_9671[19]; // @[Bitwise.scala 50:65:@7659.4]
  assign _T_9692 = _T_9671[20]; // @[Bitwise.scala 50:65:@7660.4]
  assign _T_9693 = _T_9671[21]; // @[Bitwise.scala 50:65:@7661.4]
  assign _T_9694 = _T_9671[22]; // @[Bitwise.scala 50:65:@7662.4]
  assign _T_9695 = _T_9671[23]; // @[Bitwise.scala 50:65:@7663.4]
  assign _T_9696 = _T_9671[24]; // @[Bitwise.scala 50:65:@7664.4]
  assign _T_9697 = _T_9671[25]; // @[Bitwise.scala 50:65:@7665.4]
  assign _T_9698 = _T_9671[26]; // @[Bitwise.scala 50:65:@7666.4]
  assign _T_9699 = _T_9671[27]; // @[Bitwise.scala 50:65:@7667.4]
  assign _T_9700 = _T_9671[28]; // @[Bitwise.scala 50:65:@7668.4]
  assign _T_9701 = _T_9671[29]; // @[Bitwise.scala 50:65:@7669.4]
  assign _T_9702 = _T_9671[30]; // @[Bitwise.scala 50:65:@7670.4]
  assign _T_9703 = _T_9671[31]; // @[Bitwise.scala 50:65:@7671.4]
  assign _T_9704 = _T_9671[32]; // @[Bitwise.scala 50:65:@7672.4]
  assign _T_9705 = _T_9671[33]; // @[Bitwise.scala 50:65:@7673.4]
  assign _T_9706 = _T_9671[34]; // @[Bitwise.scala 50:65:@7674.4]
  assign _T_9707 = _T_9671[35]; // @[Bitwise.scala 50:65:@7675.4]
  assign _T_9708 = _T_9671[36]; // @[Bitwise.scala 50:65:@7676.4]
  assign _T_9709 = _T_9671[37]; // @[Bitwise.scala 50:65:@7677.4]
  assign _T_9710 = _T_9671[38]; // @[Bitwise.scala 50:65:@7678.4]
  assign _T_9711 = _T_9671[39]; // @[Bitwise.scala 50:65:@7679.4]
  assign _T_9712 = _T_9671[40]; // @[Bitwise.scala 50:65:@7680.4]
  assign _T_9713 = _T_9671[41]; // @[Bitwise.scala 50:65:@7681.4]
  assign _T_9714 = _T_9671[42]; // @[Bitwise.scala 50:65:@7682.4]
  assign _T_9715 = _T_9671[43]; // @[Bitwise.scala 50:65:@7683.4]
  assign _T_9716 = _T_9671[44]; // @[Bitwise.scala 50:65:@7684.4]
  assign _T_9717 = _T_9671[45]; // @[Bitwise.scala 50:65:@7685.4]
  assign _T_9718 = _T_9671[46]; // @[Bitwise.scala 50:65:@7686.4]
  assign _T_9719 = _T_9671[47]; // @[Bitwise.scala 50:65:@7687.4]
  assign _T_9720 = _T_9671[48]; // @[Bitwise.scala 50:65:@7688.4]
  assign _T_9721 = _T_9671[49]; // @[Bitwise.scala 50:65:@7689.4]
  assign _T_9722 = _T_9671[50]; // @[Bitwise.scala 50:65:@7690.4]
  assign _T_9723 = _T_9671[51]; // @[Bitwise.scala 50:65:@7691.4]
  assign _T_9724 = _T_9671[52]; // @[Bitwise.scala 50:65:@7692.4]
  assign _T_9725 = _T_9671[53]; // @[Bitwise.scala 50:65:@7693.4]
  assign _T_9726 = _T_9671[54]; // @[Bitwise.scala 50:65:@7694.4]
  assign _T_9727 = _T_9671[55]; // @[Bitwise.scala 50:65:@7695.4]
  assign _T_9728 = _T_9671[56]; // @[Bitwise.scala 50:65:@7696.4]
  assign _T_9729 = _T_9671[57]; // @[Bitwise.scala 50:65:@7697.4]
  assign _T_9730 = _T_9671[58]; // @[Bitwise.scala 50:65:@7698.4]
  assign _T_9731 = _T_9671[59]; // @[Bitwise.scala 50:65:@7699.4]
  assign _T_9732 = _T_9671[60]; // @[Bitwise.scala 50:65:@7700.4]
  assign _T_9733 = _T_9673 + _T_9674; // @[Bitwise.scala 48:55:@7701.4]
  assign _GEN_991 = {{1'd0}, _T_9672}; // @[Bitwise.scala 48:55:@7702.4]
  assign _T_9734 = _GEN_991 + _T_9733; // @[Bitwise.scala 48:55:@7702.4]
  assign _T_9735 = _T_9675 + _T_9676; // @[Bitwise.scala 48:55:@7703.4]
  assign _T_9736 = _T_9677 + _T_9678; // @[Bitwise.scala 48:55:@7704.4]
  assign _T_9737 = _T_9735 + _T_9736; // @[Bitwise.scala 48:55:@7705.4]
  assign _T_9738 = _T_9734 + _T_9737; // @[Bitwise.scala 48:55:@7706.4]
  assign _T_9739 = _T_9679 + _T_9680; // @[Bitwise.scala 48:55:@7707.4]
  assign _T_9740 = _T_9681 + _T_9682; // @[Bitwise.scala 48:55:@7708.4]
  assign _T_9741 = _T_9739 + _T_9740; // @[Bitwise.scala 48:55:@7709.4]
  assign _T_9742 = _T_9683 + _T_9684; // @[Bitwise.scala 48:55:@7710.4]
  assign _T_9743 = _T_9685 + _T_9686; // @[Bitwise.scala 48:55:@7711.4]
  assign _T_9744 = _T_9742 + _T_9743; // @[Bitwise.scala 48:55:@7712.4]
  assign _T_9745 = _T_9741 + _T_9744; // @[Bitwise.scala 48:55:@7713.4]
  assign _T_9746 = _T_9738 + _T_9745; // @[Bitwise.scala 48:55:@7714.4]
  assign _T_9747 = _T_9688 + _T_9689; // @[Bitwise.scala 48:55:@7715.4]
  assign _GEN_992 = {{1'd0}, _T_9687}; // @[Bitwise.scala 48:55:@7716.4]
  assign _T_9748 = _GEN_992 + _T_9747; // @[Bitwise.scala 48:55:@7716.4]
  assign _T_9749 = _T_9690 + _T_9691; // @[Bitwise.scala 48:55:@7717.4]
  assign _T_9750 = _T_9692 + _T_9693; // @[Bitwise.scala 48:55:@7718.4]
  assign _T_9751 = _T_9749 + _T_9750; // @[Bitwise.scala 48:55:@7719.4]
  assign _T_9752 = _T_9748 + _T_9751; // @[Bitwise.scala 48:55:@7720.4]
  assign _T_9753 = _T_9694 + _T_9695; // @[Bitwise.scala 48:55:@7721.4]
  assign _T_9754 = _T_9696 + _T_9697; // @[Bitwise.scala 48:55:@7722.4]
  assign _T_9755 = _T_9753 + _T_9754; // @[Bitwise.scala 48:55:@7723.4]
  assign _T_9756 = _T_9698 + _T_9699; // @[Bitwise.scala 48:55:@7724.4]
  assign _T_9757 = _T_9700 + _T_9701; // @[Bitwise.scala 48:55:@7725.4]
  assign _T_9758 = _T_9756 + _T_9757; // @[Bitwise.scala 48:55:@7726.4]
  assign _T_9759 = _T_9755 + _T_9758; // @[Bitwise.scala 48:55:@7727.4]
  assign _T_9760 = _T_9752 + _T_9759; // @[Bitwise.scala 48:55:@7728.4]
  assign _T_9761 = _T_9746 + _T_9760; // @[Bitwise.scala 48:55:@7729.4]
  assign _T_9762 = _T_9703 + _T_9704; // @[Bitwise.scala 48:55:@7730.4]
  assign _GEN_993 = {{1'd0}, _T_9702}; // @[Bitwise.scala 48:55:@7731.4]
  assign _T_9763 = _GEN_993 + _T_9762; // @[Bitwise.scala 48:55:@7731.4]
  assign _T_9764 = _T_9705 + _T_9706; // @[Bitwise.scala 48:55:@7732.4]
  assign _T_9765 = _T_9707 + _T_9708; // @[Bitwise.scala 48:55:@7733.4]
  assign _T_9766 = _T_9764 + _T_9765; // @[Bitwise.scala 48:55:@7734.4]
  assign _T_9767 = _T_9763 + _T_9766; // @[Bitwise.scala 48:55:@7735.4]
  assign _T_9768 = _T_9709 + _T_9710; // @[Bitwise.scala 48:55:@7736.4]
  assign _T_9769 = _T_9711 + _T_9712; // @[Bitwise.scala 48:55:@7737.4]
  assign _T_9770 = _T_9768 + _T_9769; // @[Bitwise.scala 48:55:@7738.4]
  assign _T_9771 = _T_9713 + _T_9714; // @[Bitwise.scala 48:55:@7739.4]
  assign _T_9772 = _T_9715 + _T_9716; // @[Bitwise.scala 48:55:@7740.4]
  assign _T_9773 = _T_9771 + _T_9772; // @[Bitwise.scala 48:55:@7741.4]
  assign _T_9774 = _T_9770 + _T_9773; // @[Bitwise.scala 48:55:@7742.4]
  assign _T_9775 = _T_9767 + _T_9774; // @[Bitwise.scala 48:55:@7743.4]
  assign _T_9776 = _T_9717 + _T_9718; // @[Bitwise.scala 48:55:@7744.4]
  assign _T_9777 = _T_9719 + _T_9720; // @[Bitwise.scala 48:55:@7745.4]
  assign _T_9778 = _T_9776 + _T_9777; // @[Bitwise.scala 48:55:@7746.4]
  assign _T_9779 = _T_9721 + _T_9722; // @[Bitwise.scala 48:55:@7747.4]
  assign _T_9780 = _T_9723 + _T_9724; // @[Bitwise.scala 48:55:@7748.4]
  assign _T_9781 = _T_9779 + _T_9780; // @[Bitwise.scala 48:55:@7749.4]
  assign _T_9782 = _T_9778 + _T_9781; // @[Bitwise.scala 48:55:@7750.4]
  assign _T_9783 = _T_9725 + _T_9726; // @[Bitwise.scala 48:55:@7751.4]
  assign _T_9784 = _T_9727 + _T_9728; // @[Bitwise.scala 48:55:@7752.4]
  assign _T_9785 = _T_9783 + _T_9784; // @[Bitwise.scala 48:55:@7753.4]
  assign _T_9786 = _T_9729 + _T_9730; // @[Bitwise.scala 48:55:@7754.4]
  assign _T_9787 = _T_9731 + _T_9732; // @[Bitwise.scala 48:55:@7755.4]
  assign _T_9788 = _T_9786 + _T_9787; // @[Bitwise.scala 48:55:@7756.4]
  assign _T_9789 = _T_9785 + _T_9788; // @[Bitwise.scala 48:55:@7757.4]
  assign _T_9790 = _T_9782 + _T_9789; // @[Bitwise.scala 48:55:@7758.4]
  assign _T_9791 = _T_9775 + _T_9790; // @[Bitwise.scala 48:55:@7759.4]
  assign _T_9792 = _T_9761 + _T_9791; // @[Bitwise.scala 48:55:@7760.4]
  assign _T_9856 = _T_2230[61:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@7825.4]
  assign _T_9857 = _T_9856[0]; // @[Bitwise.scala 50:65:@7826.4]
  assign _T_9858 = _T_9856[1]; // @[Bitwise.scala 50:65:@7827.4]
  assign _T_9859 = _T_9856[2]; // @[Bitwise.scala 50:65:@7828.4]
  assign _T_9860 = _T_9856[3]; // @[Bitwise.scala 50:65:@7829.4]
  assign _T_9861 = _T_9856[4]; // @[Bitwise.scala 50:65:@7830.4]
  assign _T_9862 = _T_9856[5]; // @[Bitwise.scala 50:65:@7831.4]
  assign _T_9863 = _T_9856[6]; // @[Bitwise.scala 50:65:@7832.4]
  assign _T_9864 = _T_9856[7]; // @[Bitwise.scala 50:65:@7833.4]
  assign _T_9865 = _T_9856[8]; // @[Bitwise.scala 50:65:@7834.4]
  assign _T_9866 = _T_9856[9]; // @[Bitwise.scala 50:65:@7835.4]
  assign _T_9867 = _T_9856[10]; // @[Bitwise.scala 50:65:@7836.4]
  assign _T_9868 = _T_9856[11]; // @[Bitwise.scala 50:65:@7837.4]
  assign _T_9869 = _T_9856[12]; // @[Bitwise.scala 50:65:@7838.4]
  assign _T_9870 = _T_9856[13]; // @[Bitwise.scala 50:65:@7839.4]
  assign _T_9871 = _T_9856[14]; // @[Bitwise.scala 50:65:@7840.4]
  assign _T_9872 = _T_9856[15]; // @[Bitwise.scala 50:65:@7841.4]
  assign _T_9873 = _T_9856[16]; // @[Bitwise.scala 50:65:@7842.4]
  assign _T_9874 = _T_9856[17]; // @[Bitwise.scala 50:65:@7843.4]
  assign _T_9875 = _T_9856[18]; // @[Bitwise.scala 50:65:@7844.4]
  assign _T_9876 = _T_9856[19]; // @[Bitwise.scala 50:65:@7845.4]
  assign _T_9877 = _T_9856[20]; // @[Bitwise.scala 50:65:@7846.4]
  assign _T_9878 = _T_9856[21]; // @[Bitwise.scala 50:65:@7847.4]
  assign _T_9879 = _T_9856[22]; // @[Bitwise.scala 50:65:@7848.4]
  assign _T_9880 = _T_9856[23]; // @[Bitwise.scala 50:65:@7849.4]
  assign _T_9881 = _T_9856[24]; // @[Bitwise.scala 50:65:@7850.4]
  assign _T_9882 = _T_9856[25]; // @[Bitwise.scala 50:65:@7851.4]
  assign _T_9883 = _T_9856[26]; // @[Bitwise.scala 50:65:@7852.4]
  assign _T_9884 = _T_9856[27]; // @[Bitwise.scala 50:65:@7853.4]
  assign _T_9885 = _T_9856[28]; // @[Bitwise.scala 50:65:@7854.4]
  assign _T_9886 = _T_9856[29]; // @[Bitwise.scala 50:65:@7855.4]
  assign _T_9887 = _T_9856[30]; // @[Bitwise.scala 50:65:@7856.4]
  assign _T_9888 = _T_9856[31]; // @[Bitwise.scala 50:65:@7857.4]
  assign _T_9889 = _T_9856[32]; // @[Bitwise.scala 50:65:@7858.4]
  assign _T_9890 = _T_9856[33]; // @[Bitwise.scala 50:65:@7859.4]
  assign _T_9891 = _T_9856[34]; // @[Bitwise.scala 50:65:@7860.4]
  assign _T_9892 = _T_9856[35]; // @[Bitwise.scala 50:65:@7861.4]
  assign _T_9893 = _T_9856[36]; // @[Bitwise.scala 50:65:@7862.4]
  assign _T_9894 = _T_9856[37]; // @[Bitwise.scala 50:65:@7863.4]
  assign _T_9895 = _T_9856[38]; // @[Bitwise.scala 50:65:@7864.4]
  assign _T_9896 = _T_9856[39]; // @[Bitwise.scala 50:65:@7865.4]
  assign _T_9897 = _T_9856[40]; // @[Bitwise.scala 50:65:@7866.4]
  assign _T_9898 = _T_9856[41]; // @[Bitwise.scala 50:65:@7867.4]
  assign _T_9899 = _T_9856[42]; // @[Bitwise.scala 50:65:@7868.4]
  assign _T_9900 = _T_9856[43]; // @[Bitwise.scala 50:65:@7869.4]
  assign _T_9901 = _T_9856[44]; // @[Bitwise.scala 50:65:@7870.4]
  assign _T_9902 = _T_9856[45]; // @[Bitwise.scala 50:65:@7871.4]
  assign _T_9903 = _T_9856[46]; // @[Bitwise.scala 50:65:@7872.4]
  assign _T_9904 = _T_9856[47]; // @[Bitwise.scala 50:65:@7873.4]
  assign _T_9905 = _T_9856[48]; // @[Bitwise.scala 50:65:@7874.4]
  assign _T_9906 = _T_9856[49]; // @[Bitwise.scala 50:65:@7875.4]
  assign _T_9907 = _T_9856[50]; // @[Bitwise.scala 50:65:@7876.4]
  assign _T_9908 = _T_9856[51]; // @[Bitwise.scala 50:65:@7877.4]
  assign _T_9909 = _T_9856[52]; // @[Bitwise.scala 50:65:@7878.4]
  assign _T_9910 = _T_9856[53]; // @[Bitwise.scala 50:65:@7879.4]
  assign _T_9911 = _T_9856[54]; // @[Bitwise.scala 50:65:@7880.4]
  assign _T_9912 = _T_9856[55]; // @[Bitwise.scala 50:65:@7881.4]
  assign _T_9913 = _T_9856[56]; // @[Bitwise.scala 50:65:@7882.4]
  assign _T_9914 = _T_9856[57]; // @[Bitwise.scala 50:65:@7883.4]
  assign _T_9915 = _T_9856[58]; // @[Bitwise.scala 50:65:@7884.4]
  assign _T_9916 = _T_9856[59]; // @[Bitwise.scala 50:65:@7885.4]
  assign _T_9917 = _T_9856[60]; // @[Bitwise.scala 50:65:@7886.4]
  assign _T_9918 = _T_9856[61]; // @[Bitwise.scala 50:65:@7887.4]
  assign _T_9919 = _T_9858 + _T_9859; // @[Bitwise.scala 48:55:@7888.4]
  assign _GEN_994 = {{1'd0}, _T_9857}; // @[Bitwise.scala 48:55:@7889.4]
  assign _T_9920 = _GEN_994 + _T_9919; // @[Bitwise.scala 48:55:@7889.4]
  assign _T_9921 = _T_9860 + _T_9861; // @[Bitwise.scala 48:55:@7890.4]
  assign _T_9922 = _T_9862 + _T_9863; // @[Bitwise.scala 48:55:@7891.4]
  assign _T_9923 = _T_9921 + _T_9922; // @[Bitwise.scala 48:55:@7892.4]
  assign _T_9924 = _T_9920 + _T_9923; // @[Bitwise.scala 48:55:@7893.4]
  assign _T_9925 = _T_9864 + _T_9865; // @[Bitwise.scala 48:55:@7894.4]
  assign _T_9926 = _T_9866 + _T_9867; // @[Bitwise.scala 48:55:@7895.4]
  assign _T_9927 = _T_9925 + _T_9926; // @[Bitwise.scala 48:55:@7896.4]
  assign _T_9928 = _T_9868 + _T_9869; // @[Bitwise.scala 48:55:@7897.4]
  assign _T_9929 = _T_9870 + _T_9871; // @[Bitwise.scala 48:55:@7898.4]
  assign _T_9930 = _T_9928 + _T_9929; // @[Bitwise.scala 48:55:@7899.4]
  assign _T_9931 = _T_9927 + _T_9930; // @[Bitwise.scala 48:55:@7900.4]
  assign _T_9932 = _T_9924 + _T_9931; // @[Bitwise.scala 48:55:@7901.4]
  assign _T_9933 = _T_9872 + _T_9873; // @[Bitwise.scala 48:55:@7902.4]
  assign _T_9934 = _T_9874 + _T_9875; // @[Bitwise.scala 48:55:@7903.4]
  assign _T_9935 = _T_9933 + _T_9934; // @[Bitwise.scala 48:55:@7904.4]
  assign _T_9936 = _T_9876 + _T_9877; // @[Bitwise.scala 48:55:@7905.4]
  assign _T_9937 = _T_9878 + _T_9879; // @[Bitwise.scala 48:55:@7906.4]
  assign _T_9938 = _T_9936 + _T_9937; // @[Bitwise.scala 48:55:@7907.4]
  assign _T_9939 = _T_9935 + _T_9938; // @[Bitwise.scala 48:55:@7908.4]
  assign _T_9940 = _T_9880 + _T_9881; // @[Bitwise.scala 48:55:@7909.4]
  assign _T_9941 = _T_9882 + _T_9883; // @[Bitwise.scala 48:55:@7910.4]
  assign _T_9942 = _T_9940 + _T_9941; // @[Bitwise.scala 48:55:@7911.4]
  assign _T_9943 = _T_9884 + _T_9885; // @[Bitwise.scala 48:55:@7912.4]
  assign _T_9944 = _T_9886 + _T_9887; // @[Bitwise.scala 48:55:@7913.4]
  assign _T_9945 = _T_9943 + _T_9944; // @[Bitwise.scala 48:55:@7914.4]
  assign _T_9946 = _T_9942 + _T_9945; // @[Bitwise.scala 48:55:@7915.4]
  assign _T_9947 = _T_9939 + _T_9946; // @[Bitwise.scala 48:55:@7916.4]
  assign _T_9948 = _T_9932 + _T_9947; // @[Bitwise.scala 48:55:@7917.4]
  assign _T_9949 = _T_9889 + _T_9890; // @[Bitwise.scala 48:55:@7918.4]
  assign _GEN_995 = {{1'd0}, _T_9888}; // @[Bitwise.scala 48:55:@7919.4]
  assign _T_9950 = _GEN_995 + _T_9949; // @[Bitwise.scala 48:55:@7919.4]
  assign _T_9951 = _T_9891 + _T_9892; // @[Bitwise.scala 48:55:@7920.4]
  assign _T_9952 = _T_9893 + _T_9894; // @[Bitwise.scala 48:55:@7921.4]
  assign _T_9953 = _T_9951 + _T_9952; // @[Bitwise.scala 48:55:@7922.4]
  assign _T_9954 = _T_9950 + _T_9953; // @[Bitwise.scala 48:55:@7923.4]
  assign _T_9955 = _T_9895 + _T_9896; // @[Bitwise.scala 48:55:@7924.4]
  assign _T_9956 = _T_9897 + _T_9898; // @[Bitwise.scala 48:55:@7925.4]
  assign _T_9957 = _T_9955 + _T_9956; // @[Bitwise.scala 48:55:@7926.4]
  assign _T_9958 = _T_9899 + _T_9900; // @[Bitwise.scala 48:55:@7927.4]
  assign _T_9959 = _T_9901 + _T_9902; // @[Bitwise.scala 48:55:@7928.4]
  assign _T_9960 = _T_9958 + _T_9959; // @[Bitwise.scala 48:55:@7929.4]
  assign _T_9961 = _T_9957 + _T_9960; // @[Bitwise.scala 48:55:@7930.4]
  assign _T_9962 = _T_9954 + _T_9961; // @[Bitwise.scala 48:55:@7931.4]
  assign _T_9963 = _T_9903 + _T_9904; // @[Bitwise.scala 48:55:@7932.4]
  assign _T_9964 = _T_9905 + _T_9906; // @[Bitwise.scala 48:55:@7933.4]
  assign _T_9965 = _T_9963 + _T_9964; // @[Bitwise.scala 48:55:@7934.4]
  assign _T_9966 = _T_9907 + _T_9908; // @[Bitwise.scala 48:55:@7935.4]
  assign _T_9967 = _T_9909 + _T_9910; // @[Bitwise.scala 48:55:@7936.4]
  assign _T_9968 = _T_9966 + _T_9967; // @[Bitwise.scala 48:55:@7937.4]
  assign _T_9969 = _T_9965 + _T_9968; // @[Bitwise.scala 48:55:@7938.4]
  assign _T_9970 = _T_9911 + _T_9912; // @[Bitwise.scala 48:55:@7939.4]
  assign _T_9971 = _T_9913 + _T_9914; // @[Bitwise.scala 48:55:@7940.4]
  assign _T_9972 = _T_9970 + _T_9971; // @[Bitwise.scala 48:55:@7941.4]
  assign _T_9973 = _T_9915 + _T_9916; // @[Bitwise.scala 48:55:@7942.4]
  assign _T_9974 = _T_9917 + _T_9918; // @[Bitwise.scala 48:55:@7943.4]
  assign _T_9975 = _T_9973 + _T_9974; // @[Bitwise.scala 48:55:@7944.4]
  assign _T_9976 = _T_9972 + _T_9975; // @[Bitwise.scala 48:55:@7945.4]
  assign _T_9977 = _T_9969 + _T_9976; // @[Bitwise.scala 48:55:@7946.4]
  assign _T_9978 = _T_9962 + _T_9977; // @[Bitwise.scala 48:55:@7947.4]
  assign _T_9979 = _T_9948 + _T_9978; // @[Bitwise.scala 48:55:@7948.4]
  assign _T_10043 = _T_2230[62:0]; // @[NV_NVDLA_CSC_WL_dec.scala 60:60:@8013.4]
  assign _T_10044 = _T_10043[0]; // @[Bitwise.scala 50:65:@8014.4]
  assign _T_10045 = _T_10043[1]; // @[Bitwise.scala 50:65:@8015.4]
  assign _T_10046 = _T_10043[2]; // @[Bitwise.scala 50:65:@8016.4]
  assign _T_10047 = _T_10043[3]; // @[Bitwise.scala 50:65:@8017.4]
  assign _T_10048 = _T_10043[4]; // @[Bitwise.scala 50:65:@8018.4]
  assign _T_10049 = _T_10043[5]; // @[Bitwise.scala 50:65:@8019.4]
  assign _T_10050 = _T_10043[6]; // @[Bitwise.scala 50:65:@8020.4]
  assign _T_10051 = _T_10043[7]; // @[Bitwise.scala 50:65:@8021.4]
  assign _T_10052 = _T_10043[8]; // @[Bitwise.scala 50:65:@8022.4]
  assign _T_10053 = _T_10043[9]; // @[Bitwise.scala 50:65:@8023.4]
  assign _T_10054 = _T_10043[10]; // @[Bitwise.scala 50:65:@8024.4]
  assign _T_10055 = _T_10043[11]; // @[Bitwise.scala 50:65:@8025.4]
  assign _T_10056 = _T_10043[12]; // @[Bitwise.scala 50:65:@8026.4]
  assign _T_10057 = _T_10043[13]; // @[Bitwise.scala 50:65:@8027.4]
  assign _T_10058 = _T_10043[14]; // @[Bitwise.scala 50:65:@8028.4]
  assign _T_10059 = _T_10043[15]; // @[Bitwise.scala 50:65:@8029.4]
  assign _T_10060 = _T_10043[16]; // @[Bitwise.scala 50:65:@8030.4]
  assign _T_10061 = _T_10043[17]; // @[Bitwise.scala 50:65:@8031.4]
  assign _T_10062 = _T_10043[18]; // @[Bitwise.scala 50:65:@8032.4]
  assign _T_10063 = _T_10043[19]; // @[Bitwise.scala 50:65:@8033.4]
  assign _T_10064 = _T_10043[20]; // @[Bitwise.scala 50:65:@8034.4]
  assign _T_10065 = _T_10043[21]; // @[Bitwise.scala 50:65:@8035.4]
  assign _T_10066 = _T_10043[22]; // @[Bitwise.scala 50:65:@8036.4]
  assign _T_10067 = _T_10043[23]; // @[Bitwise.scala 50:65:@8037.4]
  assign _T_10068 = _T_10043[24]; // @[Bitwise.scala 50:65:@8038.4]
  assign _T_10069 = _T_10043[25]; // @[Bitwise.scala 50:65:@8039.4]
  assign _T_10070 = _T_10043[26]; // @[Bitwise.scala 50:65:@8040.4]
  assign _T_10071 = _T_10043[27]; // @[Bitwise.scala 50:65:@8041.4]
  assign _T_10072 = _T_10043[28]; // @[Bitwise.scala 50:65:@8042.4]
  assign _T_10073 = _T_10043[29]; // @[Bitwise.scala 50:65:@8043.4]
  assign _T_10074 = _T_10043[30]; // @[Bitwise.scala 50:65:@8044.4]
  assign _T_10075 = _T_10043[31]; // @[Bitwise.scala 50:65:@8045.4]
  assign _T_10076 = _T_10043[32]; // @[Bitwise.scala 50:65:@8046.4]
  assign _T_10077 = _T_10043[33]; // @[Bitwise.scala 50:65:@8047.4]
  assign _T_10078 = _T_10043[34]; // @[Bitwise.scala 50:65:@8048.4]
  assign _T_10079 = _T_10043[35]; // @[Bitwise.scala 50:65:@8049.4]
  assign _T_10080 = _T_10043[36]; // @[Bitwise.scala 50:65:@8050.4]
  assign _T_10081 = _T_10043[37]; // @[Bitwise.scala 50:65:@8051.4]
  assign _T_10082 = _T_10043[38]; // @[Bitwise.scala 50:65:@8052.4]
  assign _T_10083 = _T_10043[39]; // @[Bitwise.scala 50:65:@8053.4]
  assign _T_10084 = _T_10043[40]; // @[Bitwise.scala 50:65:@8054.4]
  assign _T_10085 = _T_10043[41]; // @[Bitwise.scala 50:65:@8055.4]
  assign _T_10086 = _T_10043[42]; // @[Bitwise.scala 50:65:@8056.4]
  assign _T_10087 = _T_10043[43]; // @[Bitwise.scala 50:65:@8057.4]
  assign _T_10088 = _T_10043[44]; // @[Bitwise.scala 50:65:@8058.4]
  assign _T_10089 = _T_10043[45]; // @[Bitwise.scala 50:65:@8059.4]
  assign _T_10090 = _T_10043[46]; // @[Bitwise.scala 50:65:@8060.4]
  assign _T_10091 = _T_10043[47]; // @[Bitwise.scala 50:65:@8061.4]
  assign _T_10092 = _T_10043[48]; // @[Bitwise.scala 50:65:@8062.4]
  assign _T_10093 = _T_10043[49]; // @[Bitwise.scala 50:65:@8063.4]
  assign _T_10094 = _T_10043[50]; // @[Bitwise.scala 50:65:@8064.4]
  assign _T_10095 = _T_10043[51]; // @[Bitwise.scala 50:65:@8065.4]
  assign _T_10096 = _T_10043[52]; // @[Bitwise.scala 50:65:@8066.4]
  assign _T_10097 = _T_10043[53]; // @[Bitwise.scala 50:65:@8067.4]
  assign _T_10098 = _T_10043[54]; // @[Bitwise.scala 50:65:@8068.4]
  assign _T_10099 = _T_10043[55]; // @[Bitwise.scala 50:65:@8069.4]
  assign _T_10100 = _T_10043[56]; // @[Bitwise.scala 50:65:@8070.4]
  assign _T_10101 = _T_10043[57]; // @[Bitwise.scala 50:65:@8071.4]
  assign _T_10102 = _T_10043[58]; // @[Bitwise.scala 50:65:@8072.4]
  assign _T_10103 = _T_10043[59]; // @[Bitwise.scala 50:65:@8073.4]
  assign _T_10104 = _T_10043[60]; // @[Bitwise.scala 50:65:@8074.4]
  assign _T_10105 = _T_10043[61]; // @[Bitwise.scala 50:65:@8075.4]
  assign _T_10106 = _T_10043[62]; // @[Bitwise.scala 50:65:@8076.4]
  assign _T_10107 = _T_10045 + _T_10046; // @[Bitwise.scala 48:55:@8077.4]
  assign _GEN_996 = {{1'd0}, _T_10044}; // @[Bitwise.scala 48:55:@8078.4]
  assign _T_10108 = _GEN_996 + _T_10107; // @[Bitwise.scala 48:55:@8078.4]
  assign _T_10109 = _T_10047 + _T_10048; // @[Bitwise.scala 48:55:@8079.4]
  assign _T_10110 = _T_10049 + _T_10050; // @[Bitwise.scala 48:55:@8080.4]
  assign _T_10111 = _T_10109 + _T_10110; // @[Bitwise.scala 48:55:@8081.4]
  assign _T_10112 = _T_10108 + _T_10111; // @[Bitwise.scala 48:55:@8082.4]
  assign _T_10113 = _T_10051 + _T_10052; // @[Bitwise.scala 48:55:@8083.4]
  assign _T_10114 = _T_10053 + _T_10054; // @[Bitwise.scala 48:55:@8084.4]
  assign _T_10115 = _T_10113 + _T_10114; // @[Bitwise.scala 48:55:@8085.4]
  assign _T_10116 = _T_10055 + _T_10056; // @[Bitwise.scala 48:55:@8086.4]
  assign _T_10117 = _T_10057 + _T_10058; // @[Bitwise.scala 48:55:@8087.4]
  assign _T_10118 = _T_10116 + _T_10117; // @[Bitwise.scala 48:55:@8088.4]
  assign _T_10119 = _T_10115 + _T_10118; // @[Bitwise.scala 48:55:@8089.4]
  assign _T_10120 = _T_10112 + _T_10119; // @[Bitwise.scala 48:55:@8090.4]
  assign _T_10121 = _T_10059 + _T_10060; // @[Bitwise.scala 48:55:@8091.4]
  assign _T_10122 = _T_10061 + _T_10062; // @[Bitwise.scala 48:55:@8092.4]
  assign _T_10123 = _T_10121 + _T_10122; // @[Bitwise.scala 48:55:@8093.4]
  assign _T_10124 = _T_10063 + _T_10064; // @[Bitwise.scala 48:55:@8094.4]
  assign _T_10125 = _T_10065 + _T_10066; // @[Bitwise.scala 48:55:@8095.4]
  assign _T_10126 = _T_10124 + _T_10125; // @[Bitwise.scala 48:55:@8096.4]
  assign _T_10127 = _T_10123 + _T_10126; // @[Bitwise.scala 48:55:@8097.4]
  assign _T_10128 = _T_10067 + _T_10068; // @[Bitwise.scala 48:55:@8098.4]
  assign _T_10129 = _T_10069 + _T_10070; // @[Bitwise.scala 48:55:@8099.4]
  assign _T_10130 = _T_10128 + _T_10129; // @[Bitwise.scala 48:55:@8100.4]
  assign _T_10131 = _T_10071 + _T_10072; // @[Bitwise.scala 48:55:@8101.4]
  assign _T_10132 = _T_10073 + _T_10074; // @[Bitwise.scala 48:55:@8102.4]
  assign _T_10133 = _T_10131 + _T_10132; // @[Bitwise.scala 48:55:@8103.4]
  assign _T_10134 = _T_10130 + _T_10133; // @[Bitwise.scala 48:55:@8104.4]
  assign _T_10135 = _T_10127 + _T_10134; // @[Bitwise.scala 48:55:@8105.4]
  assign _T_10136 = _T_10120 + _T_10135; // @[Bitwise.scala 48:55:@8106.4]
  assign _T_10137 = _T_10075 + _T_10076; // @[Bitwise.scala 48:55:@8107.4]
  assign _T_10138 = _T_10077 + _T_10078; // @[Bitwise.scala 48:55:@8108.4]
  assign _T_10139 = _T_10137 + _T_10138; // @[Bitwise.scala 48:55:@8109.4]
  assign _T_10140 = _T_10079 + _T_10080; // @[Bitwise.scala 48:55:@8110.4]
  assign _T_10141 = _T_10081 + _T_10082; // @[Bitwise.scala 48:55:@8111.4]
  assign _T_10142 = _T_10140 + _T_10141; // @[Bitwise.scala 48:55:@8112.4]
  assign _T_10143 = _T_10139 + _T_10142; // @[Bitwise.scala 48:55:@8113.4]
  assign _T_10144 = _T_10083 + _T_10084; // @[Bitwise.scala 48:55:@8114.4]
  assign _T_10145 = _T_10085 + _T_10086; // @[Bitwise.scala 48:55:@8115.4]
  assign _T_10146 = _T_10144 + _T_10145; // @[Bitwise.scala 48:55:@8116.4]
  assign _T_10147 = _T_10087 + _T_10088; // @[Bitwise.scala 48:55:@8117.4]
  assign _T_10148 = _T_10089 + _T_10090; // @[Bitwise.scala 48:55:@8118.4]
  assign _T_10149 = _T_10147 + _T_10148; // @[Bitwise.scala 48:55:@8119.4]
  assign _T_10150 = _T_10146 + _T_10149; // @[Bitwise.scala 48:55:@8120.4]
  assign _T_10151 = _T_10143 + _T_10150; // @[Bitwise.scala 48:55:@8121.4]
  assign _T_10152 = _T_10091 + _T_10092; // @[Bitwise.scala 48:55:@8122.4]
  assign _T_10153 = _T_10093 + _T_10094; // @[Bitwise.scala 48:55:@8123.4]
  assign _T_10154 = _T_10152 + _T_10153; // @[Bitwise.scala 48:55:@8124.4]
  assign _T_10155 = _T_10095 + _T_10096; // @[Bitwise.scala 48:55:@8125.4]
  assign _T_10156 = _T_10097 + _T_10098; // @[Bitwise.scala 48:55:@8126.4]
  assign _T_10157 = _T_10155 + _T_10156; // @[Bitwise.scala 48:55:@8127.4]
  assign _T_10158 = _T_10154 + _T_10157; // @[Bitwise.scala 48:55:@8128.4]
  assign _T_10159 = _T_10099 + _T_10100; // @[Bitwise.scala 48:55:@8129.4]
  assign _T_10160 = _T_10101 + _T_10102; // @[Bitwise.scala 48:55:@8130.4]
  assign _T_10161 = _T_10159 + _T_10160; // @[Bitwise.scala 48:55:@8131.4]
  assign _T_10162 = _T_10103 + _T_10104; // @[Bitwise.scala 48:55:@8132.4]
  assign _T_10163 = _T_10105 + _T_10106; // @[Bitwise.scala 48:55:@8133.4]
  assign _T_10164 = _T_10162 + _T_10163; // @[Bitwise.scala 48:55:@8134.4]
  assign _T_10165 = _T_10161 + _T_10164; // @[Bitwise.scala 48:55:@8135.4]
  assign _T_10166 = _T_10158 + _T_10165; // @[Bitwise.scala 48:55:@8136.4]
  assign _T_10167 = _T_10151 + _T_10166; // @[Bitwise.scala 48:55:@8137.4]
  assign _T_10168 = _T_10136 + _T_10167; // @[Bitwise.scala 48:55:@8138.4]
  assign _T_10234 = _T_2230[1]; // @[Bitwise.scala 50:65:@8205.4]
  assign _T_10235 = _T_2230[2]; // @[Bitwise.scala 50:65:@8206.4]
  assign _T_10236 = _T_2230[3]; // @[Bitwise.scala 50:65:@8207.4]
  assign _T_10237 = _T_2230[4]; // @[Bitwise.scala 50:65:@8208.4]
  assign _T_10238 = _T_2230[5]; // @[Bitwise.scala 50:65:@8209.4]
  assign _T_10239 = _T_2230[6]; // @[Bitwise.scala 50:65:@8210.4]
  assign _T_10240 = _T_2230[7]; // @[Bitwise.scala 50:65:@8211.4]
  assign _T_10241 = _T_2230[8]; // @[Bitwise.scala 50:65:@8212.4]
  assign _T_10242 = _T_2230[9]; // @[Bitwise.scala 50:65:@8213.4]
  assign _T_10243 = _T_2230[10]; // @[Bitwise.scala 50:65:@8214.4]
  assign _T_10244 = _T_2230[11]; // @[Bitwise.scala 50:65:@8215.4]
  assign _T_10245 = _T_2230[12]; // @[Bitwise.scala 50:65:@8216.4]
  assign _T_10246 = _T_2230[13]; // @[Bitwise.scala 50:65:@8217.4]
  assign _T_10247 = _T_2230[14]; // @[Bitwise.scala 50:65:@8218.4]
  assign _T_10248 = _T_2230[15]; // @[Bitwise.scala 50:65:@8219.4]
  assign _T_10249 = _T_2230[16]; // @[Bitwise.scala 50:65:@8220.4]
  assign _T_10250 = _T_2230[17]; // @[Bitwise.scala 50:65:@8221.4]
  assign _T_10251 = _T_2230[18]; // @[Bitwise.scala 50:65:@8222.4]
  assign _T_10252 = _T_2230[19]; // @[Bitwise.scala 50:65:@8223.4]
  assign _T_10253 = _T_2230[20]; // @[Bitwise.scala 50:65:@8224.4]
  assign _T_10254 = _T_2230[21]; // @[Bitwise.scala 50:65:@8225.4]
  assign _T_10255 = _T_2230[22]; // @[Bitwise.scala 50:65:@8226.4]
  assign _T_10256 = _T_2230[23]; // @[Bitwise.scala 50:65:@8227.4]
  assign _T_10257 = _T_2230[24]; // @[Bitwise.scala 50:65:@8228.4]
  assign _T_10258 = _T_2230[25]; // @[Bitwise.scala 50:65:@8229.4]
  assign _T_10259 = _T_2230[26]; // @[Bitwise.scala 50:65:@8230.4]
  assign _T_10260 = _T_2230[27]; // @[Bitwise.scala 50:65:@8231.4]
  assign _T_10261 = _T_2230[28]; // @[Bitwise.scala 50:65:@8232.4]
  assign _T_10262 = _T_2230[29]; // @[Bitwise.scala 50:65:@8233.4]
  assign _T_10263 = _T_2230[30]; // @[Bitwise.scala 50:65:@8234.4]
  assign _T_10264 = _T_2230[31]; // @[Bitwise.scala 50:65:@8235.4]
  assign _T_10265 = _T_2230[32]; // @[Bitwise.scala 50:65:@8236.4]
  assign _T_10266 = _T_2230[33]; // @[Bitwise.scala 50:65:@8237.4]
  assign _T_10267 = _T_2230[34]; // @[Bitwise.scala 50:65:@8238.4]
  assign _T_10268 = _T_2230[35]; // @[Bitwise.scala 50:65:@8239.4]
  assign _T_10269 = _T_2230[36]; // @[Bitwise.scala 50:65:@8240.4]
  assign _T_10270 = _T_2230[37]; // @[Bitwise.scala 50:65:@8241.4]
  assign _T_10271 = _T_2230[38]; // @[Bitwise.scala 50:65:@8242.4]
  assign _T_10272 = _T_2230[39]; // @[Bitwise.scala 50:65:@8243.4]
  assign _T_10273 = _T_2230[40]; // @[Bitwise.scala 50:65:@8244.4]
  assign _T_10274 = _T_2230[41]; // @[Bitwise.scala 50:65:@8245.4]
  assign _T_10275 = _T_2230[42]; // @[Bitwise.scala 50:65:@8246.4]
  assign _T_10276 = _T_2230[43]; // @[Bitwise.scala 50:65:@8247.4]
  assign _T_10277 = _T_2230[44]; // @[Bitwise.scala 50:65:@8248.4]
  assign _T_10278 = _T_2230[45]; // @[Bitwise.scala 50:65:@8249.4]
  assign _T_10279 = _T_2230[46]; // @[Bitwise.scala 50:65:@8250.4]
  assign _T_10280 = _T_2230[47]; // @[Bitwise.scala 50:65:@8251.4]
  assign _T_10281 = _T_2230[48]; // @[Bitwise.scala 50:65:@8252.4]
  assign _T_10282 = _T_2230[49]; // @[Bitwise.scala 50:65:@8253.4]
  assign _T_10283 = _T_2230[50]; // @[Bitwise.scala 50:65:@8254.4]
  assign _T_10284 = _T_2230[51]; // @[Bitwise.scala 50:65:@8255.4]
  assign _T_10285 = _T_2230[52]; // @[Bitwise.scala 50:65:@8256.4]
  assign _T_10286 = _T_2230[53]; // @[Bitwise.scala 50:65:@8257.4]
  assign _T_10287 = _T_2230[54]; // @[Bitwise.scala 50:65:@8258.4]
  assign _T_10288 = _T_2230[55]; // @[Bitwise.scala 50:65:@8259.4]
  assign _T_10289 = _T_2230[56]; // @[Bitwise.scala 50:65:@8260.4]
  assign _T_10290 = _T_2230[57]; // @[Bitwise.scala 50:65:@8261.4]
  assign _T_10291 = _T_2230[58]; // @[Bitwise.scala 50:65:@8262.4]
  assign _T_10292 = _T_2230[59]; // @[Bitwise.scala 50:65:@8263.4]
  assign _T_10293 = _T_2230[60]; // @[Bitwise.scala 50:65:@8264.4]
  assign _T_10294 = _T_2230[61]; // @[Bitwise.scala 50:65:@8265.4]
  assign _T_10295 = _T_2230[62]; // @[Bitwise.scala 50:65:@8266.4]
  assign _T_10296 = _T_2230[63]; // @[Bitwise.scala 50:65:@8267.4]
  assign _T_10297 = _T_2231 + _T_10234; // @[Bitwise.scala 48:55:@8268.4]
  assign _T_10298 = _T_10235 + _T_10236; // @[Bitwise.scala 48:55:@8269.4]
  assign _T_10299 = _T_10297 + _T_10298; // @[Bitwise.scala 48:55:@8270.4]
  assign _T_10300 = _T_10237 + _T_10238; // @[Bitwise.scala 48:55:@8271.4]
  assign _T_10301 = _T_10239 + _T_10240; // @[Bitwise.scala 48:55:@8272.4]
  assign _T_10302 = _T_10300 + _T_10301; // @[Bitwise.scala 48:55:@8273.4]
  assign _T_10303 = _T_10299 + _T_10302; // @[Bitwise.scala 48:55:@8274.4]
  assign _T_10304 = _T_10241 + _T_10242; // @[Bitwise.scala 48:55:@8275.4]
  assign _T_10305 = _T_10243 + _T_10244; // @[Bitwise.scala 48:55:@8276.4]
  assign _T_10306 = _T_10304 + _T_10305; // @[Bitwise.scala 48:55:@8277.4]
  assign _T_10307 = _T_10245 + _T_10246; // @[Bitwise.scala 48:55:@8278.4]
  assign _T_10308 = _T_10247 + _T_10248; // @[Bitwise.scala 48:55:@8279.4]
  assign _T_10309 = _T_10307 + _T_10308; // @[Bitwise.scala 48:55:@8280.4]
  assign _T_10310 = _T_10306 + _T_10309; // @[Bitwise.scala 48:55:@8281.4]
  assign _T_10311 = _T_10303 + _T_10310; // @[Bitwise.scala 48:55:@8282.4]
  assign _T_10312 = _T_10249 + _T_10250; // @[Bitwise.scala 48:55:@8283.4]
  assign _T_10313 = _T_10251 + _T_10252; // @[Bitwise.scala 48:55:@8284.4]
  assign _T_10314 = _T_10312 + _T_10313; // @[Bitwise.scala 48:55:@8285.4]
  assign _T_10315 = _T_10253 + _T_10254; // @[Bitwise.scala 48:55:@8286.4]
  assign _T_10316 = _T_10255 + _T_10256; // @[Bitwise.scala 48:55:@8287.4]
  assign _T_10317 = _T_10315 + _T_10316; // @[Bitwise.scala 48:55:@8288.4]
  assign _T_10318 = _T_10314 + _T_10317; // @[Bitwise.scala 48:55:@8289.4]
  assign _T_10319 = _T_10257 + _T_10258; // @[Bitwise.scala 48:55:@8290.4]
  assign _T_10320 = _T_10259 + _T_10260; // @[Bitwise.scala 48:55:@8291.4]
  assign _T_10321 = _T_10319 + _T_10320; // @[Bitwise.scala 48:55:@8292.4]
  assign _T_10322 = _T_10261 + _T_10262; // @[Bitwise.scala 48:55:@8293.4]
  assign _T_10323 = _T_10263 + _T_10264; // @[Bitwise.scala 48:55:@8294.4]
  assign _T_10324 = _T_10322 + _T_10323; // @[Bitwise.scala 48:55:@8295.4]
  assign _T_10325 = _T_10321 + _T_10324; // @[Bitwise.scala 48:55:@8296.4]
  assign _T_10326 = _T_10318 + _T_10325; // @[Bitwise.scala 48:55:@8297.4]
  assign _T_10327 = _T_10311 + _T_10326; // @[Bitwise.scala 48:55:@8298.4]
  assign _T_10328 = _T_10265 + _T_10266; // @[Bitwise.scala 48:55:@8299.4]
  assign _T_10329 = _T_10267 + _T_10268; // @[Bitwise.scala 48:55:@8300.4]
  assign _T_10330 = _T_10328 + _T_10329; // @[Bitwise.scala 48:55:@8301.4]
  assign _T_10331 = _T_10269 + _T_10270; // @[Bitwise.scala 48:55:@8302.4]
  assign _T_10332 = _T_10271 + _T_10272; // @[Bitwise.scala 48:55:@8303.4]
  assign _T_10333 = _T_10331 + _T_10332; // @[Bitwise.scala 48:55:@8304.4]
  assign _T_10334 = _T_10330 + _T_10333; // @[Bitwise.scala 48:55:@8305.4]
  assign _T_10335 = _T_10273 + _T_10274; // @[Bitwise.scala 48:55:@8306.4]
  assign _T_10336 = _T_10275 + _T_10276; // @[Bitwise.scala 48:55:@8307.4]
  assign _T_10337 = _T_10335 + _T_10336; // @[Bitwise.scala 48:55:@8308.4]
  assign _T_10338 = _T_10277 + _T_10278; // @[Bitwise.scala 48:55:@8309.4]
  assign _T_10339 = _T_10279 + _T_10280; // @[Bitwise.scala 48:55:@8310.4]
  assign _T_10340 = _T_10338 + _T_10339; // @[Bitwise.scala 48:55:@8311.4]
  assign _T_10341 = _T_10337 + _T_10340; // @[Bitwise.scala 48:55:@8312.4]
  assign _T_10342 = _T_10334 + _T_10341; // @[Bitwise.scala 48:55:@8313.4]
  assign _T_10343 = _T_10281 + _T_10282; // @[Bitwise.scala 48:55:@8314.4]
  assign _T_10344 = _T_10283 + _T_10284; // @[Bitwise.scala 48:55:@8315.4]
  assign _T_10345 = _T_10343 + _T_10344; // @[Bitwise.scala 48:55:@8316.4]
  assign _T_10346 = _T_10285 + _T_10286; // @[Bitwise.scala 48:55:@8317.4]
  assign _T_10347 = _T_10287 + _T_10288; // @[Bitwise.scala 48:55:@8318.4]
  assign _T_10348 = _T_10346 + _T_10347; // @[Bitwise.scala 48:55:@8319.4]
  assign _T_10349 = _T_10345 + _T_10348; // @[Bitwise.scala 48:55:@8320.4]
  assign _T_10350 = _T_10289 + _T_10290; // @[Bitwise.scala 48:55:@8321.4]
  assign _T_10351 = _T_10291 + _T_10292; // @[Bitwise.scala 48:55:@8322.4]
  assign _T_10352 = _T_10350 + _T_10351; // @[Bitwise.scala 48:55:@8323.4]
  assign _T_10353 = _T_10293 + _T_10294; // @[Bitwise.scala 48:55:@8324.4]
  assign _T_10354 = _T_10295 + _T_10296; // @[Bitwise.scala 48:55:@8325.4]
  assign _T_10355 = _T_10353 + _T_10354; // @[Bitwise.scala 48:55:@8326.4]
  assign _T_10356 = _T_10352 + _T_10355; // @[Bitwise.scala 48:55:@8327.4]
  assign _T_10357 = _T_10349 + _T_10356; // @[Bitwise.scala 48:55:@8328.4]
  assign _T_10358 = _T_10342 + _T_10357; // @[Bitwise.scala 48:55:@8329.4]
  assign _T_10359 = _T_10327 + _T_10358; // @[Bitwise.scala 48:55:@8330.4]
  assign _GEN_128 = io_input_valid ? io_input_bits_sel_0 : _T_10641_0; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_129 = io_input_valid ? io_input_bits_sel_1 : _T_10641_1; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_130 = io_input_valid ? io_input_bits_sel_2 : _T_10641_2; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_131 = io_input_valid ? io_input_bits_sel_3 : _T_10641_3; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_132 = io_input_valid ? io_input_bits_sel_4 : _T_10641_4; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_133 = io_input_valid ? io_input_bits_sel_5 : _T_10641_5; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_134 = io_input_valid ? io_input_bits_sel_6 : _T_10641_6; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_135 = io_input_valid ? io_input_bits_sel_7 : _T_10641_7; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_136 = io_input_valid ? io_input_bits_sel_8 : _T_10641_8; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_137 = io_input_valid ? io_input_bits_sel_9 : _T_10641_9; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_138 = io_input_valid ? io_input_bits_sel_10 : _T_10641_10; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_139 = io_input_valid ? io_input_bits_sel_11 : _T_10641_11; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_140 = io_input_valid ? io_input_bits_sel_12 : _T_10641_12; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_141 = io_input_valid ? io_input_bits_sel_13 : _T_10641_13; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_142 = io_input_valid ? io_input_bits_sel_14 : _T_10641_14; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_143 = io_input_valid ? io_input_bits_sel_15 : _T_10641_15; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_144 = io_input_valid ? io_input_bits_sel_16 : _T_10641_16; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_145 = io_input_valid ? io_input_bits_sel_17 : _T_10641_17; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_146 = io_input_valid ? io_input_bits_sel_18 : _T_10641_18; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_147 = io_input_valid ? io_input_bits_sel_19 : _T_10641_19; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_148 = io_input_valid ? io_input_bits_sel_20 : _T_10641_20; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_149 = io_input_valid ? io_input_bits_sel_21 : _T_10641_21; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_150 = io_input_valid ? io_input_bits_sel_22 : _T_10641_22; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_151 = io_input_valid ? io_input_bits_sel_23 : _T_10641_23; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_152 = io_input_valid ? io_input_bits_sel_24 : _T_10641_24; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_153 = io_input_valid ? io_input_bits_sel_25 : _T_10641_25; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_154 = io_input_valid ? io_input_bits_sel_26 : _T_10641_26; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_155 = io_input_valid ? io_input_bits_sel_27 : _T_10641_27; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_156 = io_input_valid ? io_input_bits_sel_28 : _T_10641_28; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_157 = io_input_valid ? io_input_bits_sel_29 : _T_10641_29; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_158 = io_input_valid ? io_input_bits_sel_30 : _T_10641_30; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _GEN_159 = io_input_valid ? io_input_bits_sel_31 : _T_10641_31; // @[NV_NVDLA_CSC_WL_dec.scala 71:25:@8499.4]
  assign _T_11318 = io_input_mask_en[0]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8661.4]
  assign _T_11319 = io_input_valid & _T_11318; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8662.4]
  assign _GEN_160 = _T_11319 ? _T_2231 : _T_11317_0; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8663.4]
  assign _GEN_161 = _T_11319 ? _T_2299 : _T_11317_1; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8668.4]
  assign _T_2167_2 = _T_2368[1:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@279.4]
  assign _GEN_162 = _T_11319 ? _T_2167_2 : _T_11317_2; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8673.4]
  assign _GEN_163 = _T_11319 ? _T_2439 : _T_11317_3; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8678.4]
  assign _T_2167_4 = _T_2512[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@425.4]
  assign _GEN_164 = _T_11319 ? _T_2167_4 : _T_11317_4; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8683.4]
  assign _T_2167_5 = _T_2587[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@501.4]
  assign _GEN_165 = _T_11319 ? _T_2167_5 : _T_11317_5; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8688.4]
  assign _T_2167_6 = _T_2664[2:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@579.4]
  assign _GEN_166 = _T_11319 ? _T_2167_6 : _T_11317_6; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8693.4]
  assign _GEN_167 = _T_11319 ? _T_2743 : _T_11317_7; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8698.4]
  assign _T_11334 = io_input_mask_en[1]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8701.4]
  assign _T_11335 = io_input_valid & _T_11334; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8702.4]
  assign _T_2167_8 = _T_2824[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@741.4]
  assign _GEN_168 = _T_11335 ? _T_2167_8 : _T_11317_8; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8703.4]
  assign _T_2167_9 = _T_2907[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@825.4]
  assign _GEN_169 = _T_11335 ? _T_2167_9 : _T_11317_9; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8708.4]
  assign _T_2167_10 = _T_2992[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@911.4]
  assign _GEN_170 = _T_11335 ? _T_2167_10 : _T_11317_10; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8713.4]
  assign _T_2167_11 = _T_3079[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@999.4]
  assign _GEN_171 = _T_11335 ? _T_2167_11 : _T_11317_11; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8718.4]
  assign _T_2167_12 = _T_3168[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1089.4]
  assign _GEN_172 = _T_11335 ? _T_2167_12 : _T_11317_12; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8723.4]
  assign _T_2167_13 = _T_3259[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1181.4]
  assign _GEN_173 = _T_11335 ? _T_2167_13 : _T_11317_13; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8728.4]
  assign _T_2167_14 = _T_3352[3:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1275.4]
  assign _GEN_174 = _T_11335 ? _T_2167_14 : _T_11317_14; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8733.4]
  assign _GEN_175 = _T_11335 ? _T_3447 : _T_11317_15; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8738.4]
  assign _T_11350 = io_input_mask_en[2]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8741.4]
  assign _T_11351 = io_input_valid & _T_11350; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8742.4]
  assign _T_2167_16 = _T_3544[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1469.4]
  assign _GEN_176 = _T_11351 ? _T_2167_16 : _T_11317_16; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8743.4]
  assign _T_2167_17 = _T_3643[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1569.4]
  assign _GEN_177 = _T_11351 ? _T_2167_17 : _T_11317_17; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8748.4]
  assign _T_2167_18 = _T_3744[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1671.4]
  assign _GEN_178 = _T_11351 ? _T_2167_18 : _T_11317_18; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8753.4]
  assign _T_2167_19 = _T_3847[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1775.4]
  assign _GEN_179 = _T_11351 ? _T_2167_19 : _T_11317_19; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8758.4]
  assign _T_2167_20 = _T_3952[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1881.4]
  assign _GEN_180 = _T_11351 ? _T_2167_20 : _T_11317_20; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8763.4]
  assign _T_2167_21 = _T_4059[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@1989.4]
  assign _GEN_181 = _T_11351 ? _T_2167_21 : _T_11317_21; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8768.4]
  assign _T_2167_22 = _T_4168[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2099.4]
  assign _GEN_182 = _T_11351 ? _T_2167_22 : _T_11317_22; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8773.4]
  assign _T_2167_23 = _T_4279[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2211.4]
  assign _GEN_183 = _T_11351 ? _T_2167_23 : _T_11317_23; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8778.4]
  assign _T_11366 = io_input_mask_en[3]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8781.4]
  assign _T_11367 = io_input_valid & _T_11366; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8782.4]
  assign _T_2167_24 = _T_4392[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2325.4]
  assign _GEN_184 = _T_11367 ? _T_2167_24 : _T_11317_24; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8783.4]
  assign _T_2167_25 = _T_4507[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2441.4]
  assign _GEN_185 = _T_11367 ? _T_2167_25 : _T_11317_25; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8788.4]
  assign _T_2167_26 = _T_4624[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2559.4]
  assign _GEN_186 = _T_11367 ? _T_2167_26 : _T_11317_26; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8793.4]
  assign _T_2167_27 = _T_4743[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2679.4]
  assign _GEN_187 = _T_11367 ? _T_2167_27 : _T_11317_27; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8798.4]
  assign _T_2167_28 = _T_4864[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2801.4]
  assign _GEN_188 = _T_11367 ? _T_2167_28 : _T_11317_28; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8803.4]
  assign _T_2167_29 = _T_4987[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@2925.4]
  assign _GEN_189 = _T_11367 ? _T_2167_29 : _T_11317_29; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8808.4]
  assign _T_2167_30 = _T_5112[4:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3051.4]
  assign _GEN_190 = _T_11367 ? _T_2167_30 : _T_11317_30; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8813.4]
  assign _GEN_191 = _T_11367 ? _T_5239 : _T_11317_31; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8818.4]
  assign _T_11382 = io_input_mask_en[4]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8821.4]
  assign _T_11383 = io_input_valid & _T_11382; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8822.4]
  assign _T_2167_32 = _T_5368[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3309.4]
  assign _GEN_192 = _T_11383 ? _T_2167_32 : _T_11317_32; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8823.4]
  assign _T_2167_33 = _T_5499[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3441.4]
  assign _GEN_193 = _T_11383 ? _T_2167_33 : _T_11317_33; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8828.4]
  assign _T_2167_34 = _T_5632[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3575.4]
  assign _GEN_194 = _T_11383 ? _T_2167_34 : _T_11317_34; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8833.4]
  assign _T_2167_35 = _T_5767[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3711.4]
  assign _GEN_195 = _T_11383 ? _T_2167_35 : _T_11317_35; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8838.4]
  assign _T_2167_36 = _T_5904[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3849.4]
  assign _GEN_196 = _T_11383 ? _T_2167_36 : _T_11317_36; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8843.4]
  assign _T_2167_37 = _T_6043[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@3989.4]
  assign _GEN_197 = _T_11383 ? _T_2167_37 : _T_11317_37; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8848.4]
  assign _T_2167_38 = _T_6184[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4131.4]
  assign _GEN_198 = _T_11383 ? _T_2167_38 : _T_11317_38; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8853.4]
  assign _T_2167_39 = _T_6327[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4275.4]
  assign _GEN_199 = _T_11383 ? _T_2167_39 : _T_11317_39; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8858.4]
  assign _T_11398 = io_input_mask_en[5]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8861.4]
  assign _T_11399 = io_input_valid & _T_11398; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8862.4]
  assign _T_2167_40 = _T_6472[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4421.4]
  assign _GEN_200 = _T_11399 ? _T_2167_40 : _T_11317_40; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8863.4]
  assign _T_2167_41 = _T_6619[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4569.4]
  assign _GEN_201 = _T_11399 ? _T_2167_41 : _T_11317_41; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8868.4]
  assign _T_2167_42 = _T_6768[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4719.4]
  assign _GEN_202 = _T_11399 ? _T_2167_42 : _T_11317_42; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8873.4]
  assign _T_2167_43 = _T_6919[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@4871.4]
  assign _GEN_203 = _T_11399 ? _T_2167_43 : _T_11317_43; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8878.4]
  assign _T_2167_44 = _T_7072[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5025.4]
  assign _GEN_204 = _T_11399 ? _T_2167_44 : _T_11317_44; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8883.4]
  assign _T_2167_45 = _T_7227[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5181.4]
  assign _GEN_205 = _T_11399 ? _T_2167_45 : _T_11317_45; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8888.4]
  assign _T_2167_46 = _T_7384[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5339.4]
  assign _GEN_206 = _T_11399 ? _T_2167_46 : _T_11317_46; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8893.4]
  assign _T_2167_47 = _T_7543[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5499.4]
  assign _GEN_207 = _T_11399 ? _T_2167_47 : _T_11317_47; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8898.4]
  assign _T_11414 = io_input_mask_en[6]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8901.4]
  assign _T_11415 = io_input_valid & _T_11414; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8902.4]
  assign _T_2167_48 = _T_7704[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5661.4]
  assign _GEN_208 = _T_11415 ? _T_2167_48 : _T_11317_48; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8903.4]
  assign _T_2167_49 = _T_7867[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5825.4]
  assign _GEN_209 = _T_11415 ? _T_2167_49 : _T_11317_49; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8908.4]
  assign _T_2167_50 = _T_8032[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@5991.4]
  assign _GEN_210 = _T_11415 ? _T_2167_50 : _T_11317_50; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8913.4]
  assign _T_2167_51 = _T_8199[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6159.4]
  assign _GEN_211 = _T_11415 ? _T_2167_51 : _T_11317_51; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8918.4]
  assign _T_2167_52 = _T_8368[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6329.4]
  assign _GEN_212 = _T_11415 ? _T_2167_52 : _T_11317_52; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8923.4]
  assign _T_2167_53 = _T_8539[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6501.4]
  assign _GEN_213 = _T_11415 ? _T_2167_53 : _T_11317_53; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8928.4]
  assign _T_2167_54 = _T_8712[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6675.4]
  assign _GEN_214 = _T_11415 ? _T_2167_54 : _T_11317_54; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8933.4]
  assign _T_2167_55 = _T_8887[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@6851.4]
  assign _GEN_215 = _T_11415 ? _T_2167_55 : _T_11317_55; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8938.4]
  assign _T_11430 = io_input_mask_en[7]; // @[NV_NVDLA_CSC_WL_dec.scala 78:47:@8941.4]
  assign _T_11431 = io_input_valid & _T_11430; // @[NV_NVDLA_CSC_WL_dec.scala 78:29:@8942.4]
  assign _T_2167_56 = _T_9064[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7029.4]
  assign _GEN_216 = _T_11431 ? _T_2167_56 : _T_11317_56; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8943.4]
  assign _T_2167_57 = _T_9243[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7209.4]
  assign _GEN_217 = _T_11431 ? _T_2167_57 : _T_11317_57; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8948.4]
  assign _T_2167_58 = _T_9424[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7391.4]
  assign _GEN_218 = _T_11431 ? _T_2167_58 : _T_11317_58; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8953.4]
  assign _T_2167_59 = _T_9607[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7575.4]
  assign _GEN_219 = _T_11431 ? _T_2167_59 : _T_11317_59; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8958.4]
  assign _T_2167_60 = _T_9792[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7761.4]
  assign _GEN_220 = _T_11431 ? _T_2167_60 : _T_11317_60; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8963.4]
  assign _T_2167_61 = _T_9979[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@7949.4]
  assign _GEN_221 = _T_11431 ? _T_2167_61 : _T_11317_61; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8968.4]
  assign _T_2167_62 = _T_10168[5:0]; // @[NV_NVDLA_CSC_WL_dec.scala 57:23:@75.4 NV_NVDLA_CSC_WL_dec.scala 60:20:@8139.4]
  assign _GEN_222 = _T_11431 ? _T_2167_62 : _T_11317_62; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8973.4]
  assign _GEN_223 = _T_11431 ? _T_10359 : _T_11317_63; // @[NV_NVDLA_CSC_WL_dec.scala 79:9:@8978.4]
  assign _T_11519 = _T_11317_0 ? _T_10366_0 : 8'h0; // @[Mux.scala 46:16:@8983.4]
  assign _T_11523 = 2'h2 == _T_11317_1; // @[Mux.scala 46:19:@8985.4]
  assign _T_11524 = _T_11523 ? _T_10366_1 : 8'h0; // @[Mux.scala 46:16:@8986.4]
  assign _T_11525 = 2'h1 == _T_11317_1; // @[Mux.scala 46:19:@8987.4]
  assign _T_11526 = _T_11525 ? _T_10366_0 : _T_11524; // @[Mux.scala 46:16:@8988.4]
  assign _T_11531 = 2'h3 == _T_11317_2; // @[Mux.scala 46:19:@8990.4]
  assign _T_11532 = _T_11531 ? _T_10366_2 : 8'h0; // @[Mux.scala 46:16:@8991.4]
  assign _T_11533 = 2'h2 == _T_11317_2; // @[Mux.scala 46:19:@8992.4]
  assign _T_11534 = _T_11533 ? _T_10366_1 : _T_11532; // @[Mux.scala 46:16:@8993.4]
  assign _T_11535 = 2'h1 == _T_11317_2; // @[Mux.scala 46:19:@8994.4]
  assign _T_11536 = _T_11535 ? _T_10366_0 : _T_11534; // @[Mux.scala 46:16:@8995.4]
  assign _T_11542 = 3'h4 == _T_11317_3; // @[Mux.scala 46:19:@8997.4]
  assign _T_11543 = _T_11542 ? _T_10366_3 : 8'h0; // @[Mux.scala 46:16:@8998.4]
  assign _T_11544 = 3'h3 == _T_11317_3; // @[Mux.scala 46:19:@8999.4]
  assign _T_11545 = _T_11544 ? _T_10366_2 : _T_11543; // @[Mux.scala 46:16:@9000.4]
  assign _T_11546 = 3'h2 == _T_11317_3; // @[Mux.scala 46:19:@9001.4]
  assign _T_11547 = _T_11546 ? _T_10366_1 : _T_11545; // @[Mux.scala 46:16:@9002.4]
  assign _T_11548 = 3'h1 == _T_11317_3; // @[Mux.scala 46:19:@9003.4]
  assign _T_11549 = _T_11548 ? _T_10366_0 : _T_11547; // @[Mux.scala 46:16:@9004.4]
  assign _T_11556 = 3'h5 == _T_11317_4; // @[Mux.scala 46:19:@9006.4]
  assign _T_11557 = _T_11556 ? _T_10366_4 : 8'h0; // @[Mux.scala 46:16:@9007.4]
  assign _T_11558 = 3'h4 == _T_11317_4; // @[Mux.scala 46:19:@9008.4]
  assign _T_11559 = _T_11558 ? _T_10366_3 : _T_11557; // @[Mux.scala 46:16:@9009.4]
  assign _T_11560 = 3'h3 == _T_11317_4; // @[Mux.scala 46:19:@9010.4]
  assign _T_11561 = _T_11560 ? _T_10366_2 : _T_11559; // @[Mux.scala 46:16:@9011.4]
  assign _T_11562 = 3'h2 == _T_11317_4; // @[Mux.scala 46:19:@9012.4]
  assign _T_11563 = _T_11562 ? _T_10366_1 : _T_11561; // @[Mux.scala 46:16:@9013.4]
  assign _T_11564 = 3'h1 == _T_11317_4; // @[Mux.scala 46:19:@9014.4]
  assign _T_11565 = _T_11564 ? _T_10366_0 : _T_11563; // @[Mux.scala 46:16:@9015.4]
  assign _T_11573 = 3'h6 == _T_11317_5; // @[Mux.scala 46:19:@9017.4]
  assign _T_11574 = _T_11573 ? _T_10366_5 : 8'h0; // @[Mux.scala 46:16:@9018.4]
  assign _T_11575 = 3'h5 == _T_11317_5; // @[Mux.scala 46:19:@9019.4]
  assign _T_11576 = _T_11575 ? _T_10366_4 : _T_11574; // @[Mux.scala 46:16:@9020.4]
  assign _T_11577 = 3'h4 == _T_11317_5; // @[Mux.scala 46:19:@9021.4]
  assign _T_11578 = _T_11577 ? _T_10366_3 : _T_11576; // @[Mux.scala 46:16:@9022.4]
  assign _T_11579 = 3'h3 == _T_11317_5; // @[Mux.scala 46:19:@9023.4]
  assign _T_11580 = _T_11579 ? _T_10366_2 : _T_11578; // @[Mux.scala 46:16:@9024.4]
  assign _T_11581 = 3'h2 == _T_11317_5; // @[Mux.scala 46:19:@9025.4]
  assign _T_11582 = _T_11581 ? _T_10366_1 : _T_11580; // @[Mux.scala 46:16:@9026.4]
  assign _T_11583 = 3'h1 == _T_11317_5; // @[Mux.scala 46:19:@9027.4]
  assign _T_11584 = _T_11583 ? _T_10366_0 : _T_11582; // @[Mux.scala 46:16:@9028.4]
  assign _T_11593 = 3'h7 == _T_11317_6; // @[Mux.scala 46:19:@9030.4]
  assign _T_11594 = _T_11593 ? _T_10366_6 : 8'h0; // @[Mux.scala 46:16:@9031.4]
  assign _T_11595 = 3'h6 == _T_11317_6; // @[Mux.scala 46:19:@9032.4]
  assign _T_11596 = _T_11595 ? _T_10366_5 : _T_11594; // @[Mux.scala 46:16:@9033.4]
  assign _T_11597 = 3'h5 == _T_11317_6; // @[Mux.scala 46:19:@9034.4]
  assign _T_11598 = _T_11597 ? _T_10366_4 : _T_11596; // @[Mux.scala 46:16:@9035.4]
  assign _T_11599 = 3'h4 == _T_11317_6; // @[Mux.scala 46:19:@9036.4]
  assign _T_11600 = _T_11599 ? _T_10366_3 : _T_11598; // @[Mux.scala 46:16:@9037.4]
  assign _T_11601 = 3'h3 == _T_11317_6; // @[Mux.scala 46:19:@9038.4]
  assign _T_11602 = _T_11601 ? _T_10366_2 : _T_11600; // @[Mux.scala 46:16:@9039.4]
  assign _T_11603 = 3'h2 == _T_11317_6; // @[Mux.scala 46:19:@9040.4]
  assign _T_11604 = _T_11603 ? _T_10366_1 : _T_11602; // @[Mux.scala 46:16:@9041.4]
  assign _T_11605 = 3'h1 == _T_11317_6; // @[Mux.scala 46:19:@9042.4]
  assign _T_11606 = _T_11605 ? _T_10366_0 : _T_11604; // @[Mux.scala 46:16:@9043.4]
  assign _T_11616 = 4'h8 == _T_11317_7; // @[Mux.scala 46:19:@9045.4]
  assign _T_11617 = _T_11616 ? _T_10366_7 : 8'h0; // @[Mux.scala 46:16:@9046.4]
  assign _T_11618 = 4'h7 == _T_11317_7; // @[Mux.scala 46:19:@9047.4]
  assign _T_11619 = _T_11618 ? _T_10366_6 : _T_11617; // @[Mux.scala 46:16:@9048.4]
  assign _T_11620 = 4'h6 == _T_11317_7; // @[Mux.scala 46:19:@9049.4]
  assign _T_11621 = _T_11620 ? _T_10366_5 : _T_11619; // @[Mux.scala 46:16:@9050.4]
  assign _T_11622 = 4'h5 == _T_11317_7; // @[Mux.scala 46:19:@9051.4]
  assign _T_11623 = _T_11622 ? _T_10366_4 : _T_11621; // @[Mux.scala 46:16:@9052.4]
  assign _T_11624 = 4'h4 == _T_11317_7; // @[Mux.scala 46:19:@9053.4]
  assign _T_11625 = _T_11624 ? _T_10366_3 : _T_11623; // @[Mux.scala 46:16:@9054.4]
  assign _T_11626 = 4'h3 == _T_11317_7; // @[Mux.scala 46:19:@9055.4]
  assign _T_11627 = _T_11626 ? _T_10366_2 : _T_11625; // @[Mux.scala 46:16:@9056.4]
  assign _T_11628 = 4'h2 == _T_11317_7; // @[Mux.scala 46:19:@9057.4]
  assign _T_11629 = _T_11628 ? _T_10366_1 : _T_11627; // @[Mux.scala 46:16:@9058.4]
  assign _T_11630 = 4'h1 == _T_11317_7; // @[Mux.scala 46:19:@9059.4]
  assign _T_11631 = _T_11630 ? _T_10366_0 : _T_11629; // @[Mux.scala 46:16:@9060.4]
  assign _T_11642 = 4'h9 == _T_11317_8; // @[Mux.scala 46:19:@9062.4]
  assign _T_11643 = _T_11642 ? _T_10366_8 : 8'h0; // @[Mux.scala 46:16:@9063.4]
  assign _T_11644 = 4'h8 == _T_11317_8; // @[Mux.scala 46:19:@9064.4]
  assign _T_11645 = _T_11644 ? _T_10366_7 : _T_11643; // @[Mux.scala 46:16:@9065.4]
  assign _T_11646 = 4'h7 == _T_11317_8; // @[Mux.scala 46:19:@9066.4]
  assign _T_11647 = _T_11646 ? _T_10366_6 : _T_11645; // @[Mux.scala 46:16:@9067.4]
  assign _T_11648 = 4'h6 == _T_11317_8; // @[Mux.scala 46:19:@9068.4]
  assign _T_11649 = _T_11648 ? _T_10366_5 : _T_11647; // @[Mux.scala 46:16:@9069.4]
  assign _T_11650 = 4'h5 == _T_11317_8; // @[Mux.scala 46:19:@9070.4]
  assign _T_11651 = _T_11650 ? _T_10366_4 : _T_11649; // @[Mux.scala 46:16:@9071.4]
  assign _T_11652 = 4'h4 == _T_11317_8; // @[Mux.scala 46:19:@9072.4]
  assign _T_11653 = _T_11652 ? _T_10366_3 : _T_11651; // @[Mux.scala 46:16:@9073.4]
  assign _T_11654 = 4'h3 == _T_11317_8; // @[Mux.scala 46:19:@9074.4]
  assign _T_11655 = _T_11654 ? _T_10366_2 : _T_11653; // @[Mux.scala 46:16:@9075.4]
  assign _T_11656 = 4'h2 == _T_11317_8; // @[Mux.scala 46:19:@9076.4]
  assign _T_11657 = _T_11656 ? _T_10366_1 : _T_11655; // @[Mux.scala 46:16:@9077.4]
  assign _T_11658 = 4'h1 == _T_11317_8; // @[Mux.scala 46:19:@9078.4]
  assign _T_11659 = _T_11658 ? _T_10366_0 : _T_11657; // @[Mux.scala 46:16:@9079.4]
  assign _T_11671 = 4'ha == _T_11317_9; // @[Mux.scala 46:19:@9081.4]
  assign _T_11672 = _T_11671 ? _T_10366_9 : 8'h0; // @[Mux.scala 46:16:@9082.4]
  assign _T_11673 = 4'h9 == _T_11317_9; // @[Mux.scala 46:19:@9083.4]
  assign _T_11674 = _T_11673 ? _T_10366_8 : _T_11672; // @[Mux.scala 46:16:@9084.4]
  assign _T_11675 = 4'h8 == _T_11317_9; // @[Mux.scala 46:19:@9085.4]
  assign _T_11676 = _T_11675 ? _T_10366_7 : _T_11674; // @[Mux.scala 46:16:@9086.4]
  assign _T_11677 = 4'h7 == _T_11317_9; // @[Mux.scala 46:19:@9087.4]
  assign _T_11678 = _T_11677 ? _T_10366_6 : _T_11676; // @[Mux.scala 46:16:@9088.4]
  assign _T_11679 = 4'h6 == _T_11317_9; // @[Mux.scala 46:19:@9089.4]
  assign _T_11680 = _T_11679 ? _T_10366_5 : _T_11678; // @[Mux.scala 46:16:@9090.4]
  assign _T_11681 = 4'h5 == _T_11317_9; // @[Mux.scala 46:19:@9091.4]
  assign _T_11682 = _T_11681 ? _T_10366_4 : _T_11680; // @[Mux.scala 46:16:@9092.4]
  assign _T_11683 = 4'h4 == _T_11317_9; // @[Mux.scala 46:19:@9093.4]
  assign _T_11684 = _T_11683 ? _T_10366_3 : _T_11682; // @[Mux.scala 46:16:@9094.4]
  assign _T_11685 = 4'h3 == _T_11317_9; // @[Mux.scala 46:19:@9095.4]
  assign _T_11686 = _T_11685 ? _T_10366_2 : _T_11684; // @[Mux.scala 46:16:@9096.4]
  assign _T_11687 = 4'h2 == _T_11317_9; // @[Mux.scala 46:19:@9097.4]
  assign _T_11688 = _T_11687 ? _T_10366_1 : _T_11686; // @[Mux.scala 46:16:@9098.4]
  assign _T_11689 = 4'h1 == _T_11317_9; // @[Mux.scala 46:19:@9099.4]
  assign _T_11690 = _T_11689 ? _T_10366_0 : _T_11688; // @[Mux.scala 46:16:@9100.4]
  assign _T_11703 = 4'hb == _T_11317_10; // @[Mux.scala 46:19:@9102.4]
  assign _T_11704 = _T_11703 ? _T_10366_10 : 8'h0; // @[Mux.scala 46:16:@9103.4]
  assign _T_11705 = 4'ha == _T_11317_10; // @[Mux.scala 46:19:@9104.4]
  assign _T_11706 = _T_11705 ? _T_10366_9 : _T_11704; // @[Mux.scala 46:16:@9105.4]
  assign _T_11707 = 4'h9 == _T_11317_10; // @[Mux.scala 46:19:@9106.4]
  assign _T_11708 = _T_11707 ? _T_10366_8 : _T_11706; // @[Mux.scala 46:16:@9107.4]
  assign _T_11709 = 4'h8 == _T_11317_10; // @[Mux.scala 46:19:@9108.4]
  assign _T_11710 = _T_11709 ? _T_10366_7 : _T_11708; // @[Mux.scala 46:16:@9109.4]
  assign _T_11711 = 4'h7 == _T_11317_10; // @[Mux.scala 46:19:@9110.4]
  assign _T_11712 = _T_11711 ? _T_10366_6 : _T_11710; // @[Mux.scala 46:16:@9111.4]
  assign _T_11713 = 4'h6 == _T_11317_10; // @[Mux.scala 46:19:@9112.4]
  assign _T_11714 = _T_11713 ? _T_10366_5 : _T_11712; // @[Mux.scala 46:16:@9113.4]
  assign _T_11715 = 4'h5 == _T_11317_10; // @[Mux.scala 46:19:@9114.4]
  assign _T_11716 = _T_11715 ? _T_10366_4 : _T_11714; // @[Mux.scala 46:16:@9115.4]
  assign _T_11717 = 4'h4 == _T_11317_10; // @[Mux.scala 46:19:@9116.4]
  assign _T_11718 = _T_11717 ? _T_10366_3 : _T_11716; // @[Mux.scala 46:16:@9117.4]
  assign _T_11719 = 4'h3 == _T_11317_10; // @[Mux.scala 46:19:@9118.4]
  assign _T_11720 = _T_11719 ? _T_10366_2 : _T_11718; // @[Mux.scala 46:16:@9119.4]
  assign _T_11721 = 4'h2 == _T_11317_10; // @[Mux.scala 46:19:@9120.4]
  assign _T_11722 = _T_11721 ? _T_10366_1 : _T_11720; // @[Mux.scala 46:16:@9121.4]
  assign _T_11723 = 4'h1 == _T_11317_10; // @[Mux.scala 46:19:@9122.4]
  assign _T_11724 = _T_11723 ? _T_10366_0 : _T_11722; // @[Mux.scala 46:16:@9123.4]
  assign _T_11738 = 4'hc == _T_11317_11; // @[Mux.scala 46:19:@9125.4]
  assign _T_11739 = _T_11738 ? _T_10366_11 : 8'h0; // @[Mux.scala 46:16:@9126.4]
  assign _T_11740 = 4'hb == _T_11317_11; // @[Mux.scala 46:19:@9127.4]
  assign _T_11741 = _T_11740 ? _T_10366_10 : _T_11739; // @[Mux.scala 46:16:@9128.4]
  assign _T_11742 = 4'ha == _T_11317_11; // @[Mux.scala 46:19:@9129.4]
  assign _T_11743 = _T_11742 ? _T_10366_9 : _T_11741; // @[Mux.scala 46:16:@9130.4]
  assign _T_11744 = 4'h9 == _T_11317_11; // @[Mux.scala 46:19:@9131.4]
  assign _T_11745 = _T_11744 ? _T_10366_8 : _T_11743; // @[Mux.scala 46:16:@9132.4]
  assign _T_11746 = 4'h8 == _T_11317_11; // @[Mux.scala 46:19:@9133.4]
  assign _T_11747 = _T_11746 ? _T_10366_7 : _T_11745; // @[Mux.scala 46:16:@9134.4]
  assign _T_11748 = 4'h7 == _T_11317_11; // @[Mux.scala 46:19:@9135.4]
  assign _T_11749 = _T_11748 ? _T_10366_6 : _T_11747; // @[Mux.scala 46:16:@9136.4]
  assign _T_11750 = 4'h6 == _T_11317_11; // @[Mux.scala 46:19:@9137.4]
  assign _T_11751 = _T_11750 ? _T_10366_5 : _T_11749; // @[Mux.scala 46:16:@9138.4]
  assign _T_11752 = 4'h5 == _T_11317_11; // @[Mux.scala 46:19:@9139.4]
  assign _T_11753 = _T_11752 ? _T_10366_4 : _T_11751; // @[Mux.scala 46:16:@9140.4]
  assign _T_11754 = 4'h4 == _T_11317_11; // @[Mux.scala 46:19:@9141.4]
  assign _T_11755 = _T_11754 ? _T_10366_3 : _T_11753; // @[Mux.scala 46:16:@9142.4]
  assign _T_11756 = 4'h3 == _T_11317_11; // @[Mux.scala 46:19:@9143.4]
  assign _T_11757 = _T_11756 ? _T_10366_2 : _T_11755; // @[Mux.scala 46:16:@9144.4]
  assign _T_11758 = 4'h2 == _T_11317_11; // @[Mux.scala 46:19:@9145.4]
  assign _T_11759 = _T_11758 ? _T_10366_1 : _T_11757; // @[Mux.scala 46:16:@9146.4]
  assign _T_11760 = 4'h1 == _T_11317_11; // @[Mux.scala 46:19:@9147.4]
  assign _T_11761 = _T_11760 ? _T_10366_0 : _T_11759; // @[Mux.scala 46:16:@9148.4]
  assign _T_11776 = 4'hd == _T_11317_12; // @[Mux.scala 46:19:@9150.4]
  assign _T_11777 = _T_11776 ? _T_10366_12 : 8'h0; // @[Mux.scala 46:16:@9151.4]
  assign _T_11778 = 4'hc == _T_11317_12; // @[Mux.scala 46:19:@9152.4]
  assign _T_11779 = _T_11778 ? _T_10366_11 : _T_11777; // @[Mux.scala 46:16:@9153.4]
  assign _T_11780 = 4'hb == _T_11317_12; // @[Mux.scala 46:19:@9154.4]
  assign _T_11781 = _T_11780 ? _T_10366_10 : _T_11779; // @[Mux.scala 46:16:@9155.4]
  assign _T_11782 = 4'ha == _T_11317_12; // @[Mux.scala 46:19:@9156.4]
  assign _T_11783 = _T_11782 ? _T_10366_9 : _T_11781; // @[Mux.scala 46:16:@9157.4]
  assign _T_11784 = 4'h9 == _T_11317_12; // @[Mux.scala 46:19:@9158.4]
  assign _T_11785 = _T_11784 ? _T_10366_8 : _T_11783; // @[Mux.scala 46:16:@9159.4]
  assign _T_11786 = 4'h8 == _T_11317_12; // @[Mux.scala 46:19:@9160.4]
  assign _T_11787 = _T_11786 ? _T_10366_7 : _T_11785; // @[Mux.scala 46:16:@9161.4]
  assign _T_11788 = 4'h7 == _T_11317_12; // @[Mux.scala 46:19:@9162.4]
  assign _T_11789 = _T_11788 ? _T_10366_6 : _T_11787; // @[Mux.scala 46:16:@9163.4]
  assign _T_11790 = 4'h6 == _T_11317_12; // @[Mux.scala 46:19:@9164.4]
  assign _T_11791 = _T_11790 ? _T_10366_5 : _T_11789; // @[Mux.scala 46:16:@9165.4]
  assign _T_11792 = 4'h5 == _T_11317_12; // @[Mux.scala 46:19:@9166.4]
  assign _T_11793 = _T_11792 ? _T_10366_4 : _T_11791; // @[Mux.scala 46:16:@9167.4]
  assign _T_11794 = 4'h4 == _T_11317_12; // @[Mux.scala 46:19:@9168.4]
  assign _T_11795 = _T_11794 ? _T_10366_3 : _T_11793; // @[Mux.scala 46:16:@9169.4]
  assign _T_11796 = 4'h3 == _T_11317_12; // @[Mux.scala 46:19:@9170.4]
  assign _T_11797 = _T_11796 ? _T_10366_2 : _T_11795; // @[Mux.scala 46:16:@9171.4]
  assign _T_11798 = 4'h2 == _T_11317_12; // @[Mux.scala 46:19:@9172.4]
  assign _T_11799 = _T_11798 ? _T_10366_1 : _T_11797; // @[Mux.scala 46:16:@9173.4]
  assign _T_11800 = 4'h1 == _T_11317_12; // @[Mux.scala 46:19:@9174.4]
  assign _T_11801 = _T_11800 ? _T_10366_0 : _T_11799; // @[Mux.scala 46:16:@9175.4]
  assign _T_11817 = 4'he == _T_11317_13; // @[Mux.scala 46:19:@9177.4]
  assign _T_11818 = _T_11817 ? _T_10366_13 : 8'h0; // @[Mux.scala 46:16:@9178.4]
  assign _T_11819 = 4'hd == _T_11317_13; // @[Mux.scala 46:19:@9179.4]
  assign _T_11820 = _T_11819 ? _T_10366_12 : _T_11818; // @[Mux.scala 46:16:@9180.4]
  assign _T_11821 = 4'hc == _T_11317_13; // @[Mux.scala 46:19:@9181.4]
  assign _T_11822 = _T_11821 ? _T_10366_11 : _T_11820; // @[Mux.scala 46:16:@9182.4]
  assign _T_11823 = 4'hb == _T_11317_13; // @[Mux.scala 46:19:@9183.4]
  assign _T_11824 = _T_11823 ? _T_10366_10 : _T_11822; // @[Mux.scala 46:16:@9184.4]
  assign _T_11825 = 4'ha == _T_11317_13; // @[Mux.scala 46:19:@9185.4]
  assign _T_11826 = _T_11825 ? _T_10366_9 : _T_11824; // @[Mux.scala 46:16:@9186.4]
  assign _T_11827 = 4'h9 == _T_11317_13; // @[Mux.scala 46:19:@9187.4]
  assign _T_11828 = _T_11827 ? _T_10366_8 : _T_11826; // @[Mux.scala 46:16:@9188.4]
  assign _T_11829 = 4'h8 == _T_11317_13; // @[Mux.scala 46:19:@9189.4]
  assign _T_11830 = _T_11829 ? _T_10366_7 : _T_11828; // @[Mux.scala 46:16:@9190.4]
  assign _T_11831 = 4'h7 == _T_11317_13; // @[Mux.scala 46:19:@9191.4]
  assign _T_11832 = _T_11831 ? _T_10366_6 : _T_11830; // @[Mux.scala 46:16:@9192.4]
  assign _T_11833 = 4'h6 == _T_11317_13; // @[Mux.scala 46:19:@9193.4]
  assign _T_11834 = _T_11833 ? _T_10366_5 : _T_11832; // @[Mux.scala 46:16:@9194.4]
  assign _T_11835 = 4'h5 == _T_11317_13; // @[Mux.scala 46:19:@9195.4]
  assign _T_11836 = _T_11835 ? _T_10366_4 : _T_11834; // @[Mux.scala 46:16:@9196.4]
  assign _T_11837 = 4'h4 == _T_11317_13; // @[Mux.scala 46:19:@9197.4]
  assign _T_11838 = _T_11837 ? _T_10366_3 : _T_11836; // @[Mux.scala 46:16:@9198.4]
  assign _T_11839 = 4'h3 == _T_11317_13; // @[Mux.scala 46:19:@9199.4]
  assign _T_11840 = _T_11839 ? _T_10366_2 : _T_11838; // @[Mux.scala 46:16:@9200.4]
  assign _T_11841 = 4'h2 == _T_11317_13; // @[Mux.scala 46:19:@9201.4]
  assign _T_11842 = _T_11841 ? _T_10366_1 : _T_11840; // @[Mux.scala 46:16:@9202.4]
  assign _T_11843 = 4'h1 == _T_11317_13; // @[Mux.scala 46:19:@9203.4]
  assign _T_11844 = _T_11843 ? _T_10366_0 : _T_11842; // @[Mux.scala 46:16:@9204.4]
  assign _T_11861 = 4'hf == _T_11317_14; // @[Mux.scala 46:19:@9206.4]
  assign _T_11862 = _T_11861 ? _T_10366_14 : 8'h0; // @[Mux.scala 46:16:@9207.4]
  assign _T_11863 = 4'he == _T_11317_14; // @[Mux.scala 46:19:@9208.4]
  assign _T_11864 = _T_11863 ? _T_10366_13 : _T_11862; // @[Mux.scala 46:16:@9209.4]
  assign _T_11865 = 4'hd == _T_11317_14; // @[Mux.scala 46:19:@9210.4]
  assign _T_11866 = _T_11865 ? _T_10366_12 : _T_11864; // @[Mux.scala 46:16:@9211.4]
  assign _T_11867 = 4'hc == _T_11317_14; // @[Mux.scala 46:19:@9212.4]
  assign _T_11868 = _T_11867 ? _T_10366_11 : _T_11866; // @[Mux.scala 46:16:@9213.4]
  assign _T_11869 = 4'hb == _T_11317_14; // @[Mux.scala 46:19:@9214.4]
  assign _T_11870 = _T_11869 ? _T_10366_10 : _T_11868; // @[Mux.scala 46:16:@9215.4]
  assign _T_11871 = 4'ha == _T_11317_14; // @[Mux.scala 46:19:@9216.4]
  assign _T_11872 = _T_11871 ? _T_10366_9 : _T_11870; // @[Mux.scala 46:16:@9217.4]
  assign _T_11873 = 4'h9 == _T_11317_14; // @[Mux.scala 46:19:@9218.4]
  assign _T_11874 = _T_11873 ? _T_10366_8 : _T_11872; // @[Mux.scala 46:16:@9219.4]
  assign _T_11875 = 4'h8 == _T_11317_14; // @[Mux.scala 46:19:@9220.4]
  assign _T_11876 = _T_11875 ? _T_10366_7 : _T_11874; // @[Mux.scala 46:16:@9221.4]
  assign _T_11877 = 4'h7 == _T_11317_14; // @[Mux.scala 46:19:@9222.4]
  assign _T_11878 = _T_11877 ? _T_10366_6 : _T_11876; // @[Mux.scala 46:16:@9223.4]
  assign _T_11879 = 4'h6 == _T_11317_14; // @[Mux.scala 46:19:@9224.4]
  assign _T_11880 = _T_11879 ? _T_10366_5 : _T_11878; // @[Mux.scala 46:16:@9225.4]
  assign _T_11881 = 4'h5 == _T_11317_14; // @[Mux.scala 46:19:@9226.4]
  assign _T_11882 = _T_11881 ? _T_10366_4 : _T_11880; // @[Mux.scala 46:16:@9227.4]
  assign _T_11883 = 4'h4 == _T_11317_14; // @[Mux.scala 46:19:@9228.4]
  assign _T_11884 = _T_11883 ? _T_10366_3 : _T_11882; // @[Mux.scala 46:16:@9229.4]
  assign _T_11885 = 4'h3 == _T_11317_14; // @[Mux.scala 46:19:@9230.4]
  assign _T_11886 = _T_11885 ? _T_10366_2 : _T_11884; // @[Mux.scala 46:16:@9231.4]
  assign _T_11887 = 4'h2 == _T_11317_14; // @[Mux.scala 46:19:@9232.4]
  assign _T_11888 = _T_11887 ? _T_10366_1 : _T_11886; // @[Mux.scala 46:16:@9233.4]
  assign _T_11889 = 4'h1 == _T_11317_14; // @[Mux.scala 46:19:@9234.4]
  assign _T_11890 = _T_11889 ? _T_10366_0 : _T_11888; // @[Mux.scala 46:16:@9235.4]
  assign _T_11908 = 5'h10 == _T_11317_15; // @[Mux.scala 46:19:@9237.4]
  assign _T_11909 = _T_11908 ? _T_10366_15 : 8'h0; // @[Mux.scala 46:16:@9238.4]
  assign _T_11910 = 5'hf == _T_11317_15; // @[Mux.scala 46:19:@9239.4]
  assign _T_11911 = _T_11910 ? _T_10366_14 : _T_11909; // @[Mux.scala 46:16:@9240.4]
  assign _T_11912 = 5'he == _T_11317_15; // @[Mux.scala 46:19:@9241.4]
  assign _T_11913 = _T_11912 ? _T_10366_13 : _T_11911; // @[Mux.scala 46:16:@9242.4]
  assign _T_11914 = 5'hd == _T_11317_15; // @[Mux.scala 46:19:@9243.4]
  assign _T_11915 = _T_11914 ? _T_10366_12 : _T_11913; // @[Mux.scala 46:16:@9244.4]
  assign _T_11916 = 5'hc == _T_11317_15; // @[Mux.scala 46:19:@9245.4]
  assign _T_11917 = _T_11916 ? _T_10366_11 : _T_11915; // @[Mux.scala 46:16:@9246.4]
  assign _T_11918 = 5'hb == _T_11317_15; // @[Mux.scala 46:19:@9247.4]
  assign _T_11919 = _T_11918 ? _T_10366_10 : _T_11917; // @[Mux.scala 46:16:@9248.4]
  assign _T_11920 = 5'ha == _T_11317_15; // @[Mux.scala 46:19:@9249.4]
  assign _T_11921 = _T_11920 ? _T_10366_9 : _T_11919; // @[Mux.scala 46:16:@9250.4]
  assign _T_11922 = 5'h9 == _T_11317_15; // @[Mux.scala 46:19:@9251.4]
  assign _T_11923 = _T_11922 ? _T_10366_8 : _T_11921; // @[Mux.scala 46:16:@9252.4]
  assign _T_11924 = 5'h8 == _T_11317_15; // @[Mux.scala 46:19:@9253.4]
  assign _T_11925 = _T_11924 ? _T_10366_7 : _T_11923; // @[Mux.scala 46:16:@9254.4]
  assign _T_11926 = 5'h7 == _T_11317_15; // @[Mux.scala 46:19:@9255.4]
  assign _T_11927 = _T_11926 ? _T_10366_6 : _T_11925; // @[Mux.scala 46:16:@9256.4]
  assign _T_11928 = 5'h6 == _T_11317_15; // @[Mux.scala 46:19:@9257.4]
  assign _T_11929 = _T_11928 ? _T_10366_5 : _T_11927; // @[Mux.scala 46:16:@9258.4]
  assign _T_11930 = 5'h5 == _T_11317_15; // @[Mux.scala 46:19:@9259.4]
  assign _T_11931 = _T_11930 ? _T_10366_4 : _T_11929; // @[Mux.scala 46:16:@9260.4]
  assign _T_11932 = 5'h4 == _T_11317_15; // @[Mux.scala 46:19:@9261.4]
  assign _T_11933 = _T_11932 ? _T_10366_3 : _T_11931; // @[Mux.scala 46:16:@9262.4]
  assign _T_11934 = 5'h3 == _T_11317_15; // @[Mux.scala 46:19:@9263.4]
  assign _T_11935 = _T_11934 ? _T_10366_2 : _T_11933; // @[Mux.scala 46:16:@9264.4]
  assign _T_11936 = 5'h2 == _T_11317_15; // @[Mux.scala 46:19:@9265.4]
  assign _T_11937 = _T_11936 ? _T_10366_1 : _T_11935; // @[Mux.scala 46:16:@9266.4]
  assign _T_11938 = 5'h1 == _T_11317_15; // @[Mux.scala 46:19:@9267.4]
  assign _T_11939 = _T_11938 ? _T_10366_0 : _T_11937; // @[Mux.scala 46:16:@9268.4]
  assign _T_11958 = 5'h11 == _T_11317_16; // @[Mux.scala 46:19:@9270.4]
  assign _T_11959 = _T_11958 ? _T_10366_16 : 8'h0; // @[Mux.scala 46:16:@9271.4]
  assign _T_11960 = 5'h10 == _T_11317_16; // @[Mux.scala 46:19:@9272.4]
  assign _T_11961 = _T_11960 ? _T_10366_15 : _T_11959; // @[Mux.scala 46:16:@9273.4]
  assign _T_11962 = 5'hf == _T_11317_16; // @[Mux.scala 46:19:@9274.4]
  assign _T_11963 = _T_11962 ? _T_10366_14 : _T_11961; // @[Mux.scala 46:16:@9275.4]
  assign _T_11964 = 5'he == _T_11317_16; // @[Mux.scala 46:19:@9276.4]
  assign _T_11965 = _T_11964 ? _T_10366_13 : _T_11963; // @[Mux.scala 46:16:@9277.4]
  assign _T_11966 = 5'hd == _T_11317_16; // @[Mux.scala 46:19:@9278.4]
  assign _T_11967 = _T_11966 ? _T_10366_12 : _T_11965; // @[Mux.scala 46:16:@9279.4]
  assign _T_11968 = 5'hc == _T_11317_16; // @[Mux.scala 46:19:@9280.4]
  assign _T_11969 = _T_11968 ? _T_10366_11 : _T_11967; // @[Mux.scala 46:16:@9281.4]
  assign _T_11970 = 5'hb == _T_11317_16; // @[Mux.scala 46:19:@9282.4]
  assign _T_11971 = _T_11970 ? _T_10366_10 : _T_11969; // @[Mux.scala 46:16:@9283.4]
  assign _T_11972 = 5'ha == _T_11317_16; // @[Mux.scala 46:19:@9284.4]
  assign _T_11973 = _T_11972 ? _T_10366_9 : _T_11971; // @[Mux.scala 46:16:@9285.4]
  assign _T_11974 = 5'h9 == _T_11317_16; // @[Mux.scala 46:19:@9286.4]
  assign _T_11975 = _T_11974 ? _T_10366_8 : _T_11973; // @[Mux.scala 46:16:@9287.4]
  assign _T_11976 = 5'h8 == _T_11317_16; // @[Mux.scala 46:19:@9288.4]
  assign _T_11977 = _T_11976 ? _T_10366_7 : _T_11975; // @[Mux.scala 46:16:@9289.4]
  assign _T_11978 = 5'h7 == _T_11317_16; // @[Mux.scala 46:19:@9290.4]
  assign _T_11979 = _T_11978 ? _T_10366_6 : _T_11977; // @[Mux.scala 46:16:@9291.4]
  assign _T_11980 = 5'h6 == _T_11317_16; // @[Mux.scala 46:19:@9292.4]
  assign _T_11981 = _T_11980 ? _T_10366_5 : _T_11979; // @[Mux.scala 46:16:@9293.4]
  assign _T_11982 = 5'h5 == _T_11317_16; // @[Mux.scala 46:19:@9294.4]
  assign _T_11983 = _T_11982 ? _T_10366_4 : _T_11981; // @[Mux.scala 46:16:@9295.4]
  assign _T_11984 = 5'h4 == _T_11317_16; // @[Mux.scala 46:19:@9296.4]
  assign _T_11985 = _T_11984 ? _T_10366_3 : _T_11983; // @[Mux.scala 46:16:@9297.4]
  assign _T_11986 = 5'h3 == _T_11317_16; // @[Mux.scala 46:19:@9298.4]
  assign _T_11987 = _T_11986 ? _T_10366_2 : _T_11985; // @[Mux.scala 46:16:@9299.4]
  assign _T_11988 = 5'h2 == _T_11317_16; // @[Mux.scala 46:19:@9300.4]
  assign _T_11989 = _T_11988 ? _T_10366_1 : _T_11987; // @[Mux.scala 46:16:@9301.4]
  assign _T_11990 = 5'h1 == _T_11317_16; // @[Mux.scala 46:19:@9302.4]
  assign _T_11991 = _T_11990 ? _T_10366_0 : _T_11989; // @[Mux.scala 46:16:@9303.4]
  assign _T_12011 = 5'h12 == _T_11317_17; // @[Mux.scala 46:19:@9305.4]
  assign _T_12012 = _T_12011 ? _T_10366_17 : 8'h0; // @[Mux.scala 46:16:@9306.4]
  assign _T_12013 = 5'h11 == _T_11317_17; // @[Mux.scala 46:19:@9307.4]
  assign _T_12014 = _T_12013 ? _T_10366_16 : _T_12012; // @[Mux.scala 46:16:@9308.4]
  assign _T_12015 = 5'h10 == _T_11317_17; // @[Mux.scala 46:19:@9309.4]
  assign _T_12016 = _T_12015 ? _T_10366_15 : _T_12014; // @[Mux.scala 46:16:@9310.4]
  assign _T_12017 = 5'hf == _T_11317_17; // @[Mux.scala 46:19:@9311.4]
  assign _T_12018 = _T_12017 ? _T_10366_14 : _T_12016; // @[Mux.scala 46:16:@9312.4]
  assign _T_12019 = 5'he == _T_11317_17; // @[Mux.scala 46:19:@9313.4]
  assign _T_12020 = _T_12019 ? _T_10366_13 : _T_12018; // @[Mux.scala 46:16:@9314.4]
  assign _T_12021 = 5'hd == _T_11317_17; // @[Mux.scala 46:19:@9315.4]
  assign _T_12022 = _T_12021 ? _T_10366_12 : _T_12020; // @[Mux.scala 46:16:@9316.4]
  assign _T_12023 = 5'hc == _T_11317_17; // @[Mux.scala 46:19:@9317.4]
  assign _T_12024 = _T_12023 ? _T_10366_11 : _T_12022; // @[Mux.scala 46:16:@9318.4]
  assign _T_12025 = 5'hb == _T_11317_17; // @[Mux.scala 46:19:@9319.4]
  assign _T_12026 = _T_12025 ? _T_10366_10 : _T_12024; // @[Mux.scala 46:16:@9320.4]
  assign _T_12027 = 5'ha == _T_11317_17; // @[Mux.scala 46:19:@9321.4]
  assign _T_12028 = _T_12027 ? _T_10366_9 : _T_12026; // @[Mux.scala 46:16:@9322.4]
  assign _T_12029 = 5'h9 == _T_11317_17; // @[Mux.scala 46:19:@9323.4]
  assign _T_12030 = _T_12029 ? _T_10366_8 : _T_12028; // @[Mux.scala 46:16:@9324.4]
  assign _T_12031 = 5'h8 == _T_11317_17; // @[Mux.scala 46:19:@9325.4]
  assign _T_12032 = _T_12031 ? _T_10366_7 : _T_12030; // @[Mux.scala 46:16:@9326.4]
  assign _T_12033 = 5'h7 == _T_11317_17; // @[Mux.scala 46:19:@9327.4]
  assign _T_12034 = _T_12033 ? _T_10366_6 : _T_12032; // @[Mux.scala 46:16:@9328.4]
  assign _T_12035 = 5'h6 == _T_11317_17; // @[Mux.scala 46:19:@9329.4]
  assign _T_12036 = _T_12035 ? _T_10366_5 : _T_12034; // @[Mux.scala 46:16:@9330.4]
  assign _T_12037 = 5'h5 == _T_11317_17; // @[Mux.scala 46:19:@9331.4]
  assign _T_12038 = _T_12037 ? _T_10366_4 : _T_12036; // @[Mux.scala 46:16:@9332.4]
  assign _T_12039 = 5'h4 == _T_11317_17; // @[Mux.scala 46:19:@9333.4]
  assign _T_12040 = _T_12039 ? _T_10366_3 : _T_12038; // @[Mux.scala 46:16:@9334.4]
  assign _T_12041 = 5'h3 == _T_11317_17; // @[Mux.scala 46:19:@9335.4]
  assign _T_12042 = _T_12041 ? _T_10366_2 : _T_12040; // @[Mux.scala 46:16:@9336.4]
  assign _T_12043 = 5'h2 == _T_11317_17; // @[Mux.scala 46:19:@9337.4]
  assign _T_12044 = _T_12043 ? _T_10366_1 : _T_12042; // @[Mux.scala 46:16:@9338.4]
  assign _T_12045 = 5'h1 == _T_11317_17; // @[Mux.scala 46:19:@9339.4]
  assign _T_12046 = _T_12045 ? _T_10366_0 : _T_12044; // @[Mux.scala 46:16:@9340.4]
  assign _T_12067 = 5'h13 == _T_11317_18; // @[Mux.scala 46:19:@9342.4]
  assign _T_12068 = _T_12067 ? _T_10366_18 : 8'h0; // @[Mux.scala 46:16:@9343.4]
  assign _T_12069 = 5'h12 == _T_11317_18; // @[Mux.scala 46:19:@9344.4]
  assign _T_12070 = _T_12069 ? _T_10366_17 : _T_12068; // @[Mux.scala 46:16:@9345.4]
  assign _T_12071 = 5'h11 == _T_11317_18; // @[Mux.scala 46:19:@9346.4]
  assign _T_12072 = _T_12071 ? _T_10366_16 : _T_12070; // @[Mux.scala 46:16:@9347.4]
  assign _T_12073 = 5'h10 == _T_11317_18; // @[Mux.scala 46:19:@9348.4]
  assign _T_12074 = _T_12073 ? _T_10366_15 : _T_12072; // @[Mux.scala 46:16:@9349.4]
  assign _T_12075 = 5'hf == _T_11317_18; // @[Mux.scala 46:19:@9350.4]
  assign _T_12076 = _T_12075 ? _T_10366_14 : _T_12074; // @[Mux.scala 46:16:@9351.4]
  assign _T_12077 = 5'he == _T_11317_18; // @[Mux.scala 46:19:@9352.4]
  assign _T_12078 = _T_12077 ? _T_10366_13 : _T_12076; // @[Mux.scala 46:16:@9353.4]
  assign _T_12079 = 5'hd == _T_11317_18; // @[Mux.scala 46:19:@9354.4]
  assign _T_12080 = _T_12079 ? _T_10366_12 : _T_12078; // @[Mux.scala 46:16:@9355.4]
  assign _T_12081 = 5'hc == _T_11317_18; // @[Mux.scala 46:19:@9356.4]
  assign _T_12082 = _T_12081 ? _T_10366_11 : _T_12080; // @[Mux.scala 46:16:@9357.4]
  assign _T_12083 = 5'hb == _T_11317_18; // @[Mux.scala 46:19:@9358.4]
  assign _T_12084 = _T_12083 ? _T_10366_10 : _T_12082; // @[Mux.scala 46:16:@9359.4]
  assign _T_12085 = 5'ha == _T_11317_18; // @[Mux.scala 46:19:@9360.4]
  assign _T_12086 = _T_12085 ? _T_10366_9 : _T_12084; // @[Mux.scala 46:16:@9361.4]
  assign _T_12087 = 5'h9 == _T_11317_18; // @[Mux.scala 46:19:@9362.4]
  assign _T_12088 = _T_12087 ? _T_10366_8 : _T_12086; // @[Mux.scala 46:16:@9363.4]
  assign _T_12089 = 5'h8 == _T_11317_18; // @[Mux.scala 46:19:@9364.4]
  assign _T_12090 = _T_12089 ? _T_10366_7 : _T_12088; // @[Mux.scala 46:16:@9365.4]
  assign _T_12091 = 5'h7 == _T_11317_18; // @[Mux.scala 46:19:@9366.4]
  assign _T_12092 = _T_12091 ? _T_10366_6 : _T_12090; // @[Mux.scala 46:16:@9367.4]
  assign _T_12093 = 5'h6 == _T_11317_18; // @[Mux.scala 46:19:@9368.4]
  assign _T_12094 = _T_12093 ? _T_10366_5 : _T_12092; // @[Mux.scala 46:16:@9369.4]
  assign _T_12095 = 5'h5 == _T_11317_18; // @[Mux.scala 46:19:@9370.4]
  assign _T_12096 = _T_12095 ? _T_10366_4 : _T_12094; // @[Mux.scala 46:16:@9371.4]
  assign _T_12097 = 5'h4 == _T_11317_18; // @[Mux.scala 46:19:@9372.4]
  assign _T_12098 = _T_12097 ? _T_10366_3 : _T_12096; // @[Mux.scala 46:16:@9373.4]
  assign _T_12099 = 5'h3 == _T_11317_18; // @[Mux.scala 46:19:@9374.4]
  assign _T_12100 = _T_12099 ? _T_10366_2 : _T_12098; // @[Mux.scala 46:16:@9375.4]
  assign _T_12101 = 5'h2 == _T_11317_18; // @[Mux.scala 46:19:@9376.4]
  assign _T_12102 = _T_12101 ? _T_10366_1 : _T_12100; // @[Mux.scala 46:16:@9377.4]
  assign _T_12103 = 5'h1 == _T_11317_18; // @[Mux.scala 46:19:@9378.4]
  assign _T_12104 = _T_12103 ? _T_10366_0 : _T_12102; // @[Mux.scala 46:16:@9379.4]
  assign _T_12126 = 5'h14 == _T_11317_19; // @[Mux.scala 46:19:@9381.4]
  assign _T_12127 = _T_12126 ? _T_10366_19 : 8'h0; // @[Mux.scala 46:16:@9382.4]
  assign _T_12128 = 5'h13 == _T_11317_19; // @[Mux.scala 46:19:@9383.4]
  assign _T_12129 = _T_12128 ? _T_10366_18 : _T_12127; // @[Mux.scala 46:16:@9384.4]
  assign _T_12130 = 5'h12 == _T_11317_19; // @[Mux.scala 46:19:@9385.4]
  assign _T_12131 = _T_12130 ? _T_10366_17 : _T_12129; // @[Mux.scala 46:16:@9386.4]
  assign _T_12132 = 5'h11 == _T_11317_19; // @[Mux.scala 46:19:@9387.4]
  assign _T_12133 = _T_12132 ? _T_10366_16 : _T_12131; // @[Mux.scala 46:16:@9388.4]
  assign _T_12134 = 5'h10 == _T_11317_19; // @[Mux.scala 46:19:@9389.4]
  assign _T_12135 = _T_12134 ? _T_10366_15 : _T_12133; // @[Mux.scala 46:16:@9390.4]
  assign _T_12136 = 5'hf == _T_11317_19; // @[Mux.scala 46:19:@9391.4]
  assign _T_12137 = _T_12136 ? _T_10366_14 : _T_12135; // @[Mux.scala 46:16:@9392.4]
  assign _T_12138 = 5'he == _T_11317_19; // @[Mux.scala 46:19:@9393.4]
  assign _T_12139 = _T_12138 ? _T_10366_13 : _T_12137; // @[Mux.scala 46:16:@9394.4]
  assign _T_12140 = 5'hd == _T_11317_19; // @[Mux.scala 46:19:@9395.4]
  assign _T_12141 = _T_12140 ? _T_10366_12 : _T_12139; // @[Mux.scala 46:16:@9396.4]
  assign _T_12142 = 5'hc == _T_11317_19; // @[Mux.scala 46:19:@9397.4]
  assign _T_12143 = _T_12142 ? _T_10366_11 : _T_12141; // @[Mux.scala 46:16:@9398.4]
  assign _T_12144 = 5'hb == _T_11317_19; // @[Mux.scala 46:19:@9399.4]
  assign _T_12145 = _T_12144 ? _T_10366_10 : _T_12143; // @[Mux.scala 46:16:@9400.4]
  assign _T_12146 = 5'ha == _T_11317_19; // @[Mux.scala 46:19:@9401.4]
  assign _T_12147 = _T_12146 ? _T_10366_9 : _T_12145; // @[Mux.scala 46:16:@9402.4]
  assign _T_12148 = 5'h9 == _T_11317_19; // @[Mux.scala 46:19:@9403.4]
  assign _T_12149 = _T_12148 ? _T_10366_8 : _T_12147; // @[Mux.scala 46:16:@9404.4]
  assign _T_12150 = 5'h8 == _T_11317_19; // @[Mux.scala 46:19:@9405.4]
  assign _T_12151 = _T_12150 ? _T_10366_7 : _T_12149; // @[Mux.scala 46:16:@9406.4]
  assign _T_12152 = 5'h7 == _T_11317_19; // @[Mux.scala 46:19:@9407.4]
  assign _T_12153 = _T_12152 ? _T_10366_6 : _T_12151; // @[Mux.scala 46:16:@9408.4]
  assign _T_12154 = 5'h6 == _T_11317_19; // @[Mux.scala 46:19:@9409.4]
  assign _T_12155 = _T_12154 ? _T_10366_5 : _T_12153; // @[Mux.scala 46:16:@9410.4]
  assign _T_12156 = 5'h5 == _T_11317_19; // @[Mux.scala 46:19:@9411.4]
  assign _T_12157 = _T_12156 ? _T_10366_4 : _T_12155; // @[Mux.scala 46:16:@9412.4]
  assign _T_12158 = 5'h4 == _T_11317_19; // @[Mux.scala 46:19:@9413.4]
  assign _T_12159 = _T_12158 ? _T_10366_3 : _T_12157; // @[Mux.scala 46:16:@9414.4]
  assign _T_12160 = 5'h3 == _T_11317_19; // @[Mux.scala 46:19:@9415.4]
  assign _T_12161 = _T_12160 ? _T_10366_2 : _T_12159; // @[Mux.scala 46:16:@9416.4]
  assign _T_12162 = 5'h2 == _T_11317_19; // @[Mux.scala 46:19:@9417.4]
  assign _T_12163 = _T_12162 ? _T_10366_1 : _T_12161; // @[Mux.scala 46:16:@9418.4]
  assign _T_12164 = 5'h1 == _T_11317_19; // @[Mux.scala 46:19:@9419.4]
  assign _T_12165 = _T_12164 ? _T_10366_0 : _T_12163; // @[Mux.scala 46:16:@9420.4]
  assign _T_12188 = 5'h15 == _T_11317_20; // @[Mux.scala 46:19:@9422.4]
  assign _T_12189 = _T_12188 ? _T_10366_20 : 8'h0; // @[Mux.scala 46:16:@9423.4]
  assign _T_12190 = 5'h14 == _T_11317_20; // @[Mux.scala 46:19:@9424.4]
  assign _T_12191 = _T_12190 ? _T_10366_19 : _T_12189; // @[Mux.scala 46:16:@9425.4]
  assign _T_12192 = 5'h13 == _T_11317_20; // @[Mux.scala 46:19:@9426.4]
  assign _T_12193 = _T_12192 ? _T_10366_18 : _T_12191; // @[Mux.scala 46:16:@9427.4]
  assign _T_12194 = 5'h12 == _T_11317_20; // @[Mux.scala 46:19:@9428.4]
  assign _T_12195 = _T_12194 ? _T_10366_17 : _T_12193; // @[Mux.scala 46:16:@9429.4]
  assign _T_12196 = 5'h11 == _T_11317_20; // @[Mux.scala 46:19:@9430.4]
  assign _T_12197 = _T_12196 ? _T_10366_16 : _T_12195; // @[Mux.scala 46:16:@9431.4]
  assign _T_12198 = 5'h10 == _T_11317_20; // @[Mux.scala 46:19:@9432.4]
  assign _T_12199 = _T_12198 ? _T_10366_15 : _T_12197; // @[Mux.scala 46:16:@9433.4]
  assign _T_12200 = 5'hf == _T_11317_20; // @[Mux.scala 46:19:@9434.4]
  assign _T_12201 = _T_12200 ? _T_10366_14 : _T_12199; // @[Mux.scala 46:16:@9435.4]
  assign _T_12202 = 5'he == _T_11317_20; // @[Mux.scala 46:19:@9436.4]
  assign _T_12203 = _T_12202 ? _T_10366_13 : _T_12201; // @[Mux.scala 46:16:@9437.4]
  assign _T_12204 = 5'hd == _T_11317_20; // @[Mux.scala 46:19:@9438.4]
  assign _T_12205 = _T_12204 ? _T_10366_12 : _T_12203; // @[Mux.scala 46:16:@9439.4]
  assign _T_12206 = 5'hc == _T_11317_20; // @[Mux.scala 46:19:@9440.4]
  assign _T_12207 = _T_12206 ? _T_10366_11 : _T_12205; // @[Mux.scala 46:16:@9441.4]
  assign _T_12208 = 5'hb == _T_11317_20; // @[Mux.scala 46:19:@9442.4]
  assign _T_12209 = _T_12208 ? _T_10366_10 : _T_12207; // @[Mux.scala 46:16:@9443.4]
  assign _T_12210 = 5'ha == _T_11317_20; // @[Mux.scala 46:19:@9444.4]
  assign _T_12211 = _T_12210 ? _T_10366_9 : _T_12209; // @[Mux.scala 46:16:@9445.4]
  assign _T_12212 = 5'h9 == _T_11317_20; // @[Mux.scala 46:19:@9446.4]
  assign _T_12213 = _T_12212 ? _T_10366_8 : _T_12211; // @[Mux.scala 46:16:@9447.4]
  assign _T_12214 = 5'h8 == _T_11317_20; // @[Mux.scala 46:19:@9448.4]
  assign _T_12215 = _T_12214 ? _T_10366_7 : _T_12213; // @[Mux.scala 46:16:@9449.4]
  assign _T_12216 = 5'h7 == _T_11317_20; // @[Mux.scala 46:19:@9450.4]
  assign _T_12217 = _T_12216 ? _T_10366_6 : _T_12215; // @[Mux.scala 46:16:@9451.4]
  assign _T_12218 = 5'h6 == _T_11317_20; // @[Mux.scala 46:19:@9452.4]
  assign _T_12219 = _T_12218 ? _T_10366_5 : _T_12217; // @[Mux.scala 46:16:@9453.4]
  assign _T_12220 = 5'h5 == _T_11317_20; // @[Mux.scala 46:19:@9454.4]
  assign _T_12221 = _T_12220 ? _T_10366_4 : _T_12219; // @[Mux.scala 46:16:@9455.4]
  assign _T_12222 = 5'h4 == _T_11317_20; // @[Mux.scala 46:19:@9456.4]
  assign _T_12223 = _T_12222 ? _T_10366_3 : _T_12221; // @[Mux.scala 46:16:@9457.4]
  assign _T_12224 = 5'h3 == _T_11317_20; // @[Mux.scala 46:19:@9458.4]
  assign _T_12225 = _T_12224 ? _T_10366_2 : _T_12223; // @[Mux.scala 46:16:@9459.4]
  assign _T_12226 = 5'h2 == _T_11317_20; // @[Mux.scala 46:19:@9460.4]
  assign _T_12227 = _T_12226 ? _T_10366_1 : _T_12225; // @[Mux.scala 46:16:@9461.4]
  assign _T_12228 = 5'h1 == _T_11317_20; // @[Mux.scala 46:19:@9462.4]
  assign _T_12229 = _T_12228 ? _T_10366_0 : _T_12227; // @[Mux.scala 46:16:@9463.4]
  assign _T_12253 = 5'h16 == _T_11317_21; // @[Mux.scala 46:19:@9465.4]
  assign _T_12254 = _T_12253 ? _T_10366_21 : 8'h0; // @[Mux.scala 46:16:@9466.4]
  assign _T_12255 = 5'h15 == _T_11317_21; // @[Mux.scala 46:19:@9467.4]
  assign _T_12256 = _T_12255 ? _T_10366_20 : _T_12254; // @[Mux.scala 46:16:@9468.4]
  assign _T_12257 = 5'h14 == _T_11317_21; // @[Mux.scala 46:19:@9469.4]
  assign _T_12258 = _T_12257 ? _T_10366_19 : _T_12256; // @[Mux.scala 46:16:@9470.4]
  assign _T_12259 = 5'h13 == _T_11317_21; // @[Mux.scala 46:19:@9471.4]
  assign _T_12260 = _T_12259 ? _T_10366_18 : _T_12258; // @[Mux.scala 46:16:@9472.4]
  assign _T_12261 = 5'h12 == _T_11317_21; // @[Mux.scala 46:19:@9473.4]
  assign _T_12262 = _T_12261 ? _T_10366_17 : _T_12260; // @[Mux.scala 46:16:@9474.4]
  assign _T_12263 = 5'h11 == _T_11317_21; // @[Mux.scala 46:19:@9475.4]
  assign _T_12264 = _T_12263 ? _T_10366_16 : _T_12262; // @[Mux.scala 46:16:@9476.4]
  assign _T_12265 = 5'h10 == _T_11317_21; // @[Mux.scala 46:19:@9477.4]
  assign _T_12266 = _T_12265 ? _T_10366_15 : _T_12264; // @[Mux.scala 46:16:@9478.4]
  assign _T_12267 = 5'hf == _T_11317_21; // @[Mux.scala 46:19:@9479.4]
  assign _T_12268 = _T_12267 ? _T_10366_14 : _T_12266; // @[Mux.scala 46:16:@9480.4]
  assign _T_12269 = 5'he == _T_11317_21; // @[Mux.scala 46:19:@9481.4]
  assign _T_12270 = _T_12269 ? _T_10366_13 : _T_12268; // @[Mux.scala 46:16:@9482.4]
  assign _T_12271 = 5'hd == _T_11317_21; // @[Mux.scala 46:19:@9483.4]
  assign _T_12272 = _T_12271 ? _T_10366_12 : _T_12270; // @[Mux.scala 46:16:@9484.4]
  assign _T_12273 = 5'hc == _T_11317_21; // @[Mux.scala 46:19:@9485.4]
  assign _T_12274 = _T_12273 ? _T_10366_11 : _T_12272; // @[Mux.scala 46:16:@9486.4]
  assign _T_12275 = 5'hb == _T_11317_21; // @[Mux.scala 46:19:@9487.4]
  assign _T_12276 = _T_12275 ? _T_10366_10 : _T_12274; // @[Mux.scala 46:16:@9488.4]
  assign _T_12277 = 5'ha == _T_11317_21; // @[Mux.scala 46:19:@9489.4]
  assign _T_12278 = _T_12277 ? _T_10366_9 : _T_12276; // @[Mux.scala 46:16:@9490.4]
  assign _T_12279 = 5'h9 == _T_11317_21; // @[Mux.scala 46:19:@9491.4]
  assign _T_12280 = _T_12279 ? _T_10366_8 : _T_12278; // @[Mux.scala 46:16:@9492.4]
  assign _T_12281 = 5'h8 == _T_11317_21; // @[Mux.scala 46:19:@9493.4]
  assign _T_12282 = _T_12281 ? _T_10366_7 : _T_12280; // @[Mux.scala 46:16:@9494.4]
  assign _T_12283 = 5'h7 == _T_11317_21; // @[Mux.scala 46:19:@9495.4]
  assign _T_12284 = _T_12283 ? _T_10366_6 : _T_12282; // @[Mux.scala 46:16:@9496.4]
  assign _T_12285 = 5'h6 == _T_11317_21; // @[Mux.scala 46:19:@9497.4]
  assign _T_12286 = _T_12285 ? _T_10366_5 : _T_12284; // @[Mux.scala 46:16:@9498.4]
  assign _T_12287 = 5'h5 == _T_11317_21; // @[Mux.scala 46:19:@9499.4]
  assign _T_12288 = _T_12287 ? _T_10366_4 : _T_12286; // @[Mux.scala 46:16:@9500.4]
  assign _T_12289 = 5'h4 == _T_11317_21; // @[Mux.scala 46:19:@9501.4]
  assign _T_12290 = _T_12289 ? _T_10366_3 : _T_12288; // @[Mux.scala 46:16:@9502.4]
  assign _T_12291 = 5'h3 == _T_11317_21; // @[Mux.scala 46:19:@9503.4]
  assign _T_12292 = _T_12291 ? _T_10366_2 : _T_12290; // @[Mux.scala 46:16:@9504.4]
  assign _T_12293 = 5'h2 == _T_11317_21; // @[Mux.scala 46:19:@9505.4]
  assign _T_12294 = _T_12293 ? _T_10366_1 : _T_12292; // @[Mux.scala 46:16:@9506.4]
  assign _T_12295 = 5'h1 == _T_11317_21; // @[Mux.scala 46:19:@9507.4]
  assign _T_12296 = _T_12295 ? _T_10366_0 : _T_12294; // @[Mux.scala 46:16:@9508.4]
  assign _T_12321 = 5'h17 == _T_11317_22; // @[Mux.scala 46:19:@9510.4]
  assign _T_12322 = _T_12321 ? _T_10366_22 : 8'h0; // @[Mux.scala 46:16:@9511.4]
  assign _T_12323 = 5'h16 == _T_11317_22; // @[Mux.scala 46:19:@9512.4]
  assign _T_12324 = _T_12323 ? _T_10366_21 : _T_12322; // @[Mux.scala 46:16:@9513.4]
  assign _T_12325 = 5'h15 == _T_11317_22; // @[Mux.scala 46:19:@9514.4]
  assign _T_12326 = _T_12325 ? _T_10366_20 : _T_12324; // @[Mux.scala 46:16:@9515.4]
  assign _T_12327 = 5'h14 == _T_11317_22; // @[Mux.scala 46:19:@9516.4]
  assign _T_12328 = _T_12327 ? _T_10366_19 : _T_12326; // @[Mux.scala 46:16:@9517.4]
  assign _T_12329 = 5'h13 == _T_11317_22; // @[Mux.scala 46:19:@9518.4]
  assign _T_12330 = _T_12329 ? _T_10366_18 : _T_12328; // @[Mux.scala 46:16:@9519.4]
  assign _T_12331 = 5'h12 == _T_11317_22; // @[Mux.scala 46:19:@9520.4]
  assign _T_12332 = _T_12331 ? _T_10366_17 : _T_12330; // @[Mux.scala 46:16:@9521.4]
  assign _T_12333 = 5'h11 == _T_11317_22; // @[Mux.scala 46:19:@9522.4]
  assign _T_12334 = _T_12333 ? _T_10366_16 : _T_12332; // @[Mux.scala 46:16:@9523.4]
  assign _T_12335 = 5'h10 == _T_11317_22; // @[Mux.scala 46:19:@9524.4]
  assign _T_12336 = _T_12335 ? _T_10366_15 : _T_12334; // @[Mux.scala 46:16:@9525.4]
  assign _T_12337 = 5'hf == _T_11317_22; // @[Mux.scala 46:19:@9526.4]
  assign _T_12338 = _T_12337 ? _T_10366_14 : _T_12336; // @[Mux.scala 46:16:@9527.4]
  assign _T_12339 = 5'he == _T_11317_22; // @[Mux.scala 46:19:@9528.4]
  assign _T_12340 = _T_12339 ? _T_10366_13 : _T_12338; // @[Mux.scala 46:16:@9529.4]
  assign _T_12341 = 5'hd == _T_11317_22; // @[Mux.scala 46:19:@9530.4]
  assign _T_12342 = _T_12341 ? _T_10366_12 : _T_12340; // @[Mux.scala 46:16:@9531.4]
  assign _T_12343 = 5'hc == _T_11317_22; // @[Mux.scala 46:19:@9532.4]
  assign _T_12344 = _T_12343 ? _T_10366_11 : _T_12342; // @[Mux.scala 46:16:@9533.4]
  assign _T_12345 = 5'hb == _T_11317_22; // @[Mux.scala 46:19:@9534.4]
  assign _T_12346 = _T_12345 ? _T_10366_10 : _T_12344; // @[Mux.scala 46:16:@9535.4]
  assign _T_12347 = 5'ha == _T_11317_22; // @[Mux.scala 46:19:@9536.4]
  assign _T_12348 = _T_12347 ? _T_10366_9 : _T_12346; // @[Mux.scala 46:16:@9537.4]
  assign _T_12349 = 5'h9 == _T_11317_22; // @[Mux.scala 46:19:@9538.4]
  assign _T_12350 = _T_12349 ? _T_10366_8 : _T_12348; // @[Mux.scala 46:16:@9539.4]
  assign _T_12351 = 5'h8 == _T_11317_22; // @[Mux.scala 46:19:@9540.4]
  assign _T_12352 = _T_12351 ? _T_10366_7 : _T_12350; // @[Mux.scala 46:16:@9541.4]
  assign _T_12353 = 5'h7 == _T_11317_22; // @[Mux.scala 46:19:@9542.4]
  assign _T_12354 = _T_12353 ? _T_10366_6 : _T_12352; // @[Mux.scala 46:16:@9543.4]
  assign _T_12355 = 5'h6 == _T_11317_22; // @[Mux.scala 46:19:@9544.4]
  assign _T_12356 = _T_12355 ? _T_10366_5 : _T_12354; // @[Mux.scala 46:16:@9545.4]
  assign _T_12357 = 5'h5 == _T_11317_22; // @[Mux.scala 46:19:@9546.4]
  assign _T_12358 = _T_12357 ? _T_10366_4 : _T_12356; // @[Mux.scala 46:16:@9547.4]
  assign _T_12359 = 5'h4 == _T_11317_22; // @[Mux.scala 46:19:@9548.4]
  assign _T_12360 = _T_12359 ? _T_10366_3 : _T_12358; // @[Mux.scala 46:16:@9549.4]
  assign _T_12361 = 5'h3 == _T_11317_22; // @[Mux.scala 46:19:@9550.4]
  assign _T_12362 = _T_12361 ? _T_10366_2 : _T_12360; // @[Mux.scala 46:16:@9551.4]
  assign _T_12363 = 5'h2 == _T_11317_22; // @[Mux.scala 46:19:@9552.4]
  assign _T_12364 = _T_12363 ? _T_10366_1 : _T_12362; // @[Mux.scala 46:16:@9553.4]
  assign _T_12365 = 5'h1 == _T_11317_22; // @[Mux.scala 46:19:@9554.4]
  assign _T_12366 = _T_12365 ? _T_10366_0 : _T_12364; // @[Mux.scala 46:16:@9555.4]
  assign _T_12392 = 5'h18 == _T_11317_23; // @[Mux.scala 46:19:@9557.4]
  assign _T_12393 = _T_12392 ? _T_10366_23 : 8'h0; // @[Mux.scala 46:16:@9558.4]
  assign _T_12394 = 5'h17 == _T_11317_23; // @[Mux.scala 46:19:@9559.4]
  assign _T_12395 = _T_12394 ? _T_10366_22 : _T_12393; // @[Mux.scala 46:16:@9560.4]
  assign _T_12396 = 5'h16 == _T_11317_23; // @[Mux.scala 46:19:@9561.4]
  assign _T_12397 = _T_12396 ? _T_10366_21 : _T_12395; // @[Mux.scala 46:16:@9562.4]
  assign _T_12398 = 5'h15 == _T_11317_23; // @[Mux.scala 46:19:@9563.4]
  assign _T_12399 = _T_12398 ? _T_10366_20 : _T_12397; // @[Mux.scala 46:16:@9564.4]
  assign _T_12400 = 5'h14 == _T_11317_23; // @[Mux.scala 46:19:@9565.4]
  assign _T_12401 = _T_12400 ? _T_10366_19 : _T_12399; // @[Mux.scala 46:16:@9566.4]
  assign _T_12402 = 5'h13 == _T_11317_23; // @[Mux.scala 46:19:@9567.4]
  assign _T_12403 = _T_12402 ? _T_10366_18 : _T_12401; // @[Mux.scala 46:16:@9568.4]
  assign _T_12404 = 5'h12 == _T_11317_23; // @[Mux.scala 46:19:@9569.4]
  assign _T_12405 = _T_12404 ? _T_10366_17 : _T_12403; // @[Mux.scala 46:16:@9570.4]
  assign _T_12406 = 5'h11 == _T_11317_23; // @[Mux.scala 46:19:@9571.4]
  assign _T_12407 = _T_12406 ? _T_10366_16 : _T_12405; // @[Mux.scala 46:16:@9572.4]
  assign _T_12408 = 5'h10 == _T_11317_23; // @[Mux.scala 46:19:@9573.4]
  assign _T_12409 = _T_12408 ? _T_10366_15 : _T_12407; // @[Mux.scala 46:16:@9574.4]
  assign _T_12410 = 5'hf == _T_11317_23; // @[Mux.scala 46:19:@9575.4]
  assign _T_12411 = _T_12410 ? _T_10366_14 : _T_12409; // @[Mux.scala 46:16:@9576.4]
  assign _T_12412 = 5'he == _T_11317_23; // @[Mux.scala 46:19:@9577.4]
  assign _T_12413 = _T_12412 ? _T_10366_13 : _T_12411; // @[Mux.scala 46:16:@9578.4]
  assign _T_12414 = 5'hd == _T_11317_23; // @[Mux.scala 46:19:@9579.4]
  assign _T_12415 = _T_12414 ? _T_10366_12 : _T_12413; // @[Mux.scala 46:16:@9580.4]
  assign _T_12416 = 5'hc == _T_11317_23; // @[Mux.scala 46:19:@9581.4]
  assign _T_12417 = _T_12416 ? _T_10366_11 : _T_12415; // @[Mux.scala 46:16:@9582.4]
  assign _T_12418 = 5'hb == _T_11317_23; // @[Mux.scala 46:19:@9583.4]
  assign _T_12419 = _T_12418 ? _T_10366_10 : _T_12417; // @[Mux.scala 46:16:@9584.4]
  assign _T_12420 = 5'ha == _T_11317_23; // @[Mux.scala 46:19:@9585.4]
  assign _T_12421 = _T_12420 ? _T_10366_9 : _T_12419; // @[Mux.scala 46:16:@9586.4]
  assign _T_12422 = 5'h9 == _T_11317_23; // @[Mux.scala 46:19:@9587.4]
  assign _T_12423 = _T_12422 ? _T_10366_8 : _T_12421; // @[Mux.scala 46:16:@9588.4]
  assign _T_12424 = 5'h8 == _T_11317_23; // @[Mux.scala 46:19:@9589.4]
  assign _T_12425 = _T_12424 ? _T_10366_7 : _T_12423; // @[Mux.scala 46:16:@9590.4]
  assign _T_12426 = 5'h7 == _T_11317_23; // @[Mux.scala 46:19:@9591.4]
  assign _T_12427 = _T_12426 ? _T_10366_6 : _T_12425; // @[Mux.scala 46:16:@9592.4]
  assign _T_12428 = 5'h6 == _T_11317_23; // @[Mux.scala 46:19:@9593.4]
  assign _T_12429 = _T_12428 ? _T_10366_5 : _T_12427; // @[Mux.scala 46:16:@9594.4]
  assign _T_12430 = 5'h5 == _T_11317_23; // @[Mux.scala 46:19:@9595.4]
  assign _T_12431 = _T_12430 ? _T_10366_4 : _T_12429; // @[Mux.scala 46:16:@9596.4]
  assign _T_12432 = 5'h4 == _T_11317_23; // @[Mux.scala 46:19:@9597.4]
  assign _T_12433 = _T_12432 ? _T_10366_3 : _T_12431; // @[Mux.scala 46:16:@9598.4]
  assign _T_12434 = 5'h3 == _T_11317_23; // @[Mux.scala 46:19:@9599.4]
  assign _T_12435 = _T_12434 ? _T_10366_2 : _T_12433; // @[Mux.scala 46:16:@9600.4]
  assign _T_12436 = 5'h2 == _T_11317_23; // @[Mux.scala 46:19:@9601.4]
  assign _T_12437 = _T_12436 ? _T_10366_1 : _T_12435; // @[Mux.scala 46:16:@9602.4]
  assign _T_12438 = 5'h1 == _T_11317_23; // @[Mux.scala 46:19:@9603.4]
  assign _T_12439 = _T_12438 ? _T_10366_0 : _T_12437; // @[Mux.scala 46:16:@9604.4]
  assign _T_12466 = 5'h19 == _T_11317_24; // @[Mux.scala 46:19:@9606.4]
  assign _T_12467 = _T_12466 ? _T_10366_24 : 8'h0; // @[Mux.scala 46:16:@9607.4]
  assign _T_12468 = 5'h18 == _T_11317_24; // @[Mux.scala 46:19:@9608.4]
  assign _T_12469 = _T_12468 ? _T_10366_23 : _T_12467; // @[Mux.scala 46:16:@9609.4]
  assign _T_12470 = 5'h17 == _T_11317_24; // @[Mux.scala 46:19:@9610.4]
  assign _T_12471 = _T_12470 ? _T_10366_22 : _T_12469; // @[Mux.scala 46:16:@9611.4]
  assign _T_12472 = 5'h16 == _T_11317_24; // @[Mux.scala 46:19:@9612.4]
  assign _T_12473 = _T_12472 ? _T_10366_21 : _T_12471; // @[Mux.scala 46:16:@9613.4]
  assign _T_12474 = 5'h15 == _T_11317_24; // @[Mux.scala 46:19:@9614.4]
  assign _T_12475 = _T_12474 ? _T_10366_20 : _T_12473; // @[Mux.scala 46:16:@9615.4]
  assign _T_12476 = 5'h14 == _T_11317_24; // @[Mux.scala 46:19:@9616.4]
  assign _T_12477 = _T_12476 ? _T_10366_19 : _T_12475; // @[Mux.scala 46:16:@9617.4]
  assign _T_12478 = 5'h13 == _T_11317_24; // @[Mux.scala 46:19:@9618.4]
  assign _T_12479 = _T_12478 ? _T_10366_18 : _T_12477; // @[Mux.scala 46:16:@9619.4]
  assign _T_12480 = 5'h12 == _T_11317_24; // @[Mux.scala 46:19:@9620.4]
  assign _T_12481 = _T_12480 ? _T_10366_17 : _T_12479; // @[Mux.scala 46:16:@9621.4]
  assign _T_12482 = 5'h11 == _T_11317_24; // @[Mux.scala 46:19:@9622.4]
  assign _T_12483 = _T_12482 ? _T_10366_16 : _T_12481; // @[Mux.scala 46:16:@9623.4]
  assign _T_12484 = 5'h10 == _T_11317_24; // @[Mux.scala 46:19:@9624.4]
  assign _T_12485 = _T_12484 ? _T_10366_15 : _T_12483; // @[Mux.scala 46:16:@9625.4]
  assign _T_12486 = 5'hf == _T_11317_24; // @[Mux.scala 46:19:@9626.4]
  assign _T_12487 = _T_12486 ? _T_10366_14 : _T_12485; // @[Mux.scala 46:16:@9627.4]
  assign _T_12488 = 5'he == _T_11317_24; // @[Mux.scala 46:19:@9628.4]
  assign _T_12489 = _T_12488 ? _T_10366_13 : _T_12487; // @[Mux.scala 46:16:@9629.4]
  assign _T_12490 = 5'hd == _T_11317_24; // @[Mux.scala 46:19:@9630.4]
  assign _T_12491 = _T_12490 ? _T_10366_12 : _T_12489; // @[Mux.scala 46:16:@9631.4]
  assign _T_12492 = 5'hc == _T_11317_24; // @[Mux.scala 46:19:@9632.4]
  assign _T_12493 = _T_12492 ? _T_10366_11 : _T_12491; // @[Mux.scala 46:16:@9633.4]
  assign _T_12494 = 5'hb == _T_11317_24; // @[Mux.scala 46:19:@9634.4]
  assign _T_12495 = _T_12494 ? _T_10366_10 : _T_12493; // @[Mux.scala 46:16:@9635.4]
  assign _T_12496 = 5'ha == _T_11317_24; // @[Mux.scala 46:19:@9636.4]
  assign _T_12497 = _T_12496 ? _T_10366_9 : _T_12495; // @[Mux.scala 46:16:@9637.4]
  assign _T_12498 = 5'h9 == _T_11317_24; // @[Mux.scala 46:19:@9638.4]
  assign _T_12499 = _T_12498 ? _T_10366_8 : _T_12497; // @[Mux.scala 46:16:@9639.4]
  assign _T_12500 = 5'h8 == _T_11317_24; // @[Mux.scala 46:19:@9640.4]
  assign _T_12501 = _T_12500 ? _T_10366_7 : _T_12499; // @[Mux.scala 46:16:@9641.4]
  assign _T_12502 = 5'h7 == _T_11317_24; // @[Mux.scala 46:19:@9642.4]
  assign _T_12503 = _T_12502 ? _T_10366_6 : _T_12501; // @[Mux.scala 46:16:@9643.4]
  assign _T_12504 = 5'h6 == _T_11317_24; // @[Mux.scala 46:19:@9644.4]
  assign _T_12505 = _T_12504 ? _T_10366_5 : _T_12503; // @[Mux.scala 46:16:@9645.4]
  assign _T_12506 = 5'h5 == _T_11317_24; // @[Mux.scala 46:19:@9646.4]
  assign _T_12507 = _T_12506 ? _T_10366_4 : _T_12505; // @[Mux.scala 46:16:@9647.4]
  assign _T_12508 = 5'h4 == _T_11317_24; // @[Mux.scala 46:19:@9648.4]
  assign _T_12509 = _T_12508 ? _T_10366_3 : _T_12507; // @[Mux.scala 46:16:@9649.4]
  assign _T_12510 = 5'h3 == _T_11317_24; // @[Mux.scala 46:19:@9650.4]
  assign _T_12511 = _T_12510 ? _T_10366_2 : _T_12509; // @[Mux.scala 46:16:@9651.4]
  assign _T_12512 = 5'h2 == _T_11317_24; // @[Mux.scala 46:19:@9652.4]
  assign _T_12513 = _T_12512 ? _T_10366_1 : _T_12511; // @[Mux.scala 46:16:@9653.4]
  assign _T_12514 = 5'h1 == _T_11317_24; // @[Mux.scala 46:19:@9654.4]
  assign _T_12515 = _T_12514 ? _T_10366_0 : _T_12513; // @[Mux.scala 46:16:@9655.4]
  assign _T_12543 = 5'h1a == _T_11317_25; // @[Mux.scala 46:19:@9657.4]
  assign _T_12544 = _T_12543 ? _T_10366_25 : 8'h0; // @[Mux.scala 46:16:@9658.4]
  assign _T_12545 = 5'h19 == _T_11317_25; // @[Mux.scala 46:19:@9659.4]
  assign _T_12546 = _T_12545 ? _T_10366_24 : _T_12544; // @[Mux.scala 46:16:@9660.4]
  assign _T_12547 = 5'h18 == _T_11317_25; // @[Mux.scala 46:19:@9661.4]
  assign _T_12548 = _T_12547 ? _T_10366_23 : _T_12546; // @[Mux.scala 46:16:@9662.4]
  assign _T_12549 = 5'h17 == _T_11317_25; // @[Mux.scala 46:19:@9663.4]
  assign _T_12550 = _T_12549 ? _T_10366_22 : _T_12548; // @[Mux.scala 46:16:@9664.4]
  assign _T_12551 = 5'h16 == _T_11317_25; // @[Mux.scala 46:19:@9665.4]
  assign _T_12552 = _T_12551 ? _T_10366_21 : _T_12550; // @[Mux.scala 46:16:@9666.4]
  assign _T_12553 = 5'h15 == _T_11317_25; // @[Mux.scala 46:19:@9667.4]
  assign _T_12554 = _T_12553 ? _T_10366_20 : _T_12552; // @[Mux.scala 46:16:@9668.4]
  assign _T_12555 = 5'h14 == _T_11317_25; // @[Mux.scala 46:19:@9669.4]
  assign _T_12556 = _T_12555 ? _T_10366_19 : _T_12554; // @[Mux.scala 46:16:@9670.4]
  assign _T_12557 = 5'h13 == _T_11317_25; // @[Mux.scala 46:19:@9671.4]
  assign _T_12558 = _T_12557 ? _T_10366_18 : _T_12556; // @[Mux.scala 46:16:@9672.4]
  assign _T_12559 = 5'h12 == _T_11317_25; // @[Mux.scala 46:19:@9673.4]
  assign _T_12560 = _T_12559 ? _T_10366_17 : _T_12558; // @[Mux.scala 46:16:@9674.4]
  assign _T_12561 = 5'h11 == _T_11317_25; // @[Mux.scala 46:19:@9675.4]
  assign _T_12562 = _T_12561 ? _T_10366_16 : _T_12560; // @[Mux.scala 46:16:@9676.4]
  assign _T_12563 = 5'h10 == _T_11317_25; // @[Mux.scala 46:19:@9677.4]
  assign _T_12564 = _T_12563 ? _T_10366_15 : _T_12562; // @[Mux.scala 46:16:@9678.4]
  assign _T_12565 = 5'hf == _T_11317_25; // @[Mux.scala 46:19:@9679.4]
  assign _T_12566 = _T_12565 ? _T_10366_14 : _T_12564; // @[Mux.scala 46:16:@9680.4]
  assign _T_12567 = 5'he == _T_11317_25; // @[Mux.scala 46:19:@9681.4]
  assign _T_12568 = _T_12567 ? _T_10366_13 : _T_12566; // @[Mux.scala 46:16:@9682.4]
  assign _T_12569 = 5'hd == _T_11317_25; // @[Mux.scala 46:19:@9683.4]
  assign _T_12570 = _T_12569 ? _T_10366_12 : _T_12568; // @[Mux.scala 46:16:@9684.4]
  assign _T_12571 = 5'hc == _T_11317_25; // @[Mux.scala 46:19:@9685.4]
  assign _T_12572 = _T_12571 ? _T_10366_11 : _T_12570; // @[Mux.scala 46:16:@9686.4]
  assign _T_12573 = 5'hb == _T_11317_25; // @[Mux.scala 46:19:@9687.4]
  assign _T_12574 = _T_12573 ? _T_10366_10 : _T_12572; // @[Mux.scala 46:16:@9688.4]
  assign _T_12575 = 5'ha == _T_11317_25; // @[Mux.scala 46:19:@9689.4]
  assign _T_12576 = _T_12575 ? _T_10366_9 : _T_12574; // @[Mux.scala 46:16:@9690.4]
  assign _T_12577 = 5'h9 == _T_11317_25; // @[Mux.scala 46:19:@9691.4]
  assign _T_12578 = _T_12577 ? _T_10366_8 : _T_12576; // @[Mux.scala 46:16:@9692.4]
  assign _T_12579 = 5'h8 == _T_11317_25; // @[Mux.scala 46:19:@9693.4]
  assign _T_12580 = _T_12579 ? _T_10366_7 : _T_12578; // @[Mux.scala 46:16:@9694.4]
  assign _T_12581 = 5'h7 == _T_11317_25; // @[Mux.scala 46:19:@9695.4]
  assign _T_12582 = _T_12581 ? _T_10366_6 : _T_12580; // @[Mux.scala 46:16:@9696.4]
  assign _T_12583 = 5'h6 == _T_11317_25; // @[Mux.scala 46:19:@9697.4]
  assign _T_12584 = _T_12583 ? _T_10366_5 : _T_12582; // @[Mux.scala 46:16:@9698.4]
  assign _T_12585 = 5'h5 == _T_11317_25; // @[Mux.scala 46:19:@9699.4]
  assign _T_12586 = _T_12585 ? _T_10366_4 : _T_12584; // @[Mux.scala 46:16:@9700.4]
  assign _T_12587 = 5'h4 == _T_11317_25; // @[Mux.scala 46:19:@9701.4]
  assign _T_12588 = _T_12587 ? _T_10366_3 : _T_12586; // @[Mux.scala 46:16:@9702.4]
  assign _T_12589 = 5'h3 == _T_11317_25; // @[Mux.scala 46:19:@9703.4]
  assign _T_12590 = _T_12589 ? _T_10366_2 : _T_12588; // @[Mux.scala 46:16:@9704.4]
  assign _T_12591 = 5'h2 == _T_11317_25; // @[Mux.scala 46:19:@9705.4]
  assign _T_12592 = _T_12591 ? _T_10366_1 : _T_12590; // @[Mux.scala 46:16:@9706.4]
  assign _T_12593 = 5'h1 == _T_11317_25; // @[Mux.scala 46:19:@9707.4]
  assign _T_12594 = _T_12593 ? _T_10366_0 : _T_12592; // @[Mux.scala 46:16:@9708.4]
  assign _T_12623 = 5'h1b == _T_11317_26; // @[Mux.scala 46:19:@9710.4]
  assign _T_12624 = _T_12623 ? _T_10366_26 : 8'h0; // @[Mux.scala 46:16:@9711.4]
  assign _T_12625 = 5'h1a == _T_11317_26; // @[Mux.scala 46:19:@9712.4]
  assign _T_12626 = _T_12625 ? _T_10366_25 : _T_12624; // @[Mux.scala 46:16:@9713.4]
  assign _T_12627 = 5'h19 == _T_11317_26; // @[Mux.scala 46:19:@9714.4]
  assign _T_12628 = _T_12627 ? _T_10366_24 : _T_12626; // @[Mux.scala 46:16:@9715.4]
  assign _T_12629 = 5'h18 == _T_11317_26; // @[Mux.scala 46:19:@9716.4]
  assign _T_12630 = _T_12629 ? _T_10366_23 : _T_12628; // @[Mux.scala 46:16:@9717.4]
  assign _T_12631 = 5'h17 == _T_11317_26; // @[Mux.scala 46:19:@9718.4]
  assign _T_12632 = _T_12631 ? _T_10366_22 : _T_12630; // @[Mux.scala 46:16:@9719.4]
  assign _T_12633 = 5'h16 == _T_11317_26; // @[Mux.scala 46:19:@9720.4]
  assign _T_12634 = _T_12633 ? _T_10366_21 : _T_12632; // @[Mux.scala 46:16:@9721.4]
  assign _T_12635 = 5'h15 == _T_11317_26; // @[Mux.scala 46:19:@9722.4]
  assign _T_12636 = _T_12635 ? _T_10366_20 : _T_12634; // @[Mux.scala 46:16:@9723.4]
  assign _T_12637 = 5'h14 == _T_11317_26; // @[Mux.scala 46:19:@9724.4]
  assign _T_12638 = _T_12637 ? _T_10366_19 : _T_12636; // @[Mux.scala 46:16:@9725.4]
  assign _T_12639 = 5'h13 == _T_11317_26; // @[Mux.scala 46:19:@9726.4]
  assign _T_12640 = _T_12639 ? _T_10366_18 : _T_12638; // @[Mux.scala 46:16:@9727.4]
  assign _T_12641 = 5'h12 == _T_11317_26; // @[Mux.scala 46:19:@9728.4]
  assign _T_12642 = _T_12641 ? _T_10366_17 : _T_12640; // @[Mux.scala 46:16:@9729.4]
  assign _T_12643 = 5'h11 == _T_11317_26; // @[Mux.scala 46:19:@9730.4]
  assign _T_12644 = _T_12643 ? _T_10366_16 : _T_12642; // @[Mux.scala 46:16:@9731.4]
  assign _T_12645 = 5'h10 == _T_11317_26; // @[Mux.scala 46:19:@9732.4]
  assign _T_12646 = _T_12645 ? _T_10366_15 : _T_12644; // @[Mux.scala 46:16:@9733.4]
  assign _T_12647 = 5'hf == _T_11317_26; // @[Mux.scala 46:19:@9734.4]
  assign _T_12648 = _T_12647 ? _T_10366_14 : _T_12646; // @[Mux.scala 46:16:@9735.4]
  assign _T_12649 = 5'he == _T_11317_26; // @[Mux.scala 46:19:@9736.4]
  assign _T_12650 = _T_12649 ? _T_10366_13 : _T_12648; // @[Mux.scala 46:16:@9737.4]
  assign _T_12651 = 5'hd == _T_11317_26; // @[Mux.scala 46:19:@9738.4]
  assign _T_12652 = _T_12651 ? _T_10366_12 : _T_12650; // @[Mux.scala 46:16:@9739.4]
  assign _T_12653 = 5'hc == _T_11317_26; // @[Mux.scala 46:19:@9740.4]
  assign _T_12654 = _T_12653 ? _T_10366_11 : _T_12652; // @[Mux.scala 46:16:@9741.4]
  assign _T_12655 = 5'hb == _T_11317_26; // @[Mux.scala 46:19:@9742.4]
  assign _T_12656 = _T_12655 ? _T_10366_10 : _T_12654; // @[Mux.scala 46:16:@9743.4]
  assign _T_12657 = 5'ha == _T_11317_26; // @[Mux.scala 46:19:@9744.4]
  assign _T_12658 = _T_12657 ? _T_10366_9 : _T_12656; // @[Mux.scala 46:16:@9745.4]
  assign _T_12659 = 5'h9 == _T_11317_26; // @[Mux.scala 46:19:@9746.4]
  assign _T_12660 = _T_12659 ? _T_10366_8 : _T_12658; // @[Mux.scala 46:16:@9747.4]
  assign _T_12661 = 5'h8 == _T_11317_26; // @[Mux.scala 46:19:@9748.4]
  assign _T_12662 = _T_12661 ? _T_10366_7 : _T_12660; // @[Mux.scala 46:16:@9749.4]
  assign _T_12663 = 5'h7 == _T_11317_26; // @[Mux.scala 46:19:@9750.4]
  assign _T_12664 = _T_12663 ? _T_10366_6 : _T_12662; // @[Mux.scala 46:16:@9751.4]
  assign _T_12665 = 5'h6 == _T_11317_26; // @[Mux.scala 46:19:@9752.4]
  assign _T_12666 = _T_12665 ? _T_10366_5 : _T_12664; // @[Mux.scala 46:16:@9753.4]
  assign _T_12667 = 5'h5 == _T_11317_26; // @[Mux.scala 46:19:@9754.4]
  assign _T_12668 = _T_12667 ? _T_10366_4 : _T_12666; // @[Mux.scala 46:16:@9755.4]
  assign _T_12669 = 5'h4 == _T_11317_26; // @[Mux.scala 46:19:@9756.4]
  assign _T_12670 = _T_12669 ? _T_10366_3 : _T_12668; // @[Mux.scala 46:16:@9757.4]
  assign _T_12671 = 5'h3 == _T_11317_26; // @[Mux.scala 46:19:@9758.4]
  assign _T_12672 = _T_12671 ? _T_10366_2 : _T_12670; // @[Mux.scala 46:16:@9759.4]
  assign _T_12673 = 5'h2 == _T_11317_26; // @[Mux.scala 46:19:@9760.4]
  assign _T_12674 = _T_12673 ? _T_10366_1 : _T_12672; // @[Mux.scala 46:16:@9761.4]
  assign _T_12675 = 5'h1 == _T_11317_26; // @[Mux.scala 46:19:@9762.4]
  assign _T_12676 = _T_12675 ? _T_10366_0 : _T_12674; // @[Mux.scala 46:16:@9763.4]
  assign _T_12706 = 5'h1c == _T_11317_27; // @[Mux.scala 46:19:@9765.4]
  assign _T_12707 = _T_12706 ? _T_10366_27 : 8'h0; // @[Mux.scala 46:16:@9766.4]
  assign _T_12708 = 5'h1b == _T_11317_27; // @[Mux.scala 46:19:@9767.4]
  assign _T_12709 = _T_12708 ? _T_10366_26 : _T_12707; // @[Mux.scala 46:16:@9768.4]
  assign _T_12710 = 5'h1a == _T_11317_27; // @[Mux.scala 46:19:@9769.4]
  assign _T_12711 = _T_12710 ? _T_10366_25 : _T_12709; // @[Mux.scala 46:16:@9770.4]
  assign _T_12712 = 5'h19 == _T_11317_27; // @[Mux.scala 46:19:@9771.4]
  assign _T_12713 = _T_12712 ? _T_10366_24 : _T_12711; // @[Mux.scala 46:16:@9772.4]
  assign _T_12714 = 5'h18 == _T_11317_27; // @[Mux.scala 46:19:@9773.4]
  assign _T_12715 = _T_12714 ? _T_10366_23 : _T_12713; // @[Mux.scala 46:16:@9774.4]
  assign _T_12716 = 5'h17 == _T_11317_27; // @[Mux.scala 46:19:@9775.4]
  assign _T_12717 = _T_12716 ? _T_10366_22 : _T_12715; // @[Mux.scala 46:16:@9776.4]
  assign _T_12718 = 5'h16 == _T_11317_27; // @[Mux.scala 46:19:@9777.4]
  assign _T_12719 = _T_12718 ? _T_10366_21 : _T_12717; // @[Mux.scala 46:16:@9778.4]
  assign _T_12720 = 5'h15 == _T_11317_27; // @[Mux.scala 46:19:@9779.4]
  assign _T_12721 = _T_12720 ? _T_10366_20 : _T_12719; // @[Mux.scala 46:16:@9780.4]
  assign _T_12722 = 5'h14 == _T_11317_27; // @[Mux.scala 46:19:@9781.4]
  assign _T_12723 = _T_12722 ? _T_10366_19 : _T_12721; // @[Mux.scala 46:16:@9782.4]
  assign _T_12724 = 5'h13 == _T_11317_27; // @[Mux.scala 46:19:@9783.4]
  assign _T_12725 = _T_12724 ? _T_10366_18 : _T_12723; // @[Mux.scala 46:16:@9784.4]
  assign _T_12726 = 5'h12 == _T_11317_27; // @[Mux.scala 46:19:@9785.4]
  assign _T_12727 = _T_12726 ? _T_10366_17 : _T_12725; // @[Mux.scala 46:16:@9786.4]
  assign _T_12728 = 5'h11 == _T_11317_27; // @[Mux.scala 46:19:@9787.4]
  assign _T_12729 = _T_12728 ? _T_10366_16 : _T_12727; // @[Mux.scala 46:16:@9788.4]
  assign _T_12730 = 5'h10 == _T_11317_27; // @[Mux.scala 46:19:@9789.4]
  assign _T_12731 = _T_12730 ? _T_10366_15 : _T_12729; // @[Mux.scala 46:16:@9790.4]
  assign _T_12732 = 5'hf == _T_11317_27; // @[Mux.scala 46:19:@9791.4]
  assign _T_12733 = _T_12732 ? _T_10366_14 : _T_12731; // @[Mux.scala 46:16:@9792.4]
  assign _T_12734 = 5'he == _T_11317_27; // @[Mux.scala 46:19:@9793.4]
  assign _T_12735 = _T_12734 ? _T_10366_13 : _T_12733; // @[Mux.scala 46:16:@9794.4]
  assign _T_12736 = 5'hd == _T_11317_27; // @[Mux.scala 46:19:@9795.4]
  assign _T_12737 = _T_12736 ? _T_10366_12 : _T_12735; // @[Mux.scala 46:16:@9796.4]
  assign _T_12738 = 5'hc == _T_11317_27; // @[Mux.scala 46:19:@9797.4]
  assign _T_12739 = _T_12738 ? _T_10366_11 : _T_12737; // @[Mux.scala 46:16:@9798.4]
  assign _T_12740 = 5'hb == _T_11317_27; // @[Mux.scala 46:19:@9799.4]
  assign _T_12741 = _T_12740 ? _T_10366_10 : _T_12739; // @[Mux.scala 46:16:@9800.4]
  assign _T_12742 = 5'ha == _T_11317_27; // @[Mux.scala 46:19:@9801.4]
  assign _T_12743 = _T_12742 ? _T_10366_9 : _T_12741; // @[Mux.scala 46:16:@9802.4]
  assign _T_12744 = 5'h9 == _T_11317_27; // @[Mux.scala 46:19:@9803.4]
  assign _T_12745 = _T_12744 ? _T_10366_8 : _T_12743; // @[Mux.scala 46:16:@9804.4]
  assign _T_12746 = 5'h8 == _T_11317_27; // @[Mux.scala 46:19:@9805.4]
  assign _T_12747 = _T_12746 ? _T_10366_7 : _T_12745; // @[Mux.scala 46:16:@9806.4]
  assign _T_12748 = 5'h7 == _T_11317_27; // @[Mux.scala 46:19:@9807.4]
  assign _T_12749 = _T_12748 ? _T_10366_6 : _T_12747; // @[Mux.scala 46:16:@9808.4]
  assign _T_12750 = 5'h6 == _T_11317_27; // @[Mux.scala 46:19:@9809.4]
  assign _T_12751 = _T_12750 ? _T_10366_5 : _T_12749; // @[Mux.scala 46:16:@9810.4]
  assign _T_12752 = 5'h5 == _T_11317_27; // @[Mux.scala 46:19:@9811.4]
  assign _T_12753 = _T_12752 ? _T_10366_4 : _T_12751; // @[Mux.scala 46:16:@9812.4]
  assign _T_12754 = 5'h4 == _T_11317_27; // @[Mux.scala 46:19:@9813.4]
  assign _T_12755 = _T_12754 ? _T_10366_3 : _T_12753; // @[Mux.scala 46:16:@9814.4]
  assign _T_12756 = 5'h3 == _T_11317_27; // @[Mux.scala 46:19:@9815.4]
  assign _T_12757 = _T_12756 ? _T_10366_2 : _T_12755; // @[Mux.scala 46:16:@9816.4]
  assign _T_12758 = 5'h2 == _T_11317_27; // @[Mux.scala 46:19:@9817.4]
  assign _T_12759 = _T_12758 ? _T_10366_1 : _T_12757; // @[Mux.scala 46:16:@9818.4]
  assign _T_12760 = 5'h1 == _T_11317_27; // @[Mux.scala 46:19:@9819.4]
  assign _T_12761 = _T_12760 ? _T_10366_0 : _T_12759; // @[Mux.scala 46:16:@9820.4]
  assign _T_12792 = 5'h1d == _T_11317_28; // @[Mux.scala 46:19:@9822.4]
  assign _T_12793 = _T_12792 ? _T_10366_28 : 8'h0; // @[Mux.scala 46:16:@9823.4]
  assign _T_12794 = 5'h1c == _T_11317_28; // @[Mux.scala 46:19:@9824.4]
  assign _T_12795 = _T_12794 ? _T_10366_27 : _T_12793; // @[Mux.scala 46:16:@9825.4]
  assign _T_12796 = 5'h1b == _T_11317_28; // @[Mux.scala 46:19:@9826.4]
  assign _T_12797 = _T_12796 ? _T_10366_26 : _T_12795; // @[Mux.scala 46:16:@9827.4]
  assign _T_12798 = 5'h1a == _T_11317_28; // @[Mux.scala 46:19:@9828.4]
  assign _T_12799 = _T_12798 ? _T_10366_25 : _T_12797; // @[Mux.scala 46:16:@9829.4]
  assign _T_12800 = 5'h19 == _T_11317_28; // @[Mux.scala 46:19:@9830.4]
  assign _T_12801 = _T_12800 ? _T_10366_24 : _T_12799; // @[Mux.scala 46:16:@9831.4]
  assign _T_12802 = 5'h18 == _T_11317_28; // @[Mux.scala 46:19:@9832.4]
  assign _T_12803 = _T_12802 ? _T_10366_23 : _T_12801; // @[Mux.scala 46:16:@9833.4]
  assign _T_12804 = 5'h17 == _T_11317_28; // @[Mux.scala 46:19:@9834.4]
  assign _T_12805 = _T_12804 ? _T_10366_22 : _T_12803; // @[Mux.scala 46:16:@9835.4]
  assign _T_12806 = 5'h16 == _T_11317_28; // @[Mux.scala 46:19:@9836.4]
  assign _T_12807 = _T_12806 ? _T_10366_21 : _T_12805; // @[Mux.scala 46:16:@9837.4]
  assign _T_12808 = 5'h15 == _T_11317_28; // @[Mux.scala 46:19:@9838.4]
  assign _T_12809 = _T_12808 ? _T_10366_20 : _T_12807; // @[Mux.scala 46:16:@9839.4]
  assign _T_12810 = 5'h14 == _T_11317_28; // @[Mux.scala 46:19:@9840.4]
  assign _T_12811 = _T_12810 ? _T_10366_19 : _T_12809; // @[Mux.scala 46:16:@9841.4]
  assign _T_12812 = 5'h13 == _T_11317_28; // @[Mux.scala 46:19:@9842.4]
  assign _T_12813 = _T_12812 ? _T_10366_18 : _T_12811; // @[Mux.scala 46:16:@9843.4]
  assign _T_12814 = 5'h12 == _T_11317_28; // @[Mux.scala 46:19:@9844.4]
  assign _T_12815 = _T_12814 ? _T_10366_17 : _T_12813; // @[Mux.scala 46:16:@9845.4]
  assign _T_12816 = 5'h11 == _T_11317_28; // @[Mux.scala 46:19:@9846.4]
  assign _T_12817 = _T_12816 ? _T_10366_16 : _T_12815; // @[Mux.scala 46:16:@9847.4]
  assign _T_12818 = 5'h10 == _T_11317_28; // @[Mux.scala 46:19:@9848.4]
  assign _T_12819 = _T_12818 ? _T_10366_15 : _T_12817; // @[Mux.scala 46:16:@9849.4]
  assign _T_12820 = 5'hf == _T_11317_28; // @[Mux.scala 46:19:@9850.4]
  assign _T_12821 = _T_12820 ? _T_10366_14 : _T_12819; // @[Mux.scala 46:16:@9851.4]
  assign _T_12822 = 5'he == _T_11317_28; // @[Mux.scala 46:19:@9852.4]
  assign _T_12823 = _T_12822 ? _T_10366_13 : _T_12821; // @[Mux.scala 46:16:@9853.4]
  assign _T_12824 = 5'hd == _T_11317_28; // @[Mux.scala 46:19:@9854.4]
  assign _T_12825 = _T_12824 ? _T_10366_12 : _T_12823; // @[Mux.scala 46:16:@9855.4]
  assign _T_12826 = 5'hc == _T_11317_28; // @[Mux.scala 46:19:@9856.4]
  assign _T_12827 = _T_12826 ? _T_10366_11 : _T_12825; // @[Mux.scala 46:16:@9857.4]
  assign _T_12828 = 5'hb == _T_11317_28; // @[Mux.scala 46:19:@9858.4]
  assign _T_12829 = _T_12828 ? _T_10366_10 : _T_12827; // @[Mux.scala 46:16:@9859.4]
  assign _T_12830 = 5'ha == _T_11317_28; // @[Mux.scala 46:19:@9860.4]
  assign _T_12831 = _T_12830 ? _T_10366_9 : _T_12829; // @[Mux.scala 46:16:@9861.4]
  assign _T_12832 = 5'h9 == _T_11317_28; // @[Mux.scala 46:19:@9862.4]
  assign _T_12833 = _T_12832 ? _T_10366_8 : _T_12831; // @[Mux.scala 46:16:@9863.4]
  assign _T_12834 = 5'h8 == _T_11317_28; // @[Mux.scala 46:19:@9864.4]
  assign _T_12835 = _T_12834 ? _T_10366_7 : _T_12833; // @[Mux.scala 46:16:@9865.4]
  assign _T_12836 = 5'h7 == _T_11317_28; // @[Mux.scala 46:19:@9866.4]
  assign _T_12837 = _T_12836 ? _T_10366_6 : _T_12835; // @[Mux.scala 46:16:@9867.4]
  assign _T_12838 = 5'h6 == _T_11317_28; // @[Mux.scala 46:19:@9868.4]
  assign _T_12839 = _T_12838 ? _T_10366_5 : _T_12837; // @[Mux.scala 46:16:@9869.4]
  assign _T_12840 = 5'h5 == _T_11317_28; // @[Mux.scala 46:19:@9870.4]
  assign _T_12841 = _T_12840 ? _T_10366_4 : _T_12839; // @[Mux.scala 46:16:@9871.4]
  assign _T_12842 = 5'h4 == _T_11317_28; // @[Mux.scala 46:19:@9872.4]
  assign _T_12843 = _T_12842 ? _T_10366_3 : _T_12841; // @[Mux.scala 46:16:@9873.4]
  assign _T_12844 = 5'h3 == _T_11317_28; // @[Mux.scala 46:19:@9874.4]
  assign _T_12845 = _T_12844 ? _T_10366_2 : _T_12843; // @[Mux.scala 46:16:@9875.4]
  assign _T_12846 = 5'h2 == _T_11317_28; // @[Mux.scala 46:19:@9876.4]
  assign _T_12847 = _T_12846 ? _T_10366_1 : _T_12845; // @[Mux.scala 46:16:@9877.4]
  assign _T_12848 = 5'h1 == _T_11317_28; // @[Mux.scala 46:19:@9878.4]
  assign _T_12849 = _T_12848 ? _T_10366_0 : _T_12847; // @[Mux.scala 46:16:@9879.4]
  assign _T_12881 = 5'h1e == _T_11317_29; // @[Mux.scala 46:19:@9881.4]
  assign _T_12882 = _T_12881 ? _T_10366_29 : 8'h0; // @[Mux.scala 46:16:@9882.4]
  assign _T_12883 = 5'h1d == _T_11317_29; // @[Mux.scala 46:19:@9883.4]
  assign _T_12884 = _T_12883 ? _T_10366_28 : _T_12882; // @[Mux.scala 46:16:@9884.4]
  assign _T_12885 = 5'h1c == _T_11317_29; // @[Mux.scala 46:19:@9885.4]
  assign _T_12886 = _T_12885 ? _T_10366_27 : _T_12884; // @[Mux.scala 46:16:@9886.4]
  assign _T_12887 = 5'h1b == _T_11317_29; // @[Mux.scala 46:19:@9887.4]
  assign _T_12888 = _T_12887 ? _T_10366_26 : _T_12886; // @[Mux.scala 46:16:@9888.4]
  assign _T_12889 = 5'h1a == _T_11317_29; // @[Mux.scala 46:19:@9889.4]
  assign _T_12890 = _T_12889 ? _T_10366_25 : _T_12888; // @[Mux.scala 46:16:@9890.4]
  assign _T_12891 = 5'h19 == _T_11317_29; // @[Mux.scala 46:19:@9891.4]
  assign _T_12892 = _T_12891 ? _T_10366_24 : _T_12890; // @[Mux.scala 46:16:@9892.4]
  assign _T_12893 = 5'h18 == _T_11317_29; // @[Mux.scala 46:19:@9893.4]
  assign _T_12894 = _T_12893 ? _T_10366_23 : _T_12892; // @[Mux.scala 46:16:@9894.4]
  assign _T_12895 = 5'h17 == _T_11317_29; // @[Mux.scala 46:19:@9895.4]
  assign _T_12896 = _T_12895 ? _T_10366_22 : _T_12894; // @[Mux.scala 46:16:@9896.4]
  assign _T_12897 = 5'h16 == _T_11317_29; // @[Mux.scala 46:19:@9897.4]
  assign _T_12898 = _T_12897 ? _T_10366_21 : _T_12896; // @[Mux.scala 46:16:@9898.4]
  assign _T_12899 = 5'h15 == _T_11317_29; // @[Mux.scala 46:19:@9899.4]
  assign _T_12900 = _T_12899 ? _T_10366_20 : _T_12898; // @[Mux.scala 46:16:@9900.4]
  assign _T_12901 = 5'h14 == _T_11317_29; // @[Mux.scala 46:19:@9901.4]
  assign _T_12902 = _T_12901 ? _T_10366_19 : _T_12900; // @[Mux.scala 46:16:@9902.4]
  assign _T_12903 = 5'h13 == _T_11317_29; // @[Mux.scala 46:19:@9903.4]
  assign _T_12904 = _T_12903 ? _T_10366_18 : _T_12902; // @[Mux.scala 46:16:@9904.4]
  assign _T_12905 = 5'h12 == _T_11317_29; // @[Mux.scala 46:19:@9905.4]
  assign _T_12906 = _T_12905 ? _T_10366_17 : _T_12904; // @[Mux.scala 46:16:@9906.4]
  assign _T_12907 = 5'h11 == _T_11317_29; // @[Mux.scala 46:19:@9907.4]
  assign _T_12908 = _T_12907 ? _T_10366_16 : _T_12906; // @[Mux.scala 46:16:@9908.4]
  assign _T_12909 = 5'h10 == _T_11317_29; // @[Mux.scala 46:19:@9909.4]
  assign _T_12910 = _T_12909 ? _T_10366_15 : _T_12908; // @[Mux.scala 46:16:@9910.4]
  assign _T_12911 = 5'hf == _T_11317_29; // @[Mux.scala 46:19:@9911.4]
  assign _T_12912 = _T_12911 ? _T_10366_14 : _T_12910; // @[Mux.scala 46:16:@9912.4]
  assign _T_12913 = 5'he == _T_11317_29; // @[Mux.scala 46:19:@9913.4]
  assign _T_12914 = _T_12913 ? _T_10366_13 : _T_12912; // @[Mux.scala 46:16:@9914.4]
  assign _T_12915 = 5'hd == _T_11317_29; // @[Mux.scala 46:19:@9915.4]
  assign _T_12916 = _T_12915 ? _T_10366_12 : _T_12914; // @[Mux.scala 46:16:@9916.4]
  assign _T_12917 = 5'hc == _T_11317_29; // @[Mux.scala 46:19:@9917.4]
  assign _T_12918 = _T_12917 ? _T_10366_11 : _T_12916; // @[Mux.scala 46:16:@9918.4]
  assign _T_12919 = 5'hb == _T_11317_29; // @[Mux.scala 46:19:@9919.4]
  assign _T_12920 = _T_12919 ? _T_10366_10 : _T_12918; // @[Mux.scala 46:16:@9920.4]
  assign _T_12921 = 5'ha == _T_11317_29; // @[Mux.scala 46:19:@9921.4]
  assign _T_12922 = _T_12921 ? _T_10366_9 : _T_12920; // @[Mux.scala 46:16:@9922.4]
  assign _T_12923 = 5'h9 == _T_11317_29; // @[Mux.scala 46:19:@9923.4]
  assign _T_12924 = _T_12923 ? _T_10366_8 : _T_12922; // @[Mux.scala 46:16:@9924.4]
  assign _T_12925 = 5'h8 == _T_11317_29; // @[Mux.scala 46:19:@9925.4]
  assign _T_12926 = _T_12925 ? _T_10366_7 : _T_12924; // @[Mux.scala 46:16:@9926.4]
  assign _T_12927 = 5'h7 == _T_11317_29; // @[Mux.scala 46:19:@9927.4]
  assign _T_12928 = _T_12927 ? _T_10366_6 : _T_12926; // @[Mux.scala 46:16:@9928.4]
  assign _T_12929 = 5'h6 == _T_11317_29; // @[Mux.scala 46:19:@9929.4]
  assign _T_12930 = _T_12929 ? _T_10366_5 : _T_12928; // @[Mux.scala 46:16:@9930.4]
  assign _T_12931 = 5'h5 == _T_11317_29; // @[Mux.scala 46:19:@9931.4]
  assign _T_12932 = _T_12931 ? _T_10366_4 : _T_12930; // @[Mux.scala 46:16:@9932.4]
  assign _T_12933 = 5'h4 == _T_11317_29; // @[Mux.scala 46:19:@9933.4]
  assign _T_12934 = _T_12933 ? _T_10366_3 : _T_12932; // @[Mux.scala 46:16:@9934.4]
  assign _T_12935 = 5'h3 == _T_11317_29; // @[Mux.scala 46:19:@9935.4]
  assign _T_12936 = _T_12935 ? _T_10366_2 : _T_12934; // @[Mux.scala 46:16:@9936.4]
  assign _T_12937 = 5'h2 == _T_11317_29; // @[Mux.scala 46:19:@9937.4]
  assign _T_12938 = _T_12937 ? _T_10366_1 : _T_12936; // @[Mux.scala 46:16:@9938.4]
  assign _T_12939 = 5'h1 == _T_11317_29; // @[Mux.scala 46:19:@9939.4]
  assign _T_12940 = _T_12939 ? _T_10366_0 : _T_12938; // @[Mux.scala 46:16:@9940.4]
  assign _T_12973 = 5'h1f == _T_11317_30; // @[Mux.scala 46:19:@9942.4]
  assign _T_12974 = _T_12973 ? _T_10366_30 : 8'h0; // @[Mux.scala 46:16:@9943.4]
  assign _T_12975 = 5'h1e == _T_11317_30; // @[Mux.scala 46:19:@9944.4]
  assign _T_12976 = _T_12975 ? _T_10366_29 : _T_12974; // @[Mux.scala 46:16:@9945.4]
  assign _T_12977 = 5'h1d == _T_11317_30; // @[Mux.scala 46:19:@9946.4]
  assign _T_12978 = _T_12977 ? _T_10366_28 : _T_12976; // @[Mux.scala 46:16:@9947.4]
  assign _T_12979 = 5'h1c == _T_11317_30; // @[Mux.scala 46:19:@9948.4]
  assign _T_12980 = _T_12979 ? _T_10366_27 : _T_12978; // @[Mux.scala 46:16:@9949.4]
  assign _T_12981 = 5'h1b == _T_11317_30; // @[Mux.scala 46:19:@9950.4]
  assign _T_12982 = _T_12981 ? _T_10366_26 : _T_12980; // @[Mux.scala 46:16:@9951.4]
  assign _T_12983 = 5'h1a == _T_11317_30; // @[Mux.scala 46:19:@9952.4]
  assign _T_12984 = _T_12983 ? _T_10366_25 : _T_12982; // @[Mux.scala 46:16:@9953.4]
  assign _T_12985 = 5'h19 == _T_11317_30; // @[Mux.scala 46:19:@9954.4]
  assign _T_12986 = _T_12985 ? _T_10366_24 : _T_12984; // @[Mux.scala 46:16:@9955.4]
  assign _T_12987 = 5'h18 == _T_11317_30; // @[Mux.scala 46:19:@9956.4]
  assign _T_12988 = _T_12987 ? _T_10366_23 : _T_12986; // @[Mux.scala 46:16:@9957.4]
  assign _T_12989 = 5'h17 == _T_11317_30; // @[Mux.scala 46:19:@9958.4]
  assign _T_12990 = _T_12989 ? _T_10366_22 : _T_12988; // @[Mux.scala 46:16:@9959.4]
  assign _T_12991 = 5'h16 == _T_11317_30; // @[Mux.scala 46:19:@9960.4]
  assign _T_12992 = _T_12991 ? _T_10366_21 : _T_12990; // @[Mux.scala 46:16:@9961.4]
  assign _T_12993 = 5'h15 == _T_11317_30; // @[Mux.scala 46:19:@9962.4]
  assign _T_12994 = _T_12993 ? _T_10366_20 : _T_12992; // @[Mux.scala 46:16:@9963.4]
  assign _T_12995 = 5'h14 == _T_11317_30; // @[Mux.scala 46:19:@9964.4]
  assign _T_12996 = _T_12995 ? _T_10366_19 : _T_12994; // @[Mux.scala 46:16:@9965.4]
  assign _T_12997 = 5'h13 == _T_11317_30; // @[Mux.scala 46:19:@9966.4]
  assign _T_12998 = _T_12997 ? _T_10366_18 : _T_12996; // @[Mux.scala 46:16:@9967.4]
  assign _T_12999 = 5'h12 == _T_11317_30; // @[Mux.scala 46:19:@9968.4]
  assign _T_13000 = _T_12999 ? _T_10366_17 : _T_12998; // @[Mux.scala 46:16:@9969.4]
  assign _T_13001 = 5'h11 == _T_11317_30; // @[Mux.scala 46:19:@9970.4]
  assign _T_13002 = _T_13001 ? _T_10366_16 : _T_13000; // @[Mux.scala 46:16:@9971.4]
  assign _T_13003 = 5'h10 == _T_11317_30; // @[Mux.scala 46:19:@9972.4]
  assign _T_13004 = _T_13003 ? _T_10366_15 : _T_13002; // @[Mux.scala 46:16:@9973.4]
  assign _T_13005 = 5'hf == _T_11317_30; // @[Mux.scala 46:19:@9974.4]
  assign _T_13006 = _T_13005 ? _T_10366_14 : _T_13004; // @[Mux.scala 46:16:@9975.4]
  assign _T_13007 = 5'he == _T_11317_30; // @[Mux.scala 46:19:@9976.4]
  assign _T_13008 = _T_13007 ? _T_10366_13 : _T_13006; // @[Mux.scala 46:16:@9977.4]
  assign _T_13009 = 5'hd == _T_11317_30; // @[Mux.scala 46:19:@9978.4]
  assign _T_13010 = _T_13009 ? _T_10366_12 : _T_13008; // @[Mux.scala 46:16:@9979.4]
  assign _T_13011 = 5'hc == _T_11317_30; // @[Mux.scala 46:19:@9980.4]
  assign _T_13012 = _T_13011 ? _T_10366_11 : _T_13010; // @[Mux.scala 46:16:@9981.4]
  assign _T_13013 = 5'hb == _T_11317_30; // @[Mux.scala 46:19:@9982.4]
  assign _T_13014 = _T_13013 ? _T_10366_10 : _T_13012; // @[Mux.scala 46:16:@9983.4]
  assign _T_13015 = 5'ha == _T_11317_30; // @[Mux.scala 46:19:@9984.4]
  assign _T_13016 = _T_13015 ? _T_10366_9 : _T_13014; // @[Mux.scala 46:16:@9985.4]
  assign _T_13017 = 5'h9 == _T_11317_30; // @[Mux.scala 46:19:@9986.4]
  assign _T_13018 = _T_13017 ? _T_10366_8 : _T_13016; // @[Mux.scala 46:16:@9987.4]
  assign _T_13019 = 5'h8 == _T_11317_30; // @[Mux.scala 46:19:@9988.4]
  assign _T_13020 = _T_13019 ? _T_10366_7 : _T_13018; // @[Mux.scala 46:16:@9989.4]
  assign _T_13021 = 5'h7 == _T_11317_30; // @[Mux.scala 46:19:@9990.4]
  assign _T_13022 = _T_13021 ? _T_10366_6 : _T_13020; // @[Mux.scala 46:16:@9991.4]
  assign _T_13023 = 5'h6 == _T_11317_30; // @[Mux.scala 46:19:@9992.4]
  assign _T_13024 = _T_13023 ? _T_10366_5 : _T_13022; // @[Mux.scala 46:16:@9993.4]
  assign _T_13025 = 5'h5 == _T_11317_30; // @[Mux.scala 46:19:@9994.4]
  assign _T_13026 = _T_13025 ? _T_10366_4 : _T_13024; // @[Mux.scala 46:16:@9995.4]
  assign _T_13027 = 5'h4 == _T_11317_30; // @[Mux.scala 46:19:@9996.4]
  assign _T_13028 = _T_13027 ? _T_10366_3 : _T_13026; // @[Mux.scala 46:16:@9997.4]
  assign _T_13029 = 5'h3 == _T_11317_30; // @[Mux.scala 46:19:@9998.4]
  assign _T_13030 = _T_13029 ? _T_10366_2 : _T_13028; // @[Mux.scala 46:16:@9999.4]
  assign _T_13031 = 5'h2 == _T_11317_30; // @[Mux.scala 46:19:@10000.4]
  assign _T_13032 = _T_13031 ? _T_10366_1 : _T_13030; // @[Mux.scala 46:16:@10001.4]
  assign _T_13033 = 5'h1 == _T_11317_30; // @[Mux.scala 46:19:@10002.4]
  assign _T_13034 = _T_13033 ? _T_10366_0 : _T_13032; // @[Mux.scala 46:16:@10003.4]
  assign _T_13068 = 6'h20 == _T_11317_31; // @[Mux.scala 46:19:@10005.4]
  assign _T_13069 = _T_13068 ? _T_10366_31 : 8'h0; // @[Mux.scala 46:16:@10006.4]
  assign _T_13070 = 6'h1f == _T_11317_31; // @[Mux.scala 46:19:@10007.4]
  assign _T_13071 = _T_13070 ? _T_10366_30 : _T_13069; // @[Mux.scala 46:16:@10008.4]
  assign _T_13072 = 6'h1e == _T_11317_31; // @[Mux.scala 46:19:@10009.4]
  assign _T_13073 = _T_13072 ? _T_10366_29 : _T_13071; // @[Mux.scala 46:16:@10010.4]
  assign _T_13074 = 6'h1d == _T_11317_31; // @[Mux.scala 46:19:@10011.4]
  assign _T_13075 = _T_13074 ? _T_10366_28 : _T_13073; // @[Mux.scala 46:16:@10012.4]
  assign _T_13076 = 6'h1c == _T_11317_31; // @[Mux.scala 46:19:@10013.4]
  assign _T_13077 = _T_13076 ? _T_10366_27 : _T_13075; // @[Mux.scala 46:16:@10014.4]
  assign _T_13078 = 6'h1b == _T_11317_31; // @[Mux.scala 46:19:@10015.4]
  assign _T_13079 = _T_13078 ? _T_10366_26 : _T_13077; // @[Mux.scala 46:16:@10016.4]
  assign _T_13080 = 6'h1a == _T_11317_31; // @[Mux.scala 46:19:@10017.4]
  assign _T_13081 = _T_13080 ? _T_10366_25 : _T_13079; // @[Mux.scala 46:16:@10018.4]
  assign _T_13082 = 6'h19 == _T_11317_31; // @[Mux.scala 46:19:@10019.4]
  assign _T_13083 = _T_13082 ? _T_10366_24 : _T_13081; // @[Mux.scala 46:16:@10020.4]
  assign _T_13084 = 6'h18 == _T_11317_31; // @[Mux.scala 46:19:@10021.4]
  assign _T_13085 = _T_13084 ? _T_10366_23 : _T_13083; // @[Mux.scala 46:16:@10022.4]
  assign _T_13086 = 6'h17 == _T_11317_31; // @[Mux.scala 46:19:@10023.4]
  assign _T_13087 = _T_13086 ? _T_10366_22 : _T_13085; // @[Mux.scala 46:16:@10024.4]
  assign _T_13088 = 6'h16 == _T_11317_31; // @[Mux.scala 46:19:@10025.4]
  assign _T_13089 = _T_13088 ? _T_10366_21 : _T_13087; // @[Mux.scala 46:16:@10026.4]
  assign _T_13090 = 6'h15 == _T_11317_31; // @[Mux.scala 46:19:@10027.4]
  assign _T_13091 = _T_13090 ? _T_10366_20 : _T_13089; // @[Mux.scala 46:16:@10028.4]
  assign _T_13092 = 6'h14 == _T_11317_31; // @[Mux.scala 46:19:@10029.4]
  assign _T_13093 = _T_13092 ? _T_10366_19 : _T_13091; // @[Mux.scala 46:16:@10030.4]
  assign _T_13094 = 6'h13 == _T_11317_31; // @[Mux.scala 46:19:@10031.4]
  assign _T_13095 = _T_13094 ? _T_10366_18 : _T_13093; // @[Mux.scala 46:16:@10032.4]
  assign _T_13096 = 6'h12 == _T_11317_31; // @[Mux.scala 46:19:@10033.4]
  assign _T_13097 = _T_13096 ? _T_10366_17 : _T_13095; // @[Mux.scala 46:16:@10034.4]
  assign _T_13098 = 6'h11 == _T_11317_31; // @[Mux.scala 46:19:@10035.4]
  assign _T_13099 = _T_13098 ? _T_10366_16 : _T_13097; // @[Mux.scala 46:16:@10036.4]
  assign _T_13100 = 6'h10 == _T_11317_31; // @[Mux.scala 46:19:@10037.4]
  assign _T_13101 = _T_13100 ? _T_10366_15 : _T_13099; // @[Mux.scala 46:16:@10038.4]
  assign _T_13102 = 6'hf == _T_11317_31; // @[Mux.scala 46:19:@10039.4]
  assign _T_13103 = _T_13102 ? _T_10366_14 : _T_13101; // @[Mux.scala 46:16:@10040.4]
  assign _T_13104 = 6'he == _T_11317_31; // @[Mux.scala 46:19:@10041.4]
  assign _T_13105 = _T_13104 ? _T_10366_13 : _T_13103; // @[Mux.scala 46:16:@10042.4]
  assign _T_13106 = 6'hd == _T_11317_31; // @[Mux.scala 46:19:@10043.4]
  assign _T_13107 = _T_13106 ? _T_10366_12 : _T_13105; // @[Mux.scala 46:16:@10044.4]
  assign _T_13108 = 6'hc == _T_11317_31; // @[Mux.scala 46:19:@10045.4]
  assign _T_13109 = _T_13108 ? _T_10366_11 : _T_13107; // @[Mux.scala 46:16:@10046.4]
  assign _T_13110 = 6'hb == _T_11317_31; // @[Mux.scala 46:19:@10047.4]
  assign _T_13111 = _T_13110 ? _T_10366_10 : _T_13109; // @[Mux.scala 46:16:@10048.4]
  assign _T_13112 = 6'ha == _T_11317_31; // @[Mux.scala 46:19:@10049.4]
  assign _T_13113 = _T_13112 ? _T_10366_9 : _T_13111; // @[Mux.scala 46:16:@10050.4]
  assign _T_13114 = 6'h9 == _T_11317_31; // @[Mux.scala 46:19:@10051.4]
  assign _T_13115 = _T_13114 ? _T_10366_8 : _T_13113; // @[Mux.scala 46:16:@10052.4]
  assign _T_13116 = 6'h8 == _T_11317_31; // @[Mux.scala 46:19:@10053.4]
  assign _T_13117 = _T_13116 ? _T_10366_7 : _T_13115; // @[Mux.scala 46:16:@10054.4]
  assign _T_13118 = 6'h7 == _T_11317_31; // @[Mux.scala 46:19:@10055.4]
  assign _T_13119 = _T_13118 ? _T_10366_6 : _T_13117; // @[Mux.scala 46:16:@10056.4]
  assign _T_13120 = 6'h6 == _T_11317_31; // @[Mux.scala 46:19:@10057.4]
  assign _T_13121 = _T_13120 ? _T_10366_5 : _T_13119; // @[Mux.scala 46:16:@10058.4]
  assign _T_13122 = 6'h5 == _T_11317_31; // @[Mux.scala 46:19:@10059.4]
  assign _T_13123 = _T_13122 ? _T_10366_4 : _T_13121; // @[Mux.scala 46:16:@10060.4]
  assign _T_13124 = 6'h4 == _T_11317_31; // @[Mux.scala 46:19:@10061.4]
  assign _T_13125 = _T_13124 ? _T_10366_3 : _T_13123; // @[Mux.scala 46:16:@10062.4]
  assign _T_13126 = 6'h3 == _T_11317_31; // @[Mux.scala 46:19:@10063.4]
  assign _T_13127 = _T_13126 ? _T_10366_2 : _T_13125; // @[Mux.scala 46:16:@10064.4]
  assign _T_13128 = 6'h2 == _T_11317_31; // @[Mux.scala 46:19:@10065.4]
  assign _T_13129 = _T_13128 ? _T_10366_1 : _T_13127; // @[Mux.scala 46:16:@10066.4]
  assign _T_13130 = 6'h1 == _T_11317_31; // @[Mux.scala 46:19:@10067.4]
  assign _T_13131 = _T_13130 ? _T_10366_0 : _T_13129; // @[Mux.scala 46:16:@10068.4]
  assign _T_13166 = 6'h21 == _T_11317_32; // @[Mux.scala 46:19:@10070.4]
  assign _T_13167 = _T_13166 ? _T_10366_32 : 8'h0; // @[Mux.scala 46:16:@10071.4]
  assign _T_13168 = 6'h20 == _T_11317_32; // @[Mux.scala 46:19:@10072.4]
  assign _T_13169 = _T_13168 ? _T_10366_31 : _T_13167; // @[Mux.scala 46:16:@10073.4]
  assign _T_13170 = 6'h1f == _T_11317_32; // @[Mux.scala 46:19:@10074.4]
  assign _T_13171 = _T_13170 ? _T_10366_30 : _T_13169; // @[Mux.scala 46:16:@10075.4]
  assign _T_13172 = 6'h1e == _T_11317_32; // @[Mux.scala 46:19:@10076.4]
  assign _T_13173 = _T_13172 ? _T_10366_29 : _T_13171; // @[Mux.scala 46:16:@10077.4]
  assign _T_13174 = 6'h1d == _T_11317_32; // @[Mux.scala 46:19:@10078.4]
  assign _T_13175 = _T_13174 ? _T_10366_28 : _T_13173; // @[Mux.scala 46:16:@10079.4]
  assign _T_13176 = 6'h1c == _T_11317_32; // @[Mux.scala 46:19:@10080.4]
  assign _T_13177 = _T_13176 ? _T_10366_27 : _T_13175; // @[Mux.scala 46:16:@10081.4]
  assign _T_13178 = 6'h1b == _T_11317_32; // @[Mux.scala 46:19:@10082.4]
  assign _T_13179 = _T_13178 ? _T_10366_26 : _T_13177; // @[Mux.scala 46:16:@10083.4]
  assign _T_13180 = 6'h1a == _T_11317_32; // @[Mux.scala 46:19:@10084.4]
  assign _T_13181 = _T_13180 ? _T_10366_25 : _T_13179; // @[Mux.scala 46:16:@10085.4]
  assign _T_13182 = 6'h19 == _T_11317_32; // @[Mux.scala 46:19:@10086.4]
  assign _T_13183 = _T_13182 ? _T_10366_24 : _T_13181; // @[Mux.scala 46:16:@10087.4]
  assign _T_13184 = 6'h18 == _T_11317_32; // @[Mux.scala 46:19:@10088.4]
  assign _T_13185 = _T_13184 ? _T_10366_23 : _T_13183; // @[Mux.scala 46:16:@10089.4]
  assign _T_13186 = 6'h17 == _T_11317_32; // @[Mux.scala 46:19:@10090.4]
  assign _T_13187 = _T_13186 ? _T_10366_22 : _T_13185; // @[Mux.scala 46:16:@10091.4]
  assign _T_13188 = 6'h16 == _T_11317_32; // @[Mux.scala 46:19:@10092.4]
  assign _T_13189 = _T_13188 ? _T_10366_21 : _T_13187; // @[Mux.scala 46:16:@10093.4]
  assign _T_13190 = 6'h15 == _T_11317_32; // @[Mux.scala 46:19:@10094.4]
  assign _T_13191 = _T_13190 ? _T_10366_20 : _T_13189; // @[Mux.scala 46:16:@10095.4]
  assign _T_13192 = 6'h14 == _T_11317_32; // @[Mux.scala 46:19:@10096.4]
  assign _T_13193 = _T_13192 ? _T_10366_19 : _T_13191; // @[Mux.scala 46:16:@10097.4]
  assign _T_13194 = 6'h13 == _T_11317_32; // @[Mux.scala 46:19:@10098.4]
  assign _T_13195 = _T_13194 ? _T_10366_18 : _T_13193; // @[Mux.scala 46:16:@10099.4]
  assign _T_13196 = 6'h12 == _T_11317_32; // @[Mux.scala 46:19:@10100.4]
  assign _T_13197 = _T_13196 ? _T_10366_17 : _T_13195; // @[Mux.scala 46:16:@10101.4]
  assign _T_13198 = 6'h11 == _T_11317_32; // @[Mux.scala 46:19:@10102.4]
  assign _T_13199 = _T_13198 ? _T_10366_16 : _T_13197; // @[Mux.scala 46:16:@10103.4]
  assign _T_13200 = 6'h10 == _T_11317_32; // @[Mux.scala 46:19:@10104.4]
  assign _T_13201 = _T_13200 ? _T_10366_15 : _T_13199; // @[Mux.scala 46:16:@10105.4]
  assign _T_13202 = 6'hf == _T_11317_32; // @[Mux.scala 46:19:@10106.4]
  assign _T_13203 = _T_13202 ? _T_10366_14 : _T_13201; // @[Mux.scala 46:16:@10107.4]
  assign _T_13204 = 6'he == _T_11317_32; // @[Mux.scala 46:19:@10108.4]
  assign _T_13205 = _T_13204 ? _T_10366_13 : _T_13203; // @[Mux.scala 46:16:@10109.4]
  assign _T_13206 = 6'hd == _T_11317_32; // @[Mux.scala 46:19:@10110.4]
  assign _T_13207 = _T_13206 ? _T_10366_12 : _T_13205; // @[Mux.scala 46:16:@10111.4]
  assign _T_13208 = 6'hc == _T_11317_32; // @[Mux.scala 46:19:@10112.4]
  assign _T_13209 = _T_13208 ? _T_10366_11 : _T_13207; // @[Mux.scala 46:16:@10113.4]
  assign _T_13210 = 6'hb == _T_11317_32; // @[Mux.scala 46:19:@10114.4]
  assign _T_13211 = _T_13210 ? _T_10366_10 : _T_13209; // @[Mux.scala 46:16:@10115.4]
  assign _T_13212 = 6'ha == _T_11317_32; // @[Mux.scala 46:19:@10116.4]
  assign _T_13213 = _T_13212 ? _T_10366_9 : _T_13211; // @[Mux.scala 46:16:@10117.4]
  assign _T_13214 = 6'h9 == _T_11317_32; // @[Mux.scala 46:19:@10118.4]
  assign _T_13215 = _T_13214 ? _T_10366_8 : _T_13213; // @[Mux.scala 46:16:@10119.4]
  assign _T_13216 = 6'h8 == _T_11317_32; // @[Mux.scala 46:19:@10120.4]
  assign _T_13217 = _T_13216 ? _T_10366_7 : _T_13215; // @[Mux.scala 46:16:@10121.4]
  assign _T_13218 = 6'h7 == _T_11317_32; // @[Mux.scala 46:19:@10122.4]
  assign _T_13219 = _T_13218 ? _T_10366_6 : _T_13217; // @[Mux.scala 46:16:@10123.4]
  assign _T_13220 = 6'h6 == _T_11317_32; // @[Mux.scala 46:19:@10124.4]
  assign _T_13221 = _T_13220 ? _T_10366_5 : _T_13219; // @[Mux.scala 46:16:@10125.4]
  assign _T_13222 = 6'h5 == _T_11317_32; // @[Mux.scala 46:19:@10126.4]
  assign _T_13223 = _T_13222 ? _T_10366_4 : _T_13221; // @[Mux.scala 46:16:@10127.4]
  assign _T_13224 = 6'h4 == _T_11317_32; // @[Mux.scala 46:19:@10128.4]
  assign _T_13225 = _T_13224 ? _T_10366_3 : _T_13223; // @[Mux.scala 46:16:@10129.4]
  assign _T_13226 = 6'h3 == _T_11317_32; // @[Mux.scala 46:19:@10130.4]
  assign _T_13227 = _T_13226 ? _T_10366_2 : _T_13225; // @[Mux.scala 46:16:@10131.4]
  assign _T_13228 = 6'h2 == _T_11317_32; // @[Mux.scala 46:19:@10132.4]
  assign _T_13229 = _T_13228 ? _T_10366_1 : _T_13227; // @[Mux.scala 46:16:@10133.4]
  assign _T_13230 = 6'h1 == _T_11317_32; // @[Mux.scala 46:19:@10134.4]
  assign _T_13231 = _T_13230 ? _T_10366_0 : _T_13229; // @[Mux.scala 46:16:@10135.4]
  assign _T_13267 = 6'h22 == _T_11317_33; // @[Mux.scala 46:19:@10137.4]
  assign _T_13268 = _T_13267 ? _T_10366_33 : 8'h0; // @[Mux.scala 46:16:@10138.4]
  assign _T_13269 = 6'h21 == _T_11317_33; // @[Mux.scala 46:19:@10139.4]
  assign _T_13270 = _T_13269 ? _T_10366_32 : _T_13268; // @[Mux.scala 46:16:@10140.4]
  assign _T_13271 = 6'h20 == _T_11317_33; // @[Mux.scala 46:19:@10141.4]
  assign _T_13272 = _T_13271 ? _T_10366_31 : _T_13270; // @[Mux.scala 46:16:@10142.4]
  assign _T_13273 = 6'h1f == _T_11317_33; // @[Mux.scala 46:19:@10143.4]
  assign _T_13274 = _T_13273 ? _T_10366_30 : _T_13272; // @[Mux.scala 46:16:@10144.4]
  assign _T_13275 = 6'h1e == _T_11317_33; // @[Mux.scala 46:19:@10145.4]
  assign _T_13276 = _T_13275 ? _T_10366_29 : _T_13274; // @[Mux.scala 46:16:@10146.4]
  assign _T_13277 = 6'h1d == _T_11317_33; // @[Mux.scala 46:19:@10147.4]
  assign _T_13278 = _T_13277 ? _T_10366_28 : _T_13276; // @[Mux.scala 46:16:@10148.4]
  assign _T_13279 = 6'h1c == _T_11317_33; // @[Mux.scala 46:19:@10149.4]
  assign _T_13280 = _T_13279 ? _T_10366_27 : _T_13278; // @[Mux.scala 46:16:@10150.4]
  assign _T_13281 = 6'h1b == _T_11317_33; // @[Mux.scala 46:19:@10151.4]
  assign _T_13282 = _T_13281 ? _T_10366_26 : _T_13280; // @[Mux.scala 46:16:@10152.4]
  assign _T_13283 = 6'h1a == _T_11317_33; // @[Mux.scala 46:19:@10153.4]
  assign _T_13284 = _T_13283 ? _T_10366_25 : _T_13282; // @[Mux.scala 46:16:@10154.4]
  assign _T_13285 = 6'h19 == _T_11317_33; // @[Mux.scala 46:19:@10155.4]
  assign _T_13286 = _T_13285 ? _T_10366_24 : _T_13284; // @[Mux.scala 46:16:@10156.4]
  assign _T_13287 = 6'h18 == _T_11317_33; // @[Mux.scala 46:19:@10157.4]
  assign _T_13288 = _T_13287 ? _T_10366_23 : _T_13286; // @[Mux.scala 46:16:@10158.4]
  assign _T_13289 = 6'h17 == _T_11317_33; // @[Mux.scala 46:19:@10159.4]
  assign _T_13290 = _T_13289 ? _T_10366_22 : _T_13288; // @[Mux.scala 46:16:@10160.4]
  assign _T_13291 = 6'h16 == _T_11317_33; // @[Mux.scala 46:19:@10161.4]
  assign _T_13292 = _T_13291 ? _T_10366_21 : _T_13290; // @[Mux.scala 46:16:@10162.4]
  assign _T_13293 = 6'h15 == _T_11317_33; // @[Mux.scala 46:19:@10163.4]
  assign _T_13294 = _T_13293 ? _T_10366_20 : _T_13292; // @[Mux.scala 46:16:@10164.4]
  assign _T_13295 = 6'h14 == _T_11317_33; // @[Mux.scala 46:19:@10165.4]
  assign _T_13296 = _T_13295 ? _T_10366_19 : _T_13294; // @[Mux.scala 46:16:@10166.4]
  assign _T_13297 = 6'h13 == _T_11317_33; // @[Mux.scala 46:19:@10167.4]
  assign _T_13298 = _T_13297 ? _T_10366_18 : _T_13296; // @[Mux.scala 46:16:@10168.4]
  assign _T_13299 = 6'h12 == _T_11317_33; // @[Mux.scala 46:19:@10169.4]
  assign _T_13300 = _T_13299 ? _T_10366_17 : _T_13298; // @[Mux.scala 46:16:@10170.4]
  assign _T_13301 = 6'h11 == _T_11317_33; // @[Mux.scala 46:19:@10171.4]
  assign _T_13302 = _T_13301 ? _T_10366_16 : _T_13300; // @[Mux.scala 46:16:@10172.4]
  assign _T_13303 = 6'h10 == _T_11317_33; // @[Mux.scala 46:19:@10173.4]
  assign _T_13304 = _T_13303 ? _T_10366_15 : _T_13302; // @[Mux.scala 46:16:@10174.4]
  assign _T_13305 = 6'hf == _T_11317_33; // @[Mux.scala 46:19:@10175.4]
  assign _T_13306 = _T_13305 ? _T_10366_14 : _T_13304; // @[Mux.scala 46:16:@10176.4]
  assign _T_13307 = 6'he == _T_11317_33; // @[Mux.scala 46:19:@10177.4]
  assign _T_13308 = _T_13307 ? _T_10366_13 : _T_13306; // @[Mux.scala 46:16:@10178.4]
  assign _T_13309 = 6'hd == _T_11317_33; // @[Mux.scala 46:19:@10179.4]
  assign _T_13310 = _T_13309 ? _T_10366_12 : _T_13308; // @[Mux.scala 46:16:@10180.4]
  assign _T_13311 = 6'hc == _T_11317_33; // @[Mux.scala 46:19:@10181.4]
  assign _T_13312 = _T_13311 ? _T_10366_11 : _T_13310; // @[Mux.scala 46:16:@10182.4]
  assign _T_13313 = 6'hb == _T_11317_33; // @[Mux.scala 46:19:@10183.4]
  assign _T_13314 = _T_13313 ? _T_10366_10 : _T_13312; // @[Mux.scala 46:16:@10184.4]
  assign _T_13315 = 6'ha == _T_11317_33; // @[Mux.scala 46:19:@10185.4]
  assign _T_13316 = _T_13315 ? _T_10366_9 : _T_13314; // @[Mux.scala 46:16:@10186.4]
  assign _T_13317 = 6'h9 == _T_11317_33; // @[Mux.scala 46:19:@10187.4]
  assign _T_13318 = _T_13317 ? _T_10366_8 : _T_13316; // @[Mux.scala 46:16:@10188.4]
  assign _T_13319 = 6'h8 == _T_11317_33; // @[Mux.scala 46:19:@10189.4]
  assign _T_13320 = _T_13319 ? _T_10366_7 : _T_13318; // @[Mux.scala 46:16:@10190.4]
  assign _T_13321 = 6'h7 == _T_11317_33; // @[Mux.scala 46:19:@10191.4]
  assign _T_13322 = _T_13321 ? _T_10366_6 : _T_13320; // @[Mux.scala 46:16:@10192.4]
  assign _T_13323 = 6'h6 == _T_11317_33; // @[Mux.scala 46:19:@10193.4]
  assign _T_13324 = _T_13323 ? _T_10366_5 : _T_13322; // @[Mux.scala 46:16:@10194.4]
  assign _T_13325 = 6'h5 == _T_11317_33; // @[Mux.scala 46:19:@10195.4]
  assign _T_13326 = _T_13325 ? _T_10366_4 : _T_13324; // @[Mux.scala 46:16:@10196.4]
  assign _T_13327 = 6'h4 == _T_11317_33; // @[Mux.scala 46:19:@10197.4]
  assign _T_13328 = _T_13327 ? _T_10366_3 : _T_13326; // @[Mux.scala 46:16:@10198.4]
  assign _T_13329 = 6'h3 == _T_11317_33; // @[Mux.scala 46:19:@10199.4]
  assign _T_13330 = _T_13329 ? _T_10366_2 : _T_13328; // @[Mux.scala 46:16:@10200.4]
  assign _T_13331 = 6'h2 == _T_11317_33; // @[Mux.scala 46:19:@10201.4]
  assign _T_13332 = _T_13331 ? _T_10366_1 : _T_13330; // @[Mux.scala 46:16:@10202.4]
  assign _T_13333 = 6'h1 == _T_11317_33; // @[Mux.scala 46:19:@10203.4]
  assign _T_13334 = _T_13333 ? _T_10366_0 : _T_13332; // @[Mux.scala 46:16:@10204.4]
  assign _T_13371 = 6'h23 == _T_11317_34; // @[Mux.scala 46:19:@10206.4]
  assign _T_13372 = _T_13371 ? _T_10366_34 : 8'h0; // @[Mux.scala 46:16:@10207.4]
  assign _T_13373 = 6'h22 == _T_11317_34; // @[Mux.scala 46:19:@10208.4]
  assign _T_13374 = _T_13373 ? _T_10366_33 : _T_13372; // @[Mux.scala 46:16:@10209.4]
  assign _T_13375 = 6'h21 == _T_11317_34; // @[Mux.scala 46:19:@10210.4]
  assign _T_13376 = _T_13375 ? _T_10366_32 : _T_13374; // @[Mux.scala 46:16:@10211.4]
  assign _T_13377 = 6'h20 == _T_11317_34; // @[Mux.scala 46:19:@10212.4]
  assign _T_13378 = _T_13377 ? _T_10366_31 : _T_13376; // @[Mux.scala 46:16:@10213.4]
  assign _T_13379 = 6'h1f == _T_11317_34; // @[Mux.scala 46:19:@10214.4]
  assign _T_13380 = _T_13379 ? _T_10366_30 : _T_13378; // @[Mux.scala 46:16:@10215.4]
  assign _T_13381 = 6'h1e == _T_11317_34; // @[Mux.scala 46:19:@10216.4]
  assign _T_13382 = _T_13381 ? _T_10366_29 : _T_13380; // @[Mux.scala 46:16:@10217.4]
  assign _T_13383 = 6'h1d == _T_11317_34; // @[Mux.scala 46:19:@10218.4]
  assign _T_13384 = _T_13383 ? _T_10366_28 : _T_13382; // @[Mux.scala 46:16:@10219.4]
  assign _T_13385 = 6'h1c == _T_11317_34; // @[Mux.scala 46:19:@10220.4]
  assign _T_13386 = _T_13385 ? _T_10366_27 : _T_13384; // @[Mux.scala 46:16:@10221.4]
  assign _T_13387 = 6'h1b == _T_11317_34; // @[Mux.scala 46:19:@10222.4]
  assign _T_13388 = _T_13387 ? _T_10366_26 : _T_13386; // @[Mux.scala 46:16:@10223.4]
  assign _T_13389 = 6'h1a == _T_11317_34; // @[Mux.scala 46:19:@10224.4]
  assign _T_13390 = _T_13389 ? _T_10366_25 : _T_13388; // @[Mux.scala 46:16:@10225.4]
  assign _T_13391 = 6'h19 == _T_11317_34; // @[Mux.scala 46:19:@10226.4]
  assign _T_13392 = _T_13391 ? _T_10366_24 : _T_13390; // @[Mux.scala 46:16:@10227.4]
  assign _T_13393 = 6'h18 == _T_11317_34; // @[Mux.scala 46:19:@10228.4]
  assign _T_13394 = _T_13393 ? _T_10366_23 : _T_13392; // @[Mux.scala 46:16:@10229.4]
  assign _T_13395 = 6'h17 == _T_11317_34; // @[Mux.scala 46:19:@10230.4]
  assign _T_13396 = _T_13395 ? _T_10366_22 : _T_13394; // @[Mux.scala 46:16:@10231.4]
  assign _T_13397 = 6'h16 == _T_11317_34; // @[Mux.scala 46:19:@10232.4]
  assign _T_13398 = _T_13397 ? _T_10366_21 : _T_13396; // @[Mux.scala 46:16:@10233.4]
  assign _T_13399 = 6'h15 == _T_11317_34; // @[Mux.scala 46:19:@10234.4]
  assign _T_13400 = _T_13399 ? _T_10366_20 : _T_13398; // @[Mux.scala 46:16:@10235.4]
  assign _T_13401 = 6'h14 == _T_11317_34; // @[Mux.scala 46:19:@10236.4]
  assign _T_13402 = _T_13401 ? _T_10366_19 : _T_13400; // @[Mux.scala 46:16:@10237.4]
  assign _T_13403 = 6'h13 == _T_11317_34; // @[Mux.scala 46:19:@10238.4]
  assign _T_13404 = _T_13403 ? _T_10366_18 : _T_13402; // @[Mux.scala 46:16:@10239.4]
  assign _T_13405 = 6'h12 == _T_11317_34; // @[Mux.scala 46:19:@10240.4]
  assign _T_13406 = _T_13405 ? _T_10366_17 : _T_13404; // @[Mux.scala 46:16:@10241.4]
  assign _T_13407 = 6'h11 == _T_11317_34; // @[Mux.scala 46:19:@10242.4]
  assign _T_13408 = _T_13407 ? _T_10366_16 : _T_13406; // @[Mux.scala 46:16:@10243.4]
  assign _T_13409 = 6'h10 == _T_11317_34; // @[Mux.scala 46:19:@10244.4]
  assign _T_13410 = _T_13409 ? _T_10366_15 : _T_13408; // @[Mux.scala 46:16:@10245.4]
  assign _T_13411 = 6'hf == _T_11317_34; // @[Mux.scala 46:19:@10246.4]
  assign _T_13412 = _T_13411 ? _T_10366_14 : _T_13410; // @[Mux.scala 46:16:@10247.4]
  assign _T_13413 = 6'he == _T_11317_34; // @[Mux.scala 46:19:@10248.4]
  assign _T_13414 = _T_13413 ? _T_10366_13 : _T_13412; // @[Mux.scala 46:16:@10249.4]
  assign _T_13415 = 6'hd == _T_11317_34; // @[Mux.scala 46:19:@10250.4]
  assign _T_13416 = _T_13415 ? _T_10366_12 : _T_13414; // @[Mux.scala 46:16:@10251.4]
  assign _T_13417 = 6'hc == _T_11317_34; // @[Mux.scala 46:19:@10252.4]
  assign _T_13418 = _T_13417 ? _T_10366_11 : _T_13416; // @[Mux.scala 46:16:@10253.4]
  assign _T_13419 = 6'hb == _T_11317_34; // @[Mux.scala 46:19:@10254.4]
  assign _T_13420 = _T_13419 ? _T_10366_10 : _T_13418; // @[Mux.scala 46:16:@10255.4]
  assign _T_13421 = 6'ha == _T_11317_34; // @[Mux.scala 46:19:@10256.4]
  assign _T_13422 = _T_13421 ? _T_10366_9 : _T_13420; // @[Mux.scala 46:16:@10257.4]
  assign _T_13423 = 6'h9 == _T_11317_34; // @[Mux.scala 46:19:@10258.4]
  assign _T_13424 = _T_13423 ? _T_10366_8 : _T_13422; // @[Mux.scala 46:16:@10259.4]
  assign _T_13425 = 6'h8 == _T_11317_34; // @[Mux.scala 46:19:@10260.4]
  assign _T_13426 = _T_13425 ? _T_10366_7 : _T_13424; // @[Mux.scala 46:16:@10261.4]
  assign _T_13427 = 6'h7 == _T_11317_34; // @[Mux.scala 46:19:@10262.4]
  assign _T_13428 = _T_13427 ? _T_10366_6 : _T_13426; // @[Mux.scala 46:16:@10263.4]
  assign _T_13429 = 6'h6 == _T_11317_34; // @[Mux.scala 46:19:@10264.4]
  assign _T_13430 = _T_13429 ? _T_10366_5 : _T_13428; // @[Mux.scala 46:16:@10265.4]
  assign _T_13431 = 6'h5 == _T_11317_34; // @[Mux.scala 46:19:@10266.4]
  assign _T_13432 = _T_13431 ? _T_10366_4 : _T_13430; // @[Mux.scala 46:16:@10267.4]
  assign _T_13433 = 6'h4 == _T_11317_34; // @[Mux.scala 46:19:@10268.4]
  assign _T_13434 = _T_13433 ? _T_10366_3 : _T_13432; // @[Mux.scala 46:16:@10269.4]
  assign _T_13435 = 6'h3 == _T_11317_34; // @[Mux.scala 46:19:@10270.4]
  assign _T_13436 = _T_13435 ? _T_10366_2 : _T_13434; // @[Mux.scala 46:16:@10271.4]
  assign _T_13437 = 6'h2 == _T_11317_34; // @[Mux.scala 46:19:@10272.4]
  assign _T_13438 = _T_13437 ? _T_10366_1 : _T_13436; // @[Mux.scala 46:16:@10273.4]
  assign _T_13439 = 6'h1 == _T_11317_34; // @[Mux.scala 46:19:@10274.4]
  assign _T_13440 = _T_13439 ? _T_10366_0 : _T_13438; // @[Mux.scala 46:16:@10275.4]
  assign _T_13478 = 6'h24 == _T_11317_35; // @[Mux.scala 46:19:@10277.4]
  assign _T_13479 = _T_13478 ? _T_10366_35 : 8'h0; // @[Mux.scala 46:16:@10278.4]
  assign _T_13480 = 6'h23 == _T_11317_35; // @[Mux.scala 46:19:@10279.4]
  assign _T_13481 = _T_13480 ? _T_10366_34 : _T_13479; // @[Mux.scala 46:16:@10280.4]
  assign _T_13482 = 6'h22 == _T_11317_35; // @[Mux.scala 46:19:@10281.4]
  assign _T_13483 = _T_13482 ? _T_10366_33 : _T_13481; // @[Mux.scala 46:16:@10282.4]
  assign _T_13484 = 6'h21 == _T_11317_35; // @[Mux.scala 46:19:@10283.4]
  assign _T_13485 = _T_13484 ? _T_10366_32 : _T_13483; // @[Mux.scala 46:16:@10284.4]
  assign _T_13486 = 6'h20 == _T_11317_35; // @[Mux.scala 46:19:@10285.4]
  assign _T_13487 = _T_13486 ? _T_10366_31 : _T_13485; // @[Mux.scala 46:16:@10286.4]
  assign _T_13488 = 6'h1f == _T_11317_35; // @[Mux.scala 46:19:@10287.4]
  assign _T_13489 = _T_13488 ? _T_10366_30 : _T_13487; // @[Mux.scala 46:16:@10288.4]
  assign _T_13490 = 6'h1e == _T_11317_35; // @[Mux.scala 46:19:@10289.4]
  assign _T_13491 = _T_13490 ? _T_10366_29 : _T_13489; // @[Mux.scala 46:16:@10290.4]
  assign _T_13492 = 6'h1d == _T_11317_35; // @[Mux.scala 46:19:@10291.4]
  assign _T_13493 = _T_13492 ? _T_10366_28 : _T_13491; // @[Mux.scala 46:16:@10292.4]
  assign _T_13494 = 6'h1c == _T_11317_35; // @[Mux.scala 46:19:@10293.4]
  assign _T_13495 = _T_13494 ? _T_10366_27 : _T_13493; // @[Mux.scala 46:16:@10294.4]
  assign _T_13496 = 6'h1b == _T_11317_35; // @[Mux.scala 46:19:@10295.4]
  assign _T_13497 = _T_13496 ? _T_10366_26 : _T_13495; // @[Mux.scala 46:16:@10296.4]
  assign _T_13498 = 6'h1a == _T_11317_35; // @[Mux.scala 46:19:@10297.4]
  assign _T_13499 = _T_13498 ? _T_10366_25 : _T_13497; // @[Mux.scala 46:16:@10298.4]
  assign _T_13500 = 6'h19 == _T_11317_35; // @[Mux.scala 46:19:@10299.4]
  assign _T_13501 = _T_13500 ? _T_10366_24 : _T_13499; // @[Mux.scala 46:16:@10300.4]
  assign _T_13502 = 6'h18 == _T_11317_35; // @[Mux.scala 46:19:@10301.4]
  assign _T_13503 = _T_13502 ? _T_10366_23 : _T_13501; // @[Mux.scala 46:16:@10302.4]
  assign _T_13504 = 6'h17 == _T_11317_35; // @[Mux.scala 46:19:@10303.4]
  assign _T_13505 = _T_13504 ? _T_10366_22 : _T_13503; // @[Mux.scala 46:16:@10304.4]
  assign _T_13506 = 6'h16 == _T_11317_35; // @[Mux.scala 46:19:@10305.4]
  assign _T_13507 = _T_13506 ? _T_10366_21 : _T_13505; // @[Mux.scala 46:16:@10306.4]
  assign _T_13508 = 6'h15 == _T_11317_35; // @[Mux.scala 46:19:@10307.4]
  assign _T_13509 = _T_13508 ? _T_10366_20 : _T_13507; // @[Mux.scala 46:16:@10308.4]
  assign _T_13510 = 6'h14 == _T_11317_35; // @[Mux.scala 46:19:@10309.4]
  assign _T_13511 = _T_13510 ? _T_10366_19 : _T_13509; // @[Mux.scala 46:16:@10310.4]
  assign _T_13512 = 6'h13 == _T_11317_35; // @[Mux.scala 46:19:@10311.4]
  assign _T_13513 = _T_13512 ? _T_10366_18 : _T_13511; // @[Mux.scala 46:16:@10312.4]
  assign _T_13514 = 6'h12 == _T_11317_35; // @[Mux.scala 46:19:@10313.4]
  assign _T_13515 = _T_13514 ? _T_10366_17 : _T_13513; // @[Mux.scala 46:16:@10314.4]
  assign _T_13516 = 6'h11 == _T_11317_35; // @[Mux.scala 46:19:@10315.4]
  assign _T_13517 = _T_13516 ? _T_10366_16 : _T_13515; // @[Mux.scala 46:16:@10316.4]
  assign _T_13518 = 6'h10 == _T_11317_35; // @[Mux.scala 46:19:@10317.4]
  assign _T_13519 = _T_13518 ? _T_10366_15 : _T_13517; // @[Mux.scala 46:16:@10318.4]
  assign _T_13520 = 6'hf == _T_11317_35; // @[Mux.scala 46:19:@10319.4]
  assign _T_13521 = _T_13520 ? _T_10366_14 : _T_13519; // @[Mux.scala 46:16:@10320.4]
  assign _T_13522 = 6'he == _T_11317_35; // @[Mux.scala 46:19:@10321.4]
  assign _T_13523 = _T_13522 ? _T_10366_13 : _T_13521; // @[Mux.scala 46:16:@10322.4]
  assign _T_13524 = 6'hd == _T_11317_35; // @[Mux.scala 46:19:@10323.4]
  assign _T_13525 = _T_13524 ? _T_10366_12 : _T_13523; // @[Mux.scala 46:16:@10324.4]
  assign _T_13526 = 6'hc == _T_11317_35; // @[Mux.scala 46:19:@10325.4]
  assign _T_13527 = _T_13526 ? _T_10366_11 : _T_13525; // @[Mux.scala 46:16:@10326.4]
  assign _T_13528 = 6'hb == _T_11317_35; // @[Mux.scala 46:19:@10327.4]
  assign _T_13529 = _T_13528 ? _T_10366_10 : _T_13527; // @[Mux.scala 46:16:@10328.4]
  assign _T_13530 = 6'ha == _T_11317_35; // @[Mux.scala 46:19:@10329.4]
  assign _T_13531 = _T_13530 ? _T_10366_9 : _T_13529; // @[Mux.scala 46:16:@10330.4]
  assign _T_13532 = 6'h9 == _T_11317_35; // @[Mux.scala 46:19:@10331.4]
  assign _T_13533 = _T_13532 ? _T_10366_8 : _T_13531; // @[Mux.scala 46:16:@10332.4]
  assign _T_13534 = 6'h8 == _T_11317_35; // @[Mux.scala 46:19:@10333.4]
  assign _T_13535 = _T_13534 ? _T_10366_7 : _T_13533; // @[Mux.scala 46:16:@10334.4]
  assign _T_13536 = 6'h7 == _T_11317_35; // @[Mux.scala 46:19:@10335.4]
  assign _T_13537 = _T_13536 ? _T_10366_6 : _T_13535; // @[Mux.scala 46:16:@10336.4]
  assign _T_13538 = 6'h6 == _T_11317_35; // @[Mux.scala 46:19:@10337.4]
  assign _T_13539 = _T_13538 ? _T_10366_5 : _T_13537; // @[Mux.scala 46:16:@10338.4]
  assign _T_13540 = 6'h5 == _T_11317_35; // @[Mux.scala 46:19:@10339.4]
  assign _T_13541 = _T_13540 ? _T_10366_4 : _T_13539; // @[Mux.scala 46:16:@10340.4]
  assign _T_13542 = 6'h4 == _T_11317_35; // @[Mux.scala 46:19:@10341.4]
  assign _T_13543 = _T_13542 ? _T_10366_3 : _T_13541; // @[Mux.scala 46:16:@10342.4]
  assign _T_13544 = 6'h3 == _T_11317_35; // @[Mux.scala 46:19:@10343.4]
  assign _T_13545 = _T_13544 ? _T_10366_2 : _T_13543; // @[Mux.scala 46:16:@10344.4]
  assign _T_13546 = 6'h2 == _T_11317_35; // @[Mux.scala 46:19:@10345.4]
  assign _T_13547 = _T_13546 ? _T_10366_1 : _T_13545; // @[Mux.scala 46:16:@10346.4]
  assign _T_13548 = 6'h1 == _T_11317_35; // @[Mux.scala 46:19:@10347.4]
  assign _T_13549 = _T_13548 ? _T_10366_0 : _T_13547; // @[Mux.scala 46:16:@10348.4]
  assign _T_13588 = 6'h25 == _T_11317_36; // @[Mux.scala 46:19:@10350.4]
  assign _T_13589 = _T_13588 ? _T_10366_36 : 8'h0; // @[Mux.scala 46:16:@10351.4]
  assign _T_13590 = 6'h24 == _T_11317_36; // @[Mux.scala 46:19:@10352.4]
  assign _T_13591 = _T_13590 ? _T_10366_35 : _T_13589; // @[Mux.scala 46:16:@10353.4]
  assign _T_13592 = 6'h23 == _T_11317_36; // @[Mux.scala 46:19:@10354.4]
  assign _T_13593 = _T_13592 ? _T_10366_34 : _T_13591; // @[Mux.scala 46:16:@10355.4]
  assign _T_13594 = 6'h22 == _T_11317_36; // @[Mux.scala 46:19:@10356.4]
  assign _T_13595 = _T_13594 ? _T_10366_33 : _T_13593; // @[Mux.scala 46:16:@10357.4]
  assign _T_13596 = 6'h21 == _T_11317_36; // @[Mux.scala 46:19:@10358.4]
  assign _T_13597 = _T_13596 ? _T_10366_32 : _T_13595; // @[Mux.scala 46:16:@10359.4]
  assign _T_13598 = 6'h20 == _T_11317_36; // @[Mux.scala 46:19:@10360.4]
  assign _T_13599 = _T_13598 ? _T_10366_31 : _T_13597; // @[Mux.scala 46:16:@10361.4]
  assign _T_13600 = 6'h1f == _T_11317_36; // @[Mux.scala 46:19:@10362.4]
  assign _T_13601 = _T_13600 ? _T_10366_30 : _T_13599; // @[Mux.scala 46:16:@10363.4]
  assign _T_13602 = 6'h1e == _T_11317_36; // @[Mux.scala 46:19:@10364.4]
  assign _T_13603 = _T_13602 ? _T_10366_29 : _T_13601; // @[Mux.scala 46:16:@10365.4]
  assign _T_13604 = 6'h1d == _T_11317_36; // @[Mux.scala 46:19:@10366.4]
  assign _T_13605 = _T_13604 ? _T_10366_28 : _T_13603; // @[Mux.scala 46:16:@10367.4]
  assign _T_13606 = 6'h1c == _T_11317_36; // @[Mux.scala 46:19:@10368.4]
  assign _T_13607 = _T_13606 ? _T_10366_27 : _T_13605; // @[Mux.scala 46:16:@10369.4]
  assign _T_13608 = 6'h1b == _T_11317_36; // @[Mux.scala 46:19:@10370.4]
  assign _T_13609 = _T_13608 ? _T_10366_26 : _T_13607; // @[Mux.scala 46:16:@10371.4]
  assign _T_13610 = 6'h1a == _T_11317_36; // @[Mux.scala 46:19:@10372.4]
  assign _T_13611 = _T_13610 ? _T_10366_25 : _T_13609; // @[Mux.scala 46:16:@10373.4]
  assign _T_13612 = 6'h19 == _T_11317_36; // @[Mux.scala 46:19:@10374.4]
  assign _T_13613 = _T_13612 ? _T_10366_24 : _T_13611; // @[Mux.scala 46:16:@10375.4]
  assign _T_13614 = 6'h18 == _T_11317_36; // @[Mux.scala 46:19:@10376.4]
  assign _T_13615 = _T_13614 ? _T_10366_23 : _T_13613; // @[Mux.scala 46:16:@10377.4]
  assign _T_13616 = 6'h17 == _T_11317_36; // @[Mux.scala 46:19:@10378.4]
  assign _T_13617 = _T_13616 ? _T_10366_22 : _T_13615; // @[Mux.scala 46:16:@10379.4]
  assign _T_13618 = 6'h16 == _T_11317_36; // @[Mux.scala 46:19:@10380.4]
  assign _T_13619 = _T_13618 ? _T_10366_21 : _T_13617; // @[Mux.scala 46:16:@10381.4]
  assign _T_13620 = 6'h15 == _T_11317_36; // @[Mux.scala 46:19:@10382.4]
  assign _T_13621 = _T_13620 ? _T_10366_20 : _T_13619; // @[Mux.scala 46:16:@10383.4]
  assign _T_13622 = 6'h14 == _T_11317_36; // @[Mux.scala 46:19:@10384.4]
  assign _T_13623 = _T_13622 ? _T_10366_19 : _T_13621; // @[Mux.scala 46:16:@10385.4]
  assign _T_13624 = 6'h13 == _T_11317_36; // @[Mux.scala 46:19:@10386.4]
  assign _T_13625 = _T_13624 ? _T_10366_18 : _T_13623; // @[Mux.scala 46:16:@10387.4]
  assign _T_13626 = 6'h12 == _T_11317_36; // @[Mux.scala 46:19:@10388.4]
  assign _T_13627 = _T_13626 ? _T_10366_17 : _T_13625; // @[Mux.scala 46:16:@10389.4]
  assign _T_13628 = 6'h11 == _T_11317_36; // @[Mux.scala 46:19:@10390.4]
  assign _T_13629 = _T_13628 ? _T_10366_16 : _T_13627; // @[Mux.scala 46:16:@10391.4]
  assign _T_13630 = 6'h10 == _T_11317_36; // @[Mux.scala 46:19:@10392.4]
  assign _T_13631 = _T_13630 ? _T_10366_15 : _T_13629; // @[Mux.scala 46:16:@10393.4]
  assign _T_13632 = 6'hf == _T_11317_36; // @[Mux.scala 46:19:@10394.4]
  assign _T_13633 = _T_13632 ? _T_10366_14 : _T_13631; // @[Mux.scala 46:16:@10395.4]
  assign _T_13634 = 6'he == _T_11317_36; // @[Mux.scala 46:19:@10396.4]
  assign _T_13635 = _T_13634 ? _T_10366_13 : _T_13633; // @[Mux.scala 46:16:@10397.4]
  assign _T_13636 = 6'hd == _T_11317_36; // @[Mux.scala 46:19:@10398.4]
  assign _T_13637 = _T_13636 ? _T_10366_12 : _T_13635; // @[Mux.scala 46:16:@10399.4]
  assign _T_13638 = 6'hc == _T_11317_36; // @[Mux.scala 46:19:@10400.4]
  assign _T_13639 = _T_13638 ? _T_10366_11 : _T_13637; // @[Mux.scala 46:16:@10401.4]
  assign _T_13640 = 6'hb == _T_11317_36; // @[Mux.scala 46:19:@10402.4]
  assign _T_13641 = _T_13640 ? _T_10366_10 : _T_13639; // @[Mux.scala 46:16:@10403.4]
  assign _T_13642 = 6'ha == _T_11317_36; // @[Mux.scala 46:19:@10404.4]
  assign _T_13643 = _T_13642 ? _T_10366_9 : _T_13641; // @[Mux.scala 46:16:@10405.4]
  assign _T_13644 = 6'h9 == _T_11317_36; // @[Mux.scala 46:19:@10406.4]
  assign _T_13645 = _T_13644 ? _T_10366_8 : _T_13643; // @[Mux.scala 46:16:@10407.4]
  assign _T_13646 = 6'h8 == _T_11317_36; // @[Mux.scala 46:19:@10408.4]
  assign _T_13647 = _T_13646 ? _T_10366_7 : _T_13645; // @[Mux.scala 46:16:@10409.4]
  assign _T_13648 = 6'h7 == _T_11317_36; // @[Mux.scala 46:19:@10410.4]
  assign _T_13649 = _T_13648 ? _T_10366_6 : _T_13647; // @[Mux.scala 46:16:@10411.4]
  assign _T_13650 = 6'h6 == _T_11317_36; // @[Mux.scala 46:19:@10412.4]
  assign _T_13651 = _T_13650 ? _T_10366_5 : _T_13649; // @[Mux.scala 46:16:@10413.4]
  assign _T_13652 = 6'h5 == _T_11317_36; // @[Mux.scala 46:19:@10414.4]
  assign _T_13653 = _T_13652 ? _T_10366_4 : _T_13651; // @[Mux.scala 46:16:@10415.4]
  assign _T_13654 = 6'h4 == _T_11317_36; // @[Mux.scala 46:19:@10416.4]
  assign _T_13655 = _T_13654 ? _T_10366_3 : _T_13653; // @[Mux.scala 46:16:@10417.4]
  assign _T_13656 = 6'h3 == _T_11317_36; // @[Mux.scala 46:19:@10418.4]
  assign _T_13657 = _T_13656 ? _T_10366_2 : _T_13655; // @[Mux.scala 46:16:@10419.4]
  assign _T_13658 = 6'h2 == _T_11317_36; // @[Mux.scala 46:19:@10420.4]
  assign _T_13659 = _T_13658 ? _T_10366_1 : _T_13657; // @[Mux.scala 46:16:@10421.4]
  assign _T_13660 = 6'h1 == _T_11317_36; // @[Mux.scala 46:19:@10422.4]
  assign _T_13661 = _T_13660 ? _T_10366_0 : _T_13659; // @[Mux.scala 46:16:@10423.4]
  assign _T_13701 = 6'h26 == _T_11317_37; // @[Mux.scala 46:19:@10425.4]
  assign _T_13702 = _T_13701 ? _T_10366_37 : 8'h0; // @[Mux.scala 46:16:@10426.4]
  assign _T_13703 = 6'h25 == _T_11317_37; // @[Mux.scala 46:19:@10427.4]
  assign _T_13704 = _T_13703 ? _T_10366_36 : _T_13702; // @[Mux.scala 46:16:@10428.4]
  assign _T_13705 = 6'h24 == _T_11317_37; // @[Mux.scala 46:19:@10429.4]
  assign _T_13706 = _T_13705 ? _T_10366_35 : _T_13704; // @[Mux.scala 46:16:@10430.4]
  assign _T_13707 = 6'h23 == _T_11317_37; // @[Mux.scala 46:19:@10431.4]
  assign _T_13708 = _T_13707 ? _T_10366_34 : _T_13706; // @[Mux.scala 46:16:@10432.4]
  assign _T_13709 = 6'h22 == _T_11317_37; // @[Mux.scala 46:19:@10433.4]
  assign _T_13710 = _T_13709 ? _T_10366_33 : _T_13708; // @[Mux.scala 46:16:@10434.4]
  assign _T_13711 = 6'h21 == _T_11317_37; // @[Mux.scala 46:19:@10435.4]
  assign _T_13712 = _T_13711 ? _T_10366_32 : _T_13710; // @[Mux.scala 46:16:@10436.4]
  assign _T_13713 = 6'h20 == _T_11317_37; // @[Mux.scala 46:19:@10437.4]
  assign _T_13714 = _T_13713 ? _T_10366_31 : _T_13712; // @[Mux.scala 46:16:@10438.4]
  assign _T_13715 = 6'h1f == _T_11317_37; // @[Mux.scala 46:19:@10439.4]
  assign _T_13716 = _T_13715 ? _T_10366_30 : _T_13714; // @[Mux.scala 46:16:@10440.4]
  assign _T_13717 = 6'h1e == _T_11317_37; // @[Mux.scala 46:19:@10441.4]
  assign _T_13718 = _T_13717 ? _T_10366_29 : _T_13716; // @[Mux.scala 46:16:@10442.4]
  assign _T_13719 = 6'h1d == _T_11317_37; // @[Mux.scala 46:19:@10443.4]
  assign _T_13720 = _T_13719 ? _T_10366_28 : _T_13718; // @[Mux.scala 46:16:@10444.4]
  assign _T_13721 = 6'h1c == _T_11317_37; // @[Mux.scala 46:19:@10445.4]
  assign _T_13722 = _T_13721 ? _T_10366_27 : _T_13720; // @[Mux.scala 46:16:@10446.4]
  assign _T_13723 = 6'h1b == _T_11317_37; // @[Mux.scala 46:19:@10447.4]
  assign _T_13724 = _T_13723 ? _T_10366_26 : _T_13722; // @[Mux.scala 46:16:@10448.4]
  assign _T_13725 = 6'h1a == _T_11317_37; // @[Mux.scala 46:19:@10449.4]
  assign _T_13726 = _T_13725 ? _T_10366_25 : _T_13724; // @[Mux.scala 46:16:@10450.4]
  assign _T_13727 = 6'h19 == _T_11317_37; // @[Mux.scala 46:19:@10451.4]
  assign _T_13728 = _T_13727 ? _T_10366_24 : _T_13726; // @[Mux.scala 46:16:@10452.4]
  assign _T_13729 = 6'h18 == _T_11317_37; // @[Mux.scala 46:19:@10453.4]
  assign _T_13730 = _T_13729 ? _T_10366_23 : _T_13728; // @[Mux.scala 46:16:@10454.4]
  assign _T_13731 = 6'h17 == _T_11317_37; // @[Mux.scala 46:19:@10455.4]
  assign _T_13732 = _T_13731 ? _T_10366_22 : _T_13730; // @[Mux.scala 46:16:@10456.4]
  assign _T_13733 = 6'h16 == _T_11317_37; // @[Mux.scala 46:19:@10457.4]
  assign _T_13734 = _T_13733 ? _T_10366_21 : _T_13732; // @[Mux.scala 46:16:@10458.4]
  assign _T_13735 = 6'h15 == _T_11317_37; // @[Mux.scala 46:19:@10459.4]
  assign _T_13736 = _T_13735 ? _T_10366_20 : _T_13734; // @[Mux.scala 46:16:@10460.4]
  assign _T_13737 = 6'h14 == _T_11317_37; // @[Mux.scala 46:19:@10461.4]
  assign _T_13738 = _T_13737 ? _T_10366_19 : _T_13736; // @[Mux.scala 46:16:@10462.4]
  assign _T_13739 = 6'h13 == _T_11317_37; // @[Mux.scala 46:19:@10463.4]
  assign _T_13740 = _T_13739 ? _T_10366_18 : _T_13738; // @[Mux.scala 46:16:@10464.4]
  assign _T_13741 = 6'h12 == _T_11317_37; // @[Mux.scala 46:19:@10465.4]
  assign _T_13742 = _T_13741 ? _T_10366_17 : _T_13740; // @[Mux.scala 46:16:@10466.4]
  assign _T_13743 = 6'h11 == _T_11317_37; // @[Mux.scala 46:19:@10467.4]
  assign _T_13744 = _T_13743 ? _T_10366_16 : _T_13742; // @[Mux.scala 46:16:@10468.4]
  assign _T_13745 = 6'h10 == _T_11317_37; // @[Mux.scala 46:19:@10469.4]
  assign _T_13746 = _T_13745 ? _T_10366_15 : _T_13744; // @[Mux.scala 46:16:@10470.4]
  assign _T_13747 = 6'hf == _T_11317_37; // @[Mux.scala 46:19:@10471.4]
  assign _T_13748 = _T_13747 ? _T_10366_14 : _T_13746; // @[Mux.scala 46:16:@10472.4]
  assign _T_13749 = 6'he == _T_11317_37; // @[Mux.scala 46:19:@10473.4]
  assign _T_13750 = _T_13749 ? _T_10366_13 : _T_13748; // @[Mux.scala 46:16:@10474.4]
  assign _T_13751 = 6'hd == _T_11317_37; // @[Mux.scala 46:19:@10475.4]
  assign _T_13752 = _T_13751 ? _T_10366_12 : _T_13750; // @[Mux.scala 46:16:@10476.4]
  assign _T_13753 = 6'hc == _T_11317_37; // @[Mux.scala 46:19:@10477.4]
  assign _T_13754 = _T_13753 ? _T_10366_11 : _T_13752; // @[Mux.scala 46:16:@10478.4]
  assign _T_13755 = 6'hb == _T_11317_37; // @[Mux.scala 46:19:@10479.4]
  assign _T_13756 = _T_13755 ? _T_10366_10 : _T_13754; // @[Mux.scala 46:16:@10480.4]
  assign _T_13757 = 6'ha == _T_11317_37; // @[Mux.scala 46:19:@10481.4]
  assign _T_13758 = _T_13757 ? _T_10366_9 : _T_13756; // @[Mux.scala 46:16:@10482.4]
  assign _T_13759 = 6'h9 == _T_11317_37; // @[Mux.scala 46:19:@10483.4]
  assign _T_13760 = _T_13759 ? _T_10366_8 : _T_13758; // @[Mux.scala 46:16:@10484.4]
  assign _T_13761 = 6'h8 == _T_11317_37; // @[Mux.scala 46:19:@10485.4]
  assign _T_13762 = _T_13761 ? _T_10366_7 : _T_13760; // @[Mux.scala 46:16:@10486.4]
  assign _T_13763 = 6'h7 == _T_11317_37; // @[Mux.scala 46:19:@10487.4]
  assign _T_13764 = _T_13763 ? _T_10366_6 : _T_13762; // @[Mux.scala 46:16:@10488.4]
  assign _T_13765 = 6'h6 == _T_11317_37; // @[Mux.scala 46:19:@10489.4]
  assign _T_13766 = _T_13765 ? _T_10366_5 : _T_13764; // @[Mux.scala 46:16:@10490.4]
  assign _T_13767 = 6'h5 == _T_11317_37; // @[Mux.scala 46:19:@10491.4]
  assign _T_13768 = _T_13767 ? _T_10366_4 : _T_13766; // @[Mux.scala 46:16:@10492.4]
  assign _T_13769 = 6'h4 == _T_11317_37; // @[Mux.scala 46:19:@10493.4]
  assign _T_13770 = _T_13769 ? _T_10366_3 : _T_13768; // @[Mux.scala 46:16:@10494.4]
  assign _T_13771 = 6'h3 == _T_11317_37; // @[Mux.scala 46:19:@10495.4]
  assign _T_13772 = _T_13771 ? _T_10366_2 : _T_13770; // @[Mux.scala 46:16:@10496.4]
  assign _T_13773 = 6'h2 == _T_11317_37; // @[Mux.scala 46:19:@10497.4]
  assign _T_13774 = _T_13773 ? _T_10366_1 : _T_13772; // @[Mux.scala 46:16:@10498.4]
  assign _T_13775 = 6'h1 == _T_11317_37; // @[Mux.scala 46:19:@10499.4]
  assign _T_13776 = _T_13775 ? _T_10366_0 : _T_13774; // @[Mux.scala 46:16:@10500.4]
  assign _T_13817 = 6'h27 == _T_11317_38; // @[Mux.scala 46:19:@10502.4]
  assign _T_13818 = _T_13817 ? _T_10366_38 : 8'h0; // @[Mux.scala 46:16:@10503.4]
  assign _T_13819 = 6'h26 == _T_11317_38; // @[Mux.scala 46:19:@10504.4]
  assign _T_13820 = _T_13819 ? _T_10366_37 : _T_13818; // @[Mux.scala 46:16:@10505.4]
  assign _T_13821 = 6'h25 == _T_11317_38; // @[Mux.scala 46:19:@10506.4]
  assign _T_13822 = _T_13821 ? _T_10366_36 : _T_13820; // @[Mux.scala 46:16:@10507.4]
  assign _T_13823 = 6'h24 == _T_11317_38; // @[Mux.scala 46:19:@10508.4]
  assign _T_13824 = _T_13823 ? _T_10366_35 : _T_13822; // @[Mux.scala 46:16:@10509.4]
  assign _T_13825 = 6'h23 == _T_11317_38; // @[Mux.scala 46:19:@10510.4]
  assign _T_13826 = _T_13825 ? _T_10366_34 : _T_13824; // @[Mux.scala 46:16:@10511.4]
  assign _T_13827 = 6'h22 == _T_11317_38; // @[Mux.scala 46:19:@10512.4]
  assign _T_13828 = _T_13827 ? _T_10366_33 : _T_13826; // @[Mux.scala 46:16:@10513.4]
  assign _T_13829 = 6'h21 == _T_11317_38; // @[Mux.scala 46:19:@10514.4]
  assign _T_13830 = _T_13829 ? _T_10366_32 : _T_13828; // @[Mux.scala 46:16:@10515.4]
  assign _T_13831 = 6'h20 == _T_11317_38; // @[Mux.scala 46:19:@10516.4]
  assign _T_13832 = _T_13831 ? _T_10366_31 : _T_13830; // @[Mux.scala 46:16:@10517.4]
  assign _T_13833 = 6'h1f == _T_11317_38; // @[Mux.scala 46:19:@10518.4]
  assign _T_13834 = _T_13833 ? _T_10366_30 : _T_13832; // @[Mux.scala 46:16:@10519.4]
  assign _T_13835 = 6'h1e == _T_11317_38; // @[Mux.scala 46:19:@10520.4]
  assign _T_13836 = _T_13835 ? _T_10366_29 : _T_13834; // @[Mux.scala 46:16:@10521.4]
  assign _T_13837 = 6'h1d == _T_11317_38; // @[Mux.scala 46:19:@10522.4]
  assign _T_13838 = _T_13837 ? _T_10366_28 : _T_13836; // @[Mux.scala 46:16:@10523.4]
  assign _T_13839 = 6'h1c == _T_11317_38; // @[Mux.scala 46:19:@10524.4]
  assign _T_13840 = _T_13839 ? _T_10366_27 : _T_13838; // @[Mux.scala 46:16:@10525.4]
  assign _T_13841 = 6'h1b == _T_11317_38; // @[Mux.scala 46:19:@10526.4]
  assign _T_13842 = _T_13841 ? _T_10366_26 : _T_13840; // @[Mux.scala 46:16:@10527.4]
  assign _T_13843 = 6'h1a == _T_11317_38; // @[Mux.scala 46:19:@10528.4]
  assign _T_13844 = _T_13843 ? _T_10366_25 : _T_13842; // @[Mux.scala 46:16:@10529.4]
  assign _T_13845 = 6'h19 == _T_11317_38; // @[Mux.scala 46:19:@10530.4]
  assign _T_13846 = _T_13845 ? _T_10366_24 : _T_13844; // @[Mux.scala 46:16:@10531.4]
  assign _T_13847 = 6'h18 == _T_11317_38; // @[Mux.scala 46:19:@10532.4]
  assign _T_13848 = _T_13847 ? _T_10366_23 : _T_13846; // @[Mux.scala 46:16:@10533.4]
  assign _T_13849 = 6'h17 == _T_11317_38; // @[Mux.scala 46:19:@10534.4]
  assign _T_13850 = _T_13849 ? _T_10366_22 : _T_13848; // @[Mux.scala 46:16:@10535.4]
  assign _T_13851 = 6'h16 == _T_11317_38; // @[Mux.scala 46:19:@10536.4]
  assign _T_13852 = _T_13851 ? _T_10366_21 : _T_13850; // @[Mux.scala 46:16:@10537.4]
  assign _T_13853 = 6'h15 == _T_11317_38; // @[Mux.scala 46:19:@10538.4]
  assign _T_13854 = _T_13853 ? _T_10366_20 : _T_13852; // @[Mux.scala 46:16:@10539.4]
  assign _T_13855 = 6'h14 == _T_11317_38; // @[Mux.scala 46:19:@10540.4]
  assign _T_13856 = _T_13855 ? _T_10366_19 : _T_13854; // @[Mux.scala 46:16:@10541.4]
  assign _T_13857 = 6'h13 == _T_11317_38; // @[Mux.scala 46:19:@10542.4]
  assign _T_13858 = _T_13857 ? _T_10366_18 : _T_13856; // @[Mux.scala 46:16:@10543.4]
  assign _T_13859 = 6'h12 == _T_11317_38; // @[Mux.scala 46:19:@10544.4]
  assign _T_13860 = _T_13859 ? _T_10366_17 : _T_13858; // @[Mux.scala 46:16:@10545.4]
  assign _T_13861 = 6'h11 == _T_11317_38; // @[Mux.scala 46:19:@10546.4]
  assign _T_13862 = _T_13861 ? _T_10366_16 : _T_13860; // @[Mux.scala 46:16:@10547.4]
  assign _T_13863 = 6'h10 == _T_11317_38; // @[Mux.scala 46:19:@10548.4]
  assign _T_13864 = _T_13863 ? _T_10366_15 : _T_13862; // @[Mux.scala 46:16:@10549.4]
  assign _T_13865 = 6'hf == _T_11317_38; // @[Mux.scala 46:19:@10550.4]
  assign _T_13866 = _T_13865 ? _T_10366_14 : _T_13864; // @[Mux.scala 46:16:@10551.4]
  assign _T_13867 = 6'he == _T_11317_38; // @[Mux.scala 46:19:@10552.4]
  assign _T_13868 = _T_13867 ? _T_10366_13 : _T_13866; // @[Mux.scala 46:16:@10553.4]
  assign _T_13869 = 6'hd == _T_11317_38; // @[Mux.scala 46:19:@10554.4]
  assign _T_13870 = _T_13869 ? _T_10366_12 : _T_13868; // @[Mux.scala 46:16:@10555.4]
  assign _T_13871 = 6'hc == _T_11317_38; // @[Mux.scala 46:19:@10556.4]
  assign _T_13872 = _T_13871 ? _T_10366_11 : _T_13870; // @[Mux.scala 46:16:@10557.4]
  assign _T_13873 = 6'hb == _T_11317_38; // @[Mux.scala 46:19:@10558.4]
  assign _T_13874 = _T_13873 ? _T_10366_10 : _T_13872; // @[Mux.scala 46:16:@10559.4]
  assign _T_13875 = 6'ha == _T_11317_38; // @[Mux.scala 46:19:@10560.4]
  assign _T_13876 = _T_13875 ? _T_10366_9 : _T_13874; // @[Mux.scala 46:16:@10561.4]
  assign _T_13877 = 6'h9 == _T_11317_38; // @[Mux.scala 46:19:@10562.4]
  assign _T_13878 = _T_13877 ? _T_10366_8 : _T_13876; // @[Mux.scala 46:16:@10563.4]
  assign _T_13879 = 6'h8 == _T_11317_38; // @[Mux.scala 46:19:@10564.4]
  assign _T_13880 = _T_13879 ? _T_10366_7 : _T_13878; // @[Mux.scala 46:16:@10565.4]
  assign _T_13881 = 6'h7 == _T_11317_38; // @[Mux.scala 46:19:@10566.4]
  assign _T_13882 = _T_13881 ? _T_10366_6 : _T_13880; // @[Mux.scala 46:16:@10567.4]
  assign _T_13883 = 6'h6 == _T_11317_38; // @[Mux.scala 46:19:@10568.4]
  assign _T_13884 = _T_13883 ? _T_10366_5 : _T_13882; // @[Mux.scala 46:16:@10569.4]
  assign _T_13885 = 6'h5 == _T_11317_38; // @[Mux.scala 46:19:@10570.4]
  assign _T_13886 = _T_13885 ? _T_10366_4 : _T_13884; // @[Mux.scala 46:16:@10571.4]
  assign _T_13887 = 6'h4 == _T_11317_38; // @[Mux.scala 46:19:@10572.4]
  assign _T_13888 = _T_13887 ? _T_10366_3 : _T_13886; // @[Mux.scala 46:16:@10573.4]
  assign _T_13889 = 6'h3 == _T_11317_38; // @[Mux.scala 46:19:@10574.4]
  assign _T_13890 = _T_13889 ? _T_10366_2 : _T_13888; // @[Mux.scala 46:16:@10575.4]
  assign _T_13891 = 6'h2 == _T_11317_38; // @[Mux.scala 46:19:@10576.4]
  assign _T_13892 = _T_13891 ? _T_10366_1 : _T_13890; // @[Mux.scala 46:16:@10577.4]
  assign _T_13893 = 6'h1 == _T_11317_38; // @[Mux.scala 46:19:@10578.4]
  assign _T_13894 = _T_13893 ? _T_10366_0 : _T_13892; // @[Mux.scala 46:16:@10579.4]
  assign _T_13936 = 6'h28 == _T_11317_39; // @[Mux.scala 46:19:@10581.4]
  assign _T_13937 = _T_13936 ? _T_10366_39 : 8'h0; // @[Mux.scala 46:16:@10582.4]
  assign _T_13938 = 6'h27 == _T_11317_39; // @[Mux.scala 46:19:@10583.4]
  assign _T_13939 = _T_13938 ? _T_10366_38 : _T_13937; // @[Mux.scala 46:16:@10584.4]
  assign _T_13940 = 6'h26 == _T_11317_39; // @[Mux.scala 46:19:@10585.4]
  assign _T_13941 = _T_13940 ? _T_10366_37 : _T_13939; // @[Mux.scala 46:16:@10586.4]
  assign _T_13942 = 6'h25 == _T_11317_39; // @[Mux.scala 46:19:@10587.4]
  assign _T_13943 = _T_13942 ? _T_10366_36 : _T_13941; // @[Mux.scala 46:16:@10588.4]
  assign _T_13944 = 6'h24 == _T_11317_39; // @[Mux.scala 46:19:@10589.4]
  assign _T_13945 = _T_13944 ? _T_10366_35 : _T_13943; // @[Mux.scala 46:16:@10590.4]
  assign _T_13946 = 6'h23 == _T_11317_39; // @[Mux.scala 46:19:@10591.4]
  assign _T_13947 = _T_13946 ? _T_10366_34 : _T_13945; // @[Mux.scala 46:16:@10592.4]
  assign _T_13948 = 6'h22 == _T_11317_39; // @[Mux.scala 46:19:@10593.4]
  assign _T_13949 = _T_13948 ? _T_10366_33 : _T_13947; // @[Mux.scala 46:16:@10594.4]
  assign _T_13950 = 6'h21 == _T_11317_39; // @[Mux.scala 46:19:@10595.4]
  assign _T_13951 = _T_13950 ? _T_10366_32 : _T_13949; // @[Mux.scala 46:16:@10596.4]
  assign _T_13952 = 6'h20 == _T_11317_39; // @[Mux.scala 46:19:@10597.4]
  assign _T_13953 = _T_13952 ? _T_10366_31 : _T_13951; // @[Mux.scala 46:16:@10598.4]
  assign _T_13954 = 6'h1f == _T_11317_39; // @[Mux.scala 46:19:@10599.4]
  assign _T_13955 = _T_13954 ? _T_10366_30 : _T_13953; // @[Mux.scala 46:16:@10600.4]
  assign _T_13956 = 6'h1e == _T_11317_39; // @[Mux.scala 46:19:@10601.4]
  assign _T_13957 = _T_13956 ? _T_10366_29 : _T_13955; // @[Mux.scala 46:16:@10602.4]
  assign _T_13958 = 6'h1d == _T_11317_39; // @[Mux.scala 46:19:@10603.4]
  assign _T_13959 = _T_13958 ? _T_10366_28 : _T_13957; // @[Mux.scala 46:16:@10604.4]
  assign _T_13960 = 6'h1c == _T_11317_39; // @[Mux.scala 46:19:@10605.4]
  assign _T_13961 = _T_13960 ? _T_10366_27 : _T_13959; // @[Mux.scala 46:16:@10606.4]
  assign _T_13962 = 6'h1b == _T_11317_39; // @[Mux.scala 46:19:@10607.4]
  assign _T_13963 = _T_13962 ? _T_10366_26 : _T_13961; // @[Mux.scala 46:16:@10608.4]
  assign _T_13964 = 6'h1a == _T_11317_39; // @[Mux.scala 46:19:@10609.4]
  assign _T_13965 = _T_13964 ? _T_10366_25 : _T_13963; // @[Mux.scala 46:16:@10610.4]
  assign _T_13966 = 6'h19 == _T_11317_39; // @[Mux.scala 46:19:@10611.4]
  assign _T_13967 = _T_13966 ? _T_10366_24 : _T_13965; // @[Mux.scala 46:16:@10612.4]
  assign _T_13968 = 6'h18 == _T_11317_39; // @[Mux.scala 46:19:@10613.4]
  assign _T_13969 = _T_13968 ? _T_10366_23 : _T_13967; // @[Mux.scala 46:16:@10614.4]
  assign _T_13970 = 6'h17 == _T_11317_39; // @[Mux.scala 46:19:@10615.4]
  assign _T_13971 = _T_13970 ? _T_10366_22 : _T_13969; // @[Mux.scala 46:16:@10616.4]
  assign _T_13972 = 6'h16 == _T_11317_39; // @[Mux.scala 46:19:@10617.4]
  assign _T_13973 = _T_13972 ? _T_10366_21 : _T_13971; // @[Mux.scala 46:16:@10618.4]
  assign _T_13974 = 6'h15 == _T_11317_39; // @[Mux.scala 46:19:@10619.4]
  assign _T_13975 = _T_13974 ? _T_10366_20 : _T_13973; // @[Mux.scala 46:16:@10620.4]
  assign _T_13976 = 6'h14 == _T_11317_39; // @[Mux.scala 46:19:@10621.4]
  assign _T_13977 = _T_13976 ? _T_10366_19 : _T_13975; // @[Mux.scala 46:16:@10622.4]
  assign _T_13978 = 6'h13 == _T_11317_39; // @[Mux.scala 46:19:@10623.4]
  assign _T_13979 = _T_13978 ? _T_10366_18 : _T_13977; // @[Mux.scala 46:16:@10624.4]
  assign _T_13980 = 6'h12 == _T_11317_39; // @[Mux.scala 46:19:@10625.4]
  assign _T_13981 = _T_13980 ? _T_10366_17 : _T_13979; // @[Mux.scala 46:16:@10626.4]
  assign _T_13982 = 6'h11 == _T_11317_39; // @[Mux.scala 46:19:@10627.4]
  assign _T_13983 = _T_13982 ? _T_10366_16 : _T_13981; // @[Mux.scala 46:16:@10628.4]
  assign _T_13984 = 6'h10 == _T_11317_39; // @[Mux.scala 46:19:@10629.4]
  assign _T_13985 = _T_13984 ? _T_10366_15 : _T_13983; // @[Mux.scala 46:16:@10630.4]
  assign _T_13986 = 6'hf == _T_11317_39; // @[Mux.scala 46:19:@10631.4]
  assign _T_13987 = _T_13986 ? _T_10366_14 : _T_13985; // @[Mux.scala 46:16:@10632.4]
  assign _T_13988 = 6'he == _T_11317_39; // @[Mux.scala 46:19:@10633.4]
  assign _T_13989 = _T_13988 ? _T_10366_13 : _T_13987; // @[Mux.scala 46:16:@10634.4]
  assign _T_13990 = 6'hd == _T_11317_39; // @[Mux.scala 46:19:@10635.4]
  assign _T_13991 = _T_13990 ? _T_10366_12 : _T_13989; // @[Mux.scala 46:16:@10636.4]
  assign _T_13992 = 6'hc == _T_11317_39; // @[Mux.scala 46:19:@10637.4]
  assign _T_13993 = _T_13992 ? _T_10366_11 : _T_13991; // @[Mux.scala 46:16:@10638.4]
  assign _T_13994 = 6'hb == _T_11317_39; // @[Mux.scala 46:19:@10639.4]
  assign _T_13995 = _T_13994 ? _T_10366_10 : _T_13993; // @[Mux.scala 46:16:@10640.4]
  assign _T_13996 = 6'ha == _T_11317_39; // @[Mux.scala 46:19:@10641.4]
  assign _T_13997 = _T_13996 ? _T_10366_9 : _T_13995; // @[Mux.scala 46:16:@10642.4]
  assign _T_13998 = 6'h9 == _T_11317_39; // @[Mux.scala 46:19:@10643.4]
  assign _T_13999 = _T_13998 ? _T_10366_8 : _T_13997; // @[Mux.scala 46:16:@10644.4]
  assign _T_14000 = 6'h8 == _T_11317_39; // @[Mux.scala 46:19:@10645.4]
  assign _T_14001 = _T_14000 ? _T_10366_7 : _T_13999; // @[Mux.scala 46:16:@10646.4]
  assign _T_14002 = 6'h7 == _T_11317_39; // @[Mux.scala 46:19:@10647.4]
  assign _T_14003 = _T_14002 ? _T_10366_6 : _T_14001; // @[Mux.scala 46:16:@10648.4]
  assign _T_14004 = 6'h6 == _T_11317_39; // @[Mux.scala 46:19:@10649.4]
  assign _T_14005 = _T_14004 ? _T_10366_5 : _T_14003; // @[Mux.scala 46:16:@10650.4]
  assign _T_14006 = 6'h5 == _T_11317_39; // @[Mux.scala 46:19:@10651.4]
  assign _T_14007 = _T_14006 ? _T_10366_4 : _T_14005; // @[Mux.scala 46:16:@10652.4]
  assign _T_14008 = 6'h4 == _T_11317_39; // @[Mux.scala 46:19:@10653.4]
  assign _T_14009 = _T_14008 ? _T_10366_3 : _T_14007; // @[Mux.scala 46:16:@10654.4]
  assign _T_14010 = 6'h3 == _T_11317_39; // @[Mux.scala 46:19:@10655.4]
  assign _T_14011 = _T_14010 ? _T_10366_2 : _T_14009; // @[Mux.scala 46:16:@10656.4]
  assign _T_14012 = 6'h2 == _T_11317_39; // @[Mux.scala 46:19:@10657.4]
  assign _T_14013 = _T_14012 ? _T_10366_1 : _T_14011; // @[Mux.scala 46:16:@10658.4]
  assign _T_14014 = 6'h1 == _T_11317_39; // @[Mux.scala 46:19:@10659.4]
  assign _T_14015 = _T_14014 ? _T_10366_0 : _T_14013; // @[Mux.scala 46:16:@10660.4]
  assign _T_14058 = 6'h29 == _T_11317_40; // @[Mux.scala 46:19:@10662.4]
  assign _T_14059 = _T_14058 ? _T_10366_40 : 8'h0; // @[Mux.scala 46:16:@10663.4]
  assign _T_14060 = 6'h28 == _T_11317_40; // @[Mux.scala 46:19:@10664.4]
  assign _T_14061 = _T_14060 ? _T_10366_39 : _T_14059; // @[Mux.scala 46:16:@10665.4]
  assign _T_14062 = 6'h27 == _T_11317_40; // @[Mux.scala 46:19:@10666.4]
  assign _T_14063 = _T_14062 ? _T_10366_38 : _T_14061; // @[Mux.scala 46:16:@10667.4]
  assign _T_14064 = 6'h26 == _T_11317_40; // @[Mux.scala 46:19:@10668.4]
  assign _T_14065 = _T_14064 ? _T_10366_37 : _T_14063; // @[Mux.scala 46:16:@10669.4]
  assign _T_14066 = 6'h25 == _T_11317_40; // @[Mux.scala 46:19:@10670.4]
  assign _T_14067 = _T_14066 ? _T_10366_36 : _T_14065; // @[Mux.scala 46:16:@10671.4]
  assign _T_14068 = 6'h24 == _T_11317_40; // @[Mux.scala 46:19:@10672.4]
  assign _T_14069 = _T_14068 ? _T_10366_35 : _T_14067; // @[Mux.scala 46:16:@10673.4]
  assign _T_14070 = 6'h23 == _T_11317_40; // @[Mux.scala 46:19:@10674.4]
  assign _T_14071 = _T_14070 ? _T_10366_34 : _T_14069; // @[Mux.scala 46:16:@10675.4]
  assign _T_14072 = 6'h22 == _T_11317_40; // @[Mux.scala 46:19:@10676.4]
  assign _T_14073 = _T_14072 ? _T_10366_33 : _T_14071; // @[Mux.scala 46:16:@10677.4]
  assign _T_14074 = 6'h21 == _T_11317_40; // @[Mux.scala 46:19:@10678.4]
  assign _T_14075 = _T_14074 ? _T_10366_32 : _T_14073; // @[Mux.scala 46:16:@10679.4]
  assign _T_14076 = 6'h20 == _T_11317_40; // @[Mux.scala 46:19:@10680.4]
  assign _T_14077 = _T_14076 ? _T_10366_31 : _T_14075; // @[Mux.scala 46:16:@10681.4]
  assign _T_14078 = 6'h1f == _T_11317_40; // @[Mux.scala 46:19:@10682.4]
  assign _T_14079 = _T_14078 ? _T_10366_30 : _T_14077; // @[Mux.scala 46:16:@10683.4]
  assign _T_14080 = 6'h1e == _T_11317_40; // @[Mux.scala 46:19:@10684.4]
  assign _T_14081 = _T_14080 ? _T_10366_29 : _T_14079; // @[Mux.scala 46:16:@10685.4]
  assign _T_14082 = 6'h1d == _T_11317_40; // @[Mux.scala 46:19:@10686.4]
  assign _T_14083 = _T_14082 ? _T_10366_28 : _T_14081; // @[Mux.scala 46:16:@10687.4]
  assign _T_14084 = 6'h1c == _T_11317_40; // @[Mux.scala 46:19:@10688.4]
  assign _T_14085 = _T_14084 ? _T_10366_27 : _T_14083; // @[Mux.scala 46:16:@10689.4]
  assign _T_14086 = 6'h1b == _T_11317_40; // @[Mux.scala 46:19:@10690.4]
  assign _T_14087 = _T_14086 ? _T_10366_26 : _T_14085; // @[Mux.scala 46:16:@10691.4]
  assign _T_14088 = 6'h1a == _T_11317_40; // @[Mux.scala 46:19:@10692.4]
  assign _T_14089 = _T_14088 ? _T_10366_25 : _T_14087; // @[Mux.scala 46:16:@10693.4]
  assign _T_14090 = 6'h19 == _T_11317_40; // @[Mux.scala 46:19:@10694.4]
  assign _T_14091 = _T_14090 ? _T_10366_24 : _T_14089; // @[Mux.scala 46:16:@10695.4]
  assign _T_14092 = 6'h18 == _T_11317_40; // @[Mux.scala 46:19:@10696.4]
  assign _T_14093 = _T_14092 ? _T_10366_23 : _T_14091; // @[Mux.scala 46:16:@10697.4]
  assign _T_14094 = 6'h17 == _T_11317_40; // @[Mux.scala 46:19:@10698.4]
  assign _T_14095 = _T_14094 ? _T_10366_22 : _T_14093; // @[Mux.scala 46:16:@10699.4]
  assign _T_14096 = 6'h16 == _T_11317_40; // @[Mux.scala 46:19:@10700.4]
  assign _T_14097 = _T_14096 ? _T_10366_21 : _T_14095; // @[Mux.scala 46:16:@10701.4]
  assign _T_14098 = 6'h15 == _T_11317_40; // @[Mux.scala 46:19:@10702.4]
  assign _T_14099 = _T_14098 ? _T_10366_20 : _T_14097; // @[Mux.scala 46:16:@10703.4]
  assign _T_14100 = 6'h14 == _T_11317_40; // @[Mux.scala 46:19:@10704.4]
  assign _T_14101 = _T_14100 ? _T_10366_19 : _T_14099; // @[Mux.scala 46:16:@10705.4]
  assign _T_14102 = 6'h13 == _T_11317_40; // @[Mux.scala 46:19:@10706.4]
  assign _T_14103 = _T_14102 ? _T_10366_18 : _T_14101; // @[Mux.scala 46:16:@10707.4]
  assign _T_14104 = 6'h12 == _T_11317_40; // @[Mux.scala 46:19:@10708.4]
  assign _T_14105 = _T_14104 ? _T_10366_17 : _T_14103; // @[Mux.scala 46:16:@10709.4]
  assign _T_14106 = 6'h11 == _T_11317_40; // @[Mux.scala 46:19:@10710.4]
  assign _T_14107 = _T_14106 ? _T_10366_16 : _T_14105; // @[Mux.scala 46:16:@10711.4]
  assign _T_14108 = 6'h10 == _T_11317_40; // @[Mux.scala 46:19:@10712.4]
  assign _T_14109 = _T_14108 ? _T_10366_15 : _T_14107; // @[Mux.scala 46:16:@10713.4]
  assign _T_14110 = 6'hf == _T_11317_40; // @[Mux.scala 46:19:@10714.4]
  assign _T_14111 = _T_14110 ? _T_10366_14 : _T_14109; // @[Mux.scala 46:16:@10715.4]
  assign _T_14112 = 6'he == _T_11317_40; // @[Mux.scala 46:19:@10716.4]
  assign _T_14113 = _T_14112 ? _T_10366_13 : _T_14111; // @[Mux.scala 46:16:@10717.4]
  assign _T_14114 = 6'hd == _T_11317_40; // @[Mux.scala 46:19:@10718.4]
  assign _T_14115 = _T_14114 ? _T_10366_12 : _T_14113; // @[Mux.scala 46:16:@10719.4]
  assign _T_14116 = 6'hc == _T_11317_40; // @[Mux.scala 46:19:@10720.4]
  assign _T_14117 = _T_14116 ? _T_10366_11 : _T_14115; // @[Mux.scala 46:16:@10721.4]
  assign _T_14118 = 6'hb == _T_11317_40; // @[Mux.scala 46:19:@10722.4]
  assign _T_14119 = _T_14118 ? _T_10366_10 : _T_14117; // @[Mux.scala 46:16:@10723.4]
  assign _T_14120 = 6'ha == _T_11317_40; // @[Mux.scala 46:19:@10724.4]
  assign _T_14121 = _T_14120 ? _T_10366_9 : _T_14119; // @[Mux.scala 46:16:@10725.4]
  assign _T_14122 = 6'h9 == _T_11317_40; // @[Mux.scala 46:19:@10726.4]
  assign _T_14123 = _T_14122 ? _T_10366_8 : _T_14121; // @[Mux.scala 46:16:@10727.4]
  assign _T_14124 = 6'h8 == _T_11317_40; // @[Mux.scala 46:19:@10728.4]
  assign _T_14125 = _T_14124 ? _T_10366_7 : _T_14123; // @[Mux.scala 46:16:@10729.4]
  assign _T_14126 = 6'h7 == _T_11317_40; // @[Mux.scala 46:19:@10730.4]
  assign _T_14127 = _T_14126 ? _T_10366_6 : _T_14125; // @[Mux.scala 46:16:@10731.4]
  assign _T_14128 = 6'h6 == _T_11317_40; // @[Mux.scala 46:19:@10732.4]
  assign _T_14129 = _T_14128 ? _T_10366_5 : _T_14127; // @[Mux.scala 46:16:@10733.4]
  assign _T_14130 = 6'h5 == _T_11317_40; // @[Mux.scala 46:19:@10734.4]
  assign _T_14131 = _T_14130 ? _T_10366_4 : _T_14129; // @[Mux.scala 46:16:@10735.4]
  assign _T_14132 = 6'h4 == _T_11317_40; // @[Mux.scala 46:19:@10736.4]
  assign _T_14133 = _T_14132 ? _T_10366_3 : _T_14131; // @[Mux.scala 46:16:@10737.4]
  assign _T_14134 = 6'h3 == _T_11317_40; // @[Mux.scala 46:19:@10738.4]
  assign _T_14135 = _T_14134 ? _T_10366_2 : _T_14133; // @[Mux.scala 46:16:@10739.4]
  assign _T_14136 = 6'h2 == _T_11317_40; // @[Mux.scala 46:19:@10740.4]
  assign _T_14137 = _T_14136 ? _T_10366_1 : _T_14135; // @[Mux.scala 46:16:@10741.4]
  assign _T_14138 = 6'h1 == _T_11317_40; // @[Mux.scala 46:19:@10742.4]
  assign _T_14139 = _T_14138 ? _T_10366_0 : _T_14137; // @[Mux.scala 46:16:@10743.4]
  assign _T_14183 = 6'h2a == _T_11317_41; // @[Mux.scala 46:19:@10745.4]
  assign _T_14184 = _T_14183 ? _T_10366_41 : 8'h0; // @[Mux.scala 46:16:@10746.4]
  assign _T_14185 = 6'h29 == _T_11317_41; // @[Mux.scala 46:19:@10747.4]
  assign _T_14186 = _T_14185 ? _T_10366_40 : _T_14184; // @[Mux.scala 46:16:@10748.4]
  assign _T_14187 = 6'h28 == _T_11317_41; // @[Mux.scala 46:19:@10749.4]
  assign _T_14188 = _T_14187 ? _T_10366_39 : _T_14186; // @[Mux.scala 46:16:@10750.4]
  assign _T_14189 = 6'h27 == _T_11317_41; // @[Mux.scala 46:19:@10751.4]
  assign _T_14190 = _T_14189 ? _T_10366_38 : _T_14188; // @[Mux.scala 46:16:@10752.4]
  assign _T_14191 = 6'h26 == _T_11317_41; // @[Mux.scala 46:19:@10753.4]
  assign _T_14192 = _T_14191 ? _T_10366_37 : _T_14190; // @[Mux.scala 46:16:@10754.4]
  assign _T_14193 = 6'h25 == _T_11317_41; // @[Mux.scala 46:19:@10755.4]
  assign _T_14194 = _T_14193 ? _T_10366_36 : _T_14192; // @[Mux.scala 46:16:@10756.4]
  assign _T_14195 = 6'h24 == _T_11317_41; // @[Mux.scala 46:19:@10757.4]
  assign _T_14196 = _T_14195 ? _T_10366_35 : _T_14194; // @[Mux.scala 46:16:@10758.4]
  assign _T_14197 = 6'h23 == _T_11317_41; // @[Mux.scala 46:19:@10759.4]
  assign _T_14198 = _T_14197 ? _T_10366_34 : _T_14196; // @[Mux.scala 46:16:@10760.4]
  assign _T_14199 = 6'h22 == _T_11317_41; // @[Mux.scala 46:19:@10761.4]
  assign _T_14200 = _T_14199 ? _T_10366_33 : _T_14198; // @[Mux.scala 46:16:@10762.4]
  assign _T_14201 = 6'h21 == _T_11317_41; // @[Mux.scala 46:19:@10763.4]
  assign _T_14202 = _T_14201 ? _T_10366_32 : _T_14200; // @[Mux.scala 46:16:@10764.4]
  assign _T_14203 = 6'h20 == _T_11317_41; // @[Mux.scala 46:19:@10765.4]
  assign _T_14204 = _T_14203 ? _T_10366_31 : _T_14202; // @[Mux.scala 46:16:@10766.4]
  assign _T_14205 = 6'h1f == _T_11317_41; // @[Mux.scala 46:19:@10767.4]
  assign _T_14206 = _T_14205 ? _T_10366_30 : _T_14204; // @[Mux.scala 46:16:@10768.4]
  assign _T_14207 = 6'h1e == _T_11317_41; // @[Mux.scala 46:19:@10769.4]
  assign _T_14208 = _T_14207 ? _T_10366_29 : _T_14206; // @[Mux.scala 46:16:@10770.4]
  assign _T_14209 = 6'h1d == _T_11317_41; // @[Mux.scala 46:19:@10771.4]
  assign _T_14210 = _T_14209 ? _T_10366_28 : _T_14208; // @[Mux.scala 46:16:@10772.4]
  assign _T_14211 = 6'h1c == _T_11317_41; // @[Mux.scala 46:19:@10773.4]
  assign _T_14212 = _T_14211 ? _T_10366_27 : _T_14210; // @[Mux.scala 46:16:@10774.4]
  assign _T_14213 = 6'h1b == _T_11317_41; // @[Mux.scala 46:19:@10775.4]
  assign _T_14214 = _T_14213 ? _T_10366_26 : _T_14212; // @[Mux.scala 46:16:@10776.4]
  assign _T_14215 = 6'h1a == _T_11317_41; // @[Mux.scala 46:19:@10777.4]
  assign _T_14216 = _T_14215 ? _T_10366_25 : _T_14214; // @[Mux.scala 46:16:@10778.4]
  assign _T_14217 = 6'h19 == _T_11317_41; // @[Mux.scala 46:19:@10779.4]
  assign _T_14218 = _T_14217 ? _T_10366_24 : _T_14216; // @[Mux.scala 46:16:@10780.4]
  assign _T_14219 = 6'h18 == _T_11317_41; // @[Mux.scala 46:19:@10781.4]
  assign _T_14220 = _T_14219 ? _T_10366_23 : _T_14218; // @[Mux.scala 46:16:@10782.4]
  assign _T_14221 = 6'h17 == _T_11317_41; // @[Mux.scala 46:19:@10783.4]
  assign _T_14222 = _T_14221 ? _T_10366_22 : _T_14220; // @[Mux.scala 46:16:@10784.4]
  assign _T_14223 = 6'h16 == _T_11317_41; // @[Mux.scala 46:19:@10785.4]
  assign _T_14224 = _T_14223 ? _T_10366_21 : _T_14222; // @[Mux.scala 46:16:@10786.4]
  assign _T_14225 = 6'h15 == _T_11317_41; // @[Mux.scala 46:19:@10787.4]
  assign _T_14226 = _T_14225 ? _T_10366_20 : _T_14224; // @[Mux.scala 46:16:@10788.4]
  assign _T_14227 = 6'h14 == _T_11317_41; // @[Mux.scala 46:19:@10789.4]
  assign _T_14228 = _T_14227 ? _T_10366_19 : _T_14226; // @[Mux.scala 46:16:@10790.4]
  assign _T_14229 = 6'h13 == _T_11317_41; // @[Mux.scala 46:19:@10791.4]
  assign _T_14230 = _T_14229 ? _T_10366_18 : _T_14228; // @[Mux.scala 46:16:@10792.4]
  assign _T_14231 = 6'h12 == _T_11317_41; // @[Mux.scala 46:19:@10793.4]
  assign _T_14232 = _T_14231 ? _T_10366_17 : _T_14230; // @[Mux.scala 46:16:@10794.4]
  assign _T_14233 = 6'h11 == _T_11317_41; // @[Mux.scala 46:19:@10795.4]
  assign _T_14234 = _T_14233 ? _T_10366_16 : _T_14232; // @[Mux.scala 46:16:@10796.4]
  assign _T_14235 = 6'h10 == _T_11317_41; // @[Mux.scala 46:19:@10797.4]
  assign _T_14236 = _T_14235 ? _T_10366_15 : _T_14234; // @[Mux.scala 46:16:@10798.4]
  assign _T_14237 = 6'hf == _T_11317_41; // @[Mux.scala 46:19:@10799.4]
  assign _T_14238 = _T_14237 ? _T_10366_14 : _T_14236; // @[Mux.scala 46:16:@10800.4]
  assign _T_14239 = 6'he == _T_11317_41; // @[Mux.scala 46:19:@10801.4]
  assign _T_14240 = _T_14239 ? _T_10366_13 : _T_14238; // @[Mux.scala 46:16:@10802.4]
  assign _T_14241 = 6'hd == _T_11317_41; // @[Mux.scala 46:19:@10803.4]
  assign _T_14242 = _T_14241 ? _T_10366_12 : _T_14240; // @[Mux.scala 46:16:@10804.4]
  assign _T_14243 = 6'hc == _T_11317_41; // @[Mux.scala 46:19:@10805.4]
  assign _T_14244 = _T_14243 ? _T_10366_11 : _T_14242; // @[Mux.scala 46:16:@10806.4]
  assign _T_14245 = 6'hb == _T_11317_41; // @[Mux.scala 46:19:@10807.4]
  assign _T_14246 = _T_14245 ? _T_10366_10 : _T_14244; // @[Mux.scala 46:16:@10808.4]
  assign _T_14247 = 6'ha == _T_11317_41; // @[Mux.scala 46:19:@10809.4]
  assign _T_14248 = _T_14247 ? _T_10366_9 : _T_14246; // @[Mux.scala 46:16:@10810.4]
  assign _T_14249 = 6'h9 == _T_11317_41; // @[Mux.scala 46:19:@10811.4]
  assign _T_14250 = _T_14249 ? _T_10366_8 : _T_14248; // @[Mux.scala 46:16:@10812.4]
  assign _T_14251 = 6'h8 == _T_11317_41; // @[Mux.scala 46:19:@10813.4]
  assign _T_14252 = _T_14251 ? _T_10366_7 : _T_14250; // @[Mux.scala 46:16:@10814.4]
  assign _T_14253 = 6'h7 == _T_11317_41; // @[Mux.scala 46:19:@10815.4]
  assign _T_14254 = _T_14253 ? _T_10366_6 : _T_14252; // @[Mux.scala 46:16:@10816.4]
  assign _T_14255 = 6'h6 == _T_11317_41; // @[Mux.scala 46:19:@10817.4]
  assign _T_14256 = _T_14255 ? _T_10366_5 : _T_14254; // @[Mux.scala 46:16:@10818.4]
  assign _T_14257 = 6'h5 == _T_11317_41; // @[Mux.scala 46:19:@10819.4]
  assign _T_14258 = _T_14257 ? _T_10366_4 : _T_14256; // @[Mux.scala 46:16:@10820.4]
  assign _T_14259 = 6'h4 == _T_11317_41; // @[Mux.scala 46:19:@10821.4]
  assign _T_14260 = _T_14259 ? _T_10366_3 : _T_14258; // @[Mux.scala 46:16:@10822.4]
  assign _T_14261 = 6'h3 == _T_11317_41; // @[Mux.scala 46:19:@10823.4]
  assign _T_14262 = _T_14261 ? _T_10366_2 : _T_14260; // @[Mux.scala 46:16:@10824.4]
  assign _T_14263 = 6'h2 == _T_11317_41; // @[Mux.scala 46:19:@10825.4]
  assign _T_14264 = _T_14263 ? _T_10366_1 : _T_14262; // @[Mux.scala 46:16:@10826.4]
  assign _T_14265 = 6'h1 == _T_11317_41; // @[Mux.scala 46:19:@10827.4]
  assign _T_14266 = _T_14265 ? _T_10366_0 : _T_14264; // @[Mux.scala 46:16:@10828.4]
  assign _T_14311 = 6'h2b == _T_11317_42; // @[Mux.scala 46:19:@10830.4]
  assign _T_14312 = _T_14311 ? _T_10366_42 : 8'h0; // @[Mux.scala 46:16:@10831.4]
  assign _T_14313 = 6'h2a == _T_11317_42; // @[Mux.scala 46:19:@10832.4]
  assign _T_14314 = _T_14313 ? _T_10366_41 : _T_14312; // @[Mux.scala 46:16:@10833.4]
  assign _T_14315 = 6'h29 == _T_11317_42; // @[Mux.scala 46:19:@10834.4]
  assign _T_14316 = _T_14315 ? _T_10366_40 : _T_14314; // @[Mux.scala 46:16:@10835.4]
  assign _T_14317 = 6'h28 == _T_11317_42; // @[Mux.scala 46:19:@10836.4]
  assign _T_14318 = _T_14317 ? _T_10366_39 : _T_14316; // @[Mux.scala 46:16:@10837.4]
  assign _T_14319 = 6'h27 == _T_11317_42; // @[Mux.scala 46:19:@10838.4]
  assign _T_14320 = _T_14319 ? _T_10366_38 : _T_14318; // @[Mux.scala 46:16:@10839.4]
  assign _T_14321 = 6'h26 == _T_11317_42; // @[Mux.scala 46:19:@10840.4]
  assign _T_14322 = _T_14321 ? _T_10366_37 : _T_14320; // @[Mux.scala 46:16:@10841.4]
  assign _T_14323 = 6'h25 == _T_11317_42; // @[Mux.scala 46:19:@10842.4]
  assign _T_14324 = _T_14323 ? _T_10366_36 : _T_14322; // @[Mux.scala 46:16:@10843.4]
  assign _T_14325 = 6'h24 == _T_11317_42; // @[Mux.scala 46:19:@10844.4]
  assign _T_14326 = _T_14325 ? _T_10366_35 : _T_14324; // @[Mux.scala 46:16:@10845.4]
  assign _T_14327 = 6'h23 == _T_11317_42; // @[Mux.scala 46:19:@10846.4]
  assign _T_14328 = _T_14327 ? _T_10366_34 : _T_14326; // @[Mux.scala 46:16:@10847.4]
  assign _T_14329 = 6'h22 == _T_11317_42; // @[Mux.scala 46:19:@10848.4]
  assign _T_14330 = _T_14329 ? _T_10366_33 : _T_14328; // @[Mux.scala 46:16:@10849.4]
  assign _T_14331 = 6'h21 == _T_11317_42; // @[Mux.scala 46:19:@10850.4]
  assign _T_14332 = _T_14331 ? _T_10366_32 : _T_14330; // @[Mux.scala 46:16:@10851.4]
  assign _T_14333 = 6'h20 == _T_11317_42; // @[Mux.scala 46:19:@10852.4]
  assign _T_14334 = _T_14333 ? _T_10366_31 : _T_14332; // @[Mux.scala 46:16:@10853.4]
  assign _T_14335 = 6'h1f == _T_11317_42; // @[Mux.scala 46:19:@10854.4]
  assign _T_14336 = _T_14335 ? _T_10366_30 : _T_14334; // @[Mux.scala 46:16:@10855.4]
  assign _T_14337 = 6'h1e == _T_11317_42; // @[Mux.scala 46:19:@10856.4]
  assign _T_14338 = _T_14337 ? _T_10366_29 : _T_14336; // @[Mux.scala 46:16:@10857.4]
  assign _T_14339 = 6'h1d == _T_11317_42; // @[Mux.scala 46:19:@10858.4]
  assign _T_14340 = _T_14339 ? _T_10366_28 : _T_14338; // @[Mux.scala 46:16:@10859.4]
  assign _T_14341 = 6'h1c == _T_11317_42; // @[Mux.scala 46:19:@10860.4]
  assign _T_14342 = _T_14341 ? _T_10366_27 : _T_14340; // @[Mux.scala 46:16:@10861.4]
  assign _T_14343 = 6'h1b == _T_11317_42; // @[Mux.scala 46:19:@10862.4]
  assign _T_14344 = _T_14343 ? _T_10366_26 : _T_14342; // @[Mux.scala 46:16:@10863.4]
  assign _T_14345 = 6'h1a == _T_11317_42; // @[Mux.scala 46:19:@10864.4]
  assign _T_14346 = _T_14345 ? _T_10366_25 : _T_14344; // @[Mux.scala 46:16:@10865.4]
  assign _T_14347 = 6'h19 == _T_11317_42; // @[Mux.scala 46:19:@10866.4]
  assign _T_14348 = _T_14347 ? _T_10366_24 : _T_14346; // @[Mux.scala 46:16:@10867.4]
  assign _T_14349 = 6'h18 == _T_11317_42; // @[Mux.scala 46:19:@10868.4]
  assign _T_14350 = _T_14349 ? _T_10366_23 : _T_14348; // @[Mux.scala 46:16:@10869.4]
  assign _T_14351 = 6'h17 == _T_11317_42; // @[Mux.scala 46:19:@10870.4]
  assign _T_14352 = _T_14351 ? _T_10366_22 : _T_14350; // @[Mux.scala 46:16:@10871.4]
  assign _T_14353 = 6'h16 == _T_11317_42; // @[Mux.scala 46:19:@10872.4]
  assign _T_14354 = _T_14353 ? _T_10366_21 : _T_14352; // @[Mux.scala 46:16:@10873.4]
  assign _T_14355 = 6'h15 == _T_11317_42; // @[Mux.scala 46:19:@10874.4]
  assign _T_14356 = _T_14355 ? _T_10366_20 : _T_14354; // @[Mux.scala 46:16:@10875.4]
  assign _T_14357 = 6'h14 == _T_11317_42; // @[Mux.scala 46:19:@10876.4]
  assign _T_14358 = _T_14357 ? _T_10366_19 : _T_14356; // @[Mux.scala 46:16:@10877.4]
  assign _T_14359 = 6'h13 == _T_11317_42; // @[Mux.scala 46:19:@10878.4]
  assign _T_14360 = _T_14359 ? _T_10366_18 : _T_14358; // @[Mux.scala 46:16:@10879.4]
  assign _T_14361 = 6'h12 == _T_11317_42; // @[Mux.scala 46:19:@10880.4]
  assign _T_14362 = _T_14361 ? _T_10366_17 : _T_14360; // @[Mux.scala 46:16:@10881.4]
  assign _T_14363 = 6'h11 == _T_11317_42; // @[Mux.scala 46:19:@10882.4]
  assign _T_14364 = _T_14363 ? _T_10366_16 : _T_14362; // @[Mux.scala 46:16:@10883.4]
  assign _T_14365 = 6'h10 == _T_11317_42; // @[Mux.scala 46:19:@10884.4]
  assign _T_14366 = _T_14365 ? _T_10366_15 : _T_14364; // @[Mux.scala 46:16:@10885.4]
  assign _T_14367 = 6'hf == _T_11317_42; // @[Mux.scala 46:19:@10886.4]
  assign _T_14368 = _T_14367 ? _T_10366_14 : _T_14366; // @[Mux.scala 46:16:@10887.4]
  assign _T_14369 = 6'he == _T_11317_42; // @[Mux.scala 46:19:@10888.4]
  assign _T_14370 = _T_14369 ? _T_10366_13 : _T_14368; // @[Mux.scala 46:16:@10889.4]
  assign _T_14371 = 6'hd == _T_11317_42; // @[Mux.scala 46:19:@10890.4]
  assign _T_14372 = _T_14371 ? _T_10366_12 : _T_14370; // @[Mux.scala 46:16:@10891.4]
  assign _T_14373 = 6'hc == _T_11317_42; // @[Mux.scala 46:19:@10892.4]
  assign _T_14374 = _T_14373 ? _T_10366_11 : _T_14372; // @[Mux.scala 46:16:@10893.4]
  assign _T_14375 = 6'hb == _T_11317_42; // @[Mux.scala 46:19:@10894.4]
  assign _T_14376 = _T_14375 ? _T_10366_10 : _T_14374; // @[Mux.scala 46:16:@10895.4]
  assign _T_14377 = 6'ha == _T_11317_42; // @[Mux.scala 46:19:@10896.4]
  assign _T_14378 = _T_14377 ? _T_10366_9 : _T_14376; // @[Mux.scala 46:16:@10897.4]
  assign _T_14379 = 6'h9 == _T_11317_42; // @[Mux.scala 46:19:@10898.4]
  assign _T_14380 = _T_14379 ? _T_10366_8 : _T_14378; // @[Mux.scala 46:16:@10899.4]
  assign _T_14381 = 6'h8 == _T_11317_42; // @[Mux.scala 46:19:@10900.4]
  assign _T_14382 = _T_14381 ? _T_10366_7 : _T_14380; // @[Mux.scala 46:16:@10901.4]
  assign _T_14383 = 6'h7 == _T_11317_42; // @[Mux.scala 46:19:@10902.4]
  assign _T_14384 = _T_14383 ? _T_10366_6 : _T_14382; // @[Mux.scala 46:16:@10903.4]
  assign _T_14385 = 6'h6 == _T_11317_42; // @[Mux.scala 46:19:@10904.4]
  assign _T_14386 = _T_14385 ? _T_10366_5 : _T_14384; // @[Mux.scala 46:16:@10905.4]
  assign _T_14387 = 6'h5 == _T_11317_42; // @[Mux.scala 46:19:@10906.4]
  assign _T_14388 = _T_14387 ? _T_10366_4 : _T_14386; // @[Mux.scala 46:16:@10907.4]
  assign _T_14389 = 6'h4 == _T_11317_42; // @[Mux.scala 46:19:@10908.4]
  assign _T_14390 = _T_14389 ? _T_10366_3 : _T_14388; // @[Mux.scala 46:16:@10909.4]
  assign _T_14391 = 6'h3 == _T_11317_42; // @[Mux.scala 46:19:@10910.4]
  assign _T_14392 = _T_14391 ? _T_10366_2 : _T_14390; // @[Mux.scala 46:16:@10911.4]
  assign _T_14393 = 6'h2 == _T_11317_42; // @[Mux.scala 46:19:@10912.4]
  assign _T_14394 = _T_14393 ? _T_10366_1 : _T_14392; // @[Mux.scala 46:16:@10913.4]
  assign _T_14395 = 6'h1 == _T_11317_42; // @[Mux.scala 46:19:@10914.4]
  assign _T_14396 = _T_14395 ? _T_10366_0 : _T_14394; // @[Mux.scala 46:16:@10915.4]
  assign _T_14442 = 6'h2c == _T_11317_43; // @[Mux.scala 46:19:@10917.4]
  assign _T_14443 = _T_14442 ? _T_10366_43 : 8'h0; // @[Mux.scala 46:16:@10918.4]
  assign _T_14444 = 6'h2b == _T_11317_43; // @[Mux.scala 46:19:@10919.4]
  assign _T_14445 = _T_14444 ? _T_10366_42 : _T_14443; // @[Mux.scala 46:16:@10920.4]
  assign _T_14446 = 6'h2a == _T_11317_43; // @[Mux.scala 46:19:@10921.4]
  assign _T_14447 = _T_14446 ? _T_10366_41 : _T_14445; // @[Mux.scala 46:16:@10922.4]
  assign _T_14448 = 6'h29 == _T_11317_43; // @[Mux.scala 46:19:@10923.4]
  assign _T_14449 = _T_14448 ? _T_10366_40 : _T_14447; // @[Mux.scala 46:16:@10924.4]
  assign _T_14450 = 6'h28 == _T_11317_43; // @[Mux.scala 46:19:@10925.4]
  assign _T_14451 = _T_14450 ? _T_10366_39 : _T_14449; // @[Mux.scala 46:16:@10926.4]
  assign _T_14452 = 6'h27 == _T_11317_43; // @[Mux.scala 46:19:@10927.4]
  assign _T_14453 = _T_14452 ? _T_10366_38 : _T_14451; // @[Mux.scala 46:16:@10928.4]
  assign _T_14454 = 6'h26 == _T_11317_43; // @[Mux.scala 46:19:@10929.4]
  assign _T_14455 = _T_14454 ? _T_10366_37 : _T_14453; // @[Mux.scala 46:16:@10930.4]
  assign _T_14456 = 6'h25 == _T_11317_43; // @[Mux.scala 46:19:@10931.4]
  assign _T_14457 = _T_14456 ? _T_10366_36 : _T_14455; // @[Mux.scala 46:16:@10932.4]
  assign _T_14458 = 6'h24 == _T_11317_43; // @[Mux.scala 46:19:@10933.4]
  assign _T_14459 = _T_14458 ? _T_10366_35 : _T_14457; // @[Mux.scala 46:16:@10934.4]
  assign _T_14460 = 6'h23 == _T_11317_43; // @[Mux.scala 46:19:@10935.4]
  assign _T_14461 = _T_14460 ? _T_10366_34 : _T_14459; // @[Mux.scala 46:16:@10936.4]
  assign _T_14462 = 6'h22 == _T_11317_43; // @[Mux.scala 46:19:@10937.4]
  assign _T_14463 = _T_14462 ? _T_10366_33 : _T_14461; // @[Mux.scala 46:16:@10938.4]
  assign _T_14464 = 6'h21 == _T_11317_43; // @[Mux.scala 46:19:@10939.4]
  assign _T_14465 = _T_14464 ? _T_10366_32 : _T_14463; // @[Mux.scala 46:16:@10940.4]
  assign _T_14466 = 6'h20 == _T_11317_43; // @[Mux.scala 46:19:@10941.4]
  assign _T_14467 = _T_14466 ? _T_10366_31 : _T_14465; // @[Mux.scala 46:16:@10942.4]
  assign _T_14468 = 6'h1f == _T_11317_43; // @[Mux.scala 46:19:@10943.4]
  assign _T_14469 = _T_14468 ? _T_10366_30 : _T_14467; // @[Mux.scala 46:16:@10944.4]
  assign _T_14470 = 6'h1e == _T_11317_43; // @[Mux.scala 46:19:@10945.4]
  assign _T_14471 = _T_14470 ? _T_10366_29 : _T_14469; // @[Mux.scala 46:16:@10946.4]
  assign _T_14472 = 6'h1d == _T_11317_43; // @[Mux.scala 46:19:@10947.4]
  assign _T_14473 = _T_14472 ? _T_10366_28 : _T_14471; // @[Mux.scala 46:16:@10948.4]
  assign _T_14474 = 6'h1c == _T_11317_43; // @[Mux.scala 46:19:@10949.4]
  assign _T_14475 = _T_14474 ? _T_10366_27 : _T_14473; // @[Mux.scala 46:16:@10950.4]
  assign _T_14476 = 6'h1b == _T_11317_43; // @[Mux.scala 46:19:@10951.4]
  assign _T_14477 = _T_14476 ? _T_10366_26 : _T_14475; // @[Mux.scala 46:16:@10952.4]
  assign _T_14478 = 6'h1a == _T_11317_43; // @[Mux.scala 46:19:@10953.4]
  assign _T_14479 = _T_14478 ? _T_10366_25 : _T_14477; // @[Mux.scala 46:16:@10954.4]
  assign _T_14480 = 6'h19 == _T_11317_43; // @[Mux.scala 46:19:@10955.4]
  assign _T_14481 = _T_14480 ? _T_10366_24 : _T_14479; // @[Mux.scala 46:16:@10956.4]
  assign _T_14482 = 6'h18 == _T_11317_43; // @[Mux.scala 46:19:@10957.4]
  assign _T_14483 = _T_14482 ? _T_10366_23 : _T_14481; // @[Mux.scala 46:16:@10958.4]
  assign _T_14484 = 6'h17 == _T_11317_43; // @[Mux.scala 46:19:@10959.4]
  assign _T_14485 = _T_14484 ? _T_10366_22 : _T_14483; // @[Mux.scala 46:16:@10960.4]
  assign _T_14486 = 6'h16 == _T_11317_43; // @[Mux.scala 46:19:@10961.4]
  assign _T_14487 = _T_14486 ? _T_10366_21 : _T_14485; // @[Mux.scala 46:16:@10962.4]
  assign _T_14488 = 6'h15 == _T_11317_43; // @[Mux.scala 46:19:@10963.4]
  assign _T_14489 = _T_14488 ? _T_10366_20 : _T_14487; // @[Mux.scala 46:16:@10964.4]
  assign _T_14490 = 6'h14 == _T_11317_43; // @[Mux.scala 46:19:@10965.4]
  assign _T_14491 = _T_14490 ? _T_10366_19 : _T_14489; // @[Mux.scala 46:16:@10966.4]
  assign _T_14492 = 6'h13 == _T_11317_43; // @[Mux.scala 46:19:@10967.4]
  assign _T_14493 = _T_14492 ? _T_10366_18 : _T_14491; // @[Mux.scala 46:16:@10968.4]
  assign _T_14494 = 6'h12 == _T_11317_43; // @[Mux.scala 46:19:@10969.4]
  assign _T_14495 = _T_14494 ? _T_10366_17 : _T_14493; // @[Mux.scala 46:16:@10970.4]
  assign _T_14496 = 6'h11 == _T_11317_43; // @[Mux.scala 46:19:@10971.4]
  assign _T_14497 = _T_14496 ? _T_10366_16 : _T_14495; // @[Mux.scala 46:16:@10972.4]
  assign _T_14498 = 6'h10 == _T_11317_43; // @[Mux.scala 46:19:@10973.4]
  assign _T_14499 = _T_14498 ? _T_10366_15 : _T_14497; // @[Mux.scala 46:16:@10974.4]
  assign _T_14500 = 6'hf == _T_11317_43; // @[Mux.scala 46:19:@10975.4]
  assign _T_14501 = _T_14500 ? _T_10366_14 : _T_14499; // @[Mux.scala 46:16:@10976.4]
  assign _T_14502 = 6'he == _T_11317_43; // @[Mux.scala 46:19:@10977.4]
  assign _T_14503 = _T_14502 ? _T_10366_13 : _T_14501; // @[Mux.scala 46:16:@10978.4]
  assign _T_14504 = 6'hd == _T_11317_43; // @[Mux.scala 46:19:@10979.4]
  assign _T_14505 = _T_14504 ? _T_10366_12 : _T_14503; // @[Mux.scala 46:16:@10980.4]
  assign _T_14506 = 6'hc == _T_11317_43; // @[Mux.scala 46:19:@10981.4]
  assign _T_14507 = _T_14506 ? _T_10366_11 : _T_14505; // @[Mux.scala 46:16:@10982.4]
  assign _T_14508 = 6'hb == _T_11317_43; // @[Mux.scala 46:19:@10983.4]
  assign _T_14509 = _T_14508 ? _T_10366_10 : _T_14507; // @[Mux.scala 46:16:@10984.4]
  assign _T_14510 = 6'ha == _T_11317_43; // @[Mux.scala 46:19:@10985.4]
  assign _T_14511 = _T_14510 ? _T_10366_9 : _T_14509; // @[Mux.scala 46:16:@10986.4]
  assign _T_14512 = 6'h9 == _T_11317_43; // @[Mux.scala 46:19:@10987.4]
  assign _T_14513 = _T_14512 ? _T_10366_8 : _T_14511; // @[Mux.scala 46:16:@10988.4]
  assign _T_14514 = 6'h8 == _T_11317_43; // @[Mux.scala 46:19:@10989.4]
  assign _T_14515 = _T_14514 ? _T_10366_7 : _T_14513; // @[Mux.scala 46:16:@10990.4]
  assign _T_14516 = 6'h7 == _T_11317_43; // @[Mux.scala 46:19:@10991.4]
  assign _T_14517 = _T_14516 ? _T_10366_6 : _T_14515; // @[Mux.scala 46:16:@10992.4]
  assign _T_14518 = 6'h6 == _T_11317_43; // @[Mux.scala 46:19:@10993.4]
  assign _T_14519 = _T_14518 ? _T_10366_5 : _T_14517; // @[Mux.scala 46:16:@10994.4]
  assign _T_14520 = 6'h5 == _T_11317_43; // @[Mux.scala 46:19:@10995.4]
  assign _T_14521 = _T_14520 ? _T_10366_4 : _T_14519; // @[Mux.scala 46:16:@10996.4]
  assign _T_14522 = 6'h4 == _T_11317_43; // @[Mux.scala 46:19:@10997.4]
  assign _T_14523 = _T_14522 ? _T_10366_3 : _T_14521; // @[Mux.scala 46:16:@10998.4]
  assign _T_14524 = 6'h3 == _T_11317_43; // @[Mux.scala 46:19:@10999.4]
  assign _T_14525 = _T_14524 ? _T_10366_2 : _T_14523; // @[Mux.scala 46:16:@11000.4]
  assign _T_14526 = 6'h2 == _T_11317_43; // @[Mux.scala 46:19:@11001.4]
  assign _T_14527 = _T_14526 ? _T_10366_1 : _T_14525; // @[Mux.scala 46:16:@11002.4]
  assign _T_14528 = 6'h1 == _T_11317_43; // @[Mux.scala 46:19:@11003.4]
  assign _T_14529 = _T_14528 ? _T_10366_0 : _T_14527; // @[Mux.scala 46:16:@11004.4]
  assign _T_14576 = 6'h2d == _T_11317_44; // @[Mux.scala 46:19:@11006.4]
  assign _T_14577 = _T_14576 ? _T_10366_44 : 8'h0; // @[Mux.scala 46:16:@11007.4]
  assign _T_14578 = 6'h2c == _T_11317_44; // @[Mux.scala 46:19:@11008.4]
  assign _T_14579 = _T_14578 ? _T_10366_43 : _T_14577; // @[Mux.scala 46:16:@11009.4]
  assign _T_14580 = 6'h2b == _T_11317_44; // @[Mux.scala 46:19:@11010.4]
  assign _T_14581 = _T_14580 ? _T_10366_42 : _T_14579; // @[Mux.scala 46:16:@11011.4]
  assign _T_14582 = 6'h2a == _T_11317_44; // @[Mux.scala 46:19:@11012.4]
  assign _T_14583 = _T_14582 ? _T_10366_41 : _T_14581; // @[Mux.scala 46:16:@11013.4]
  assign _T_14584 = 6'h29 == _T_11317_44; // @[Mux.scala 46:19:@11014.4]
  assign _T_14585 = _T_14584 ? _T_10366_40 : _T_14583; // @[Mux.scala 46:16:@11015.4]
  assign _T_14586 = 6'h28 == _T_11317_44; // @[Mux.scala 46:19:@11016.4]
  assign _T_14587 = _T_14586 ? _T_10366_39 : _T_14585; // @[Mux.scala 46:16:@11017.4]
  assign _T_14588 = 6'h27 == _T_11317_44; // @[Mux.scala 46:19:@11018.4]
  assign _T_14589 = _T_14588 ? _T_10366_38 : _T_14587; // @[Mux.scala 46:16:@11019.4]
  assign _T_14590 = 6'h26 == _T_11317_44; // @[Mux.scala 46:19:@11020.4]
  assign _T_14591 = _T_14590 ? _T_10366_37 : _T_14589; // @[Mux.scala 46:16:@11021.4]
  assign _T_14592 = 6'h25 == _T_11317_44; // @[Mux.scala 46:19:@11022.4]
  assign _T_14593 = _T_14592 ? _T_10366_36 : _T_14591; // @[Mux.scala 46:16:@11023.4]
  assign _T_14594 = 6'h24 == _T_11317_44; // @[Mux.scala 46:19:@11024.4]
  assign _T_14595 = _T_14594 ? _T_10366_35 : _T_14593; // @[Mux.scala 46:16:@11025.4]
  assign _T_14596 = 6'h23 == _T_11317_44; // @[Mux.scala 46:19:@11026.4]
  assign _T_14597 = _T_14596 ? _T_10366_34 : _T_14595; // @[Mux.scala 46:16:@11027.4]
  assign _T_14598 = 6'h22 == _T_11317_44; // @[Mux.scala 46:19:@11028.4]
  assign _T_14599 = _T_14598 ? _T_10366_33 : _T_14597; // @[Mux.scala 46:16:@11029.4]
  assign _T_14600 = 6'h21 == _T_11317_44; // @[Mux.scala 46:19:@11030.4]
  assign _T_14601 = _T_14600 ? _T_10366_32 : _T_14599; // @[Mux.scala 46:16:@11031.4]
  assign _T_14602 = 6'h20 == _T_11317_44; // @[Mux.scala 46:19:@11032.4]
  assign _T_14603 = _T_14602 ? _T_10366_31 : _T_14601; // @[Mux.scala 46:16:@11033.4]
  assign _T_14604 = 6'h1f == _T_11317_44; // @[Mux.scala 46:19:@11034.4]
  assign _T_14605 = _T_14604 ? _T_10366_30 : _T_14603; // @[Mux.scala 46:16:@11035.4]
  assign _T_14606 = 6'h1e == _T_11317_44; // @[Mux.scala 46:19:@11036.4]
  assign _T_14607 = _T_14606 ? _T_10366_29 : _T_14605; // @[Mux.scala 46:16:@11037.4]
  assign _T_14608 = 6'h1d == _T_11317_44; // @[Mux.scala 46:19:@11038.4]
  assign _T_14609 = _T_14608 ? _T_10366_28 : _T_14607; // @[Mux.scala 46:16:@11039.4]
  assign _T_14610 = 6'h1c == _T_11317_44; // @[Mux.scala 46:19:@11040.4]
  assign _T_14611 = _T_14610 ? _T_10366_27 : _T_14609; // @[Mux.scala 46:16:@11041.4]
  assign _T_14612 = 6'h1b == _T_11317_44; // @[Mux.scala 46:19:@11042.4]
  assign _T_14613 = _T_14612 ? _T_10366_26 : _T_14611; // @[Mux.scala 46:16:@11043.4]
  assign _T_14614 = 6'h1a == _T_11317_44; // @[Mux.scala 46:19:@11044.4]
  assign _T_14615 = _T_14614 ? _T_10366_25 : _T_14613; // @[Mux.scala 46:16:@11045.4]
  assign _T_14616 = 6'h19 == _T_11317_44; // @[Mux.scala 46:19:@11046.4]
  assign _T_14617 = _T_14616 ? _T_10366_24 : _T_14615; // @[Mux.scala 46:16:@11047.4]
  assign _T_14618 = 6'h18 == _T_11317_44; // @[Mux.scala 46:19:@11048.4]
  assign _T_14619 = _T_14618 ? _T_10366_23 : _T_14617; // @[Mux.scala 46:16:@11049.4]
  assign _T_14620 = 6'h17 == _T_11317_44; // @[Mux.scala 46:19:@11050.4]
  assign _T_14621 = _T_14620 ? _T_10366_22 : _T_14619; // @[Mux.scala 46:16:@11051.4]
  assign _T_14622 = 6'h16 == _T_11317_44; // @[Mux.scala 46:19:@11052.4]
  assign _T_14623 = _T_14622 ? _T_10366_21 : _T_14621; // @[Mux.scala 46:16:@11053.4]
  assign _T_14624 = 6'h15 == _T_11317_44; // @[Mux.scala 46:19:@11054.4]
  assign _T_14625 = _T_14624 ? _T_10366_20 : _T_14623; // @[Mux.scala 46:16:@11055.4]
  assign _T_14626 = 6'h14 == _T_11317_44; // @[Mux.scala 46:19:@11056.4]
  assign _T_14627 = _T_14626 ? _T_10366_19 : _T_14625; // @[Mux.scala 46:16:@11057.4]
  assign _T_14628 = 6'h13 == _T_11317_44; // @[Mux.scala 46:19:@11058.4]
  assign _T_14629 = _T_14628 ? _T_10366_18 : _T_14627; // @[Mux.scala 46:16:@11059.4]
  assign _T_14630 = 6'h12 == _T_11317_44; // @[Mux.scala 46:19:@11060.4]
  assign _T_14631 = _T_14630 ? _T_10366_17 : _T_14629; // @[Mux.scala 46:16:@11061.4]
  assign _T_14632 = 6'h11 == _T_11317_44; // @[Mux.scala 46:19:@11062.4]
  assign _T_14633 = _T_14632 ? _T_10366_16 : _T_14631; // @[Mux.scala 46:16:@11063.4]
  assign _T_14634 = 6'h10 == _T_11317_44; // @[Mux.scala 46:19:@11064.4]
  assign _T_14635 = _T_14634 ? _T_10366_15 : _T_14633; // @[Mux.scala 46:16:@11065.4]
  assign _T_14636 = 6'hf == _T_11317_44; // @[Mux.scala 46:19:@11066.4]
  assign _T_14637 = _T_14636 ? _T_10366_14 : _T_14635; // @[Mux.scala 46:16:@11067.4]
  assign _T_14638 = 6'he == _T_11317_44; // @[Mux.scala 46:19:@11068.4]
  assign _T_14639 = _T_14638 ? _T_10366_13 : _T_14637; // @[Mux.scala 46:16:@11069.4]
  assign _T_14640 = 6'hd == _T_11317_44; // @[Mux.scala 46:19:@11070.4]
  assign _T_14641 = _T_14640 ? _T_10366_12 : _T_14639; // @[Mux.scala 46:16:@11071.4]
  assign _T_14642 = 6'hc == _T_11317_44; // @[Mux.scala 46:19:@11072.4]
  assign _T_14643 = _T_14642 ? _T_10366_11 : _T_14641; // @[Mux.scala 46:16:@11073.4]
  assign _T_14644 = 6'hb == _T_11317_44; // @[Mux.scala 46:19:@11074.4]
  assign _T_14645 = _T_14644 ? _T_10366_10 : _T_14643; // @[Mux.scala 46:16:@11075.4]
  assign _T_14646 = 6'ha == _T_11317_44; // @[Mux.scala 46:19:@11076.4]
  assign _T_14647 = _T_14646 ? _T_10366_9 : _T_14645; // @[Mux.scala 46:16:@11077.4]
  assign _T_14648 = 6'h9 == _T_11317_44; // @[Mux.scala 46:19:@11078.4]
  assign _T_14649 = _T_14648 ? _T_10366_8 : _T_14647; // @[Mux.scala 46:16:@11079.4]
  assign _T_14650 = 6'h8 == _T_11317_44; // @[Mux.scala 46:19:@11080.4]
  assign _T_14651 = _T_14650 ? _T_10366_7 : _T_14649; // @[Mux.scala 46:16:@11081.4]
  assign _T_14652 = 6'h7 == _T_11317_44; // @[Mux.scala 46:19:@11082.4]
  assign _T_14653 = _T_14652 ? _T_10366_6 : _T_14651; // @[Mux.scala 46:16:@11083.4]
  assign _T_14654 = 6'h6 == _T_11317_44; // @[Mux.scala 46:19:@11084.4]
  assign _T_14655 = _T_14654 ? _T_10366_5 : _T_14653; // @[Mux.scala 46:16:@11085.4]
  assign _T_14656 = 6'h5 == _T_11317_44; // @[Mux.scala 46:19:@11086.4]
  assign _T_14657 = _T_14656 ? _T_10366_4 : _T_14655; // @[Mux.scala 46:16:@11087.4]
  assign _T_14658 = 6'h4 == _T_11317_44; // @[Mux.scala 46:19:@11088.4]
  assign _T_14659 = _T_14658 ? _T_10366_3 : _T_14657; // @[Mux.scala 46:16:@11089.4]
  assign _T_14660 = 6'h3 == _T_11317_44; // @[Mux.scala 46:19:@11090.4]
  assign _T_14661 = _T_14660 ? _T_10366_2 : _T_14659; // @[Mux.scala 46:16:@11091.4]
  assign _T_14662 = 6'h2 == _T_11317_44; // @[Mux.scala 46:19:@11092.4]
  assign _T_14663 = _T_14662 ? _T_10366_1 : _T_14661; // @[Mux.scala 46:16:@11093.4]
  assign _T_14664 = 6'h1 == _T_11317_44; // @[Mux.scala 46:19:@11094.4]
  assign _T_14665 = _T_14664 ? _T_10366_0 : _T_14663; // @[Mux.scala 46:16:@11095.4]
  assign _T_14713 = 6'h2e == _T_11317_45; // @[Mux.scala 46:19:@11097.4]
  assign _T_14714 = _T_14713 ? _T_10366_45 : 8'h0; // @[Mux.scala 46:16:@11098.4]
  assign _T_14715 = 6'h2d == _T_11317_45; // @[Mux.scala 46:19:@11099.4]
  assign _T_14716 = _T_14715 ? _T_10366_44 : _T_14714; // @[Mux.scala 46:16:@11100.4]
  assign _T_14717 = 6'h2c == _T_11317_45; // @[Mux.scala 46:19:@11101.4]
  assign _T_14718 = _T_14717 ? _T_10366_43 : _T_14716; // @[Mux.scala 46:16:@11102.4]
  assign _T_14719 = 6'h2b == _T_11317_45; // @[Mux.scala 46:19:@11103.4]
  assign _T_14720 = _T_14719 ? _T_10366_42 : _T_14718; // @[Mux.scala 46:16:@11104.4]
  assign _T_14721 = 6'h2a == _T_11317_45; // @[Mux.scala 46:19:@11105.4]
  assign _T_14722 = _T_14721 ? _T_10366_41 : _T_14720; // @[Mux.scala 46:16:@11106.4]
  assign _T_14723 = 6'h29 == _T_11317_45; // @[Mux.scala 46:19:@11107.4]
  assign _T_14724 = _T_14723 ? _T_10366_40 : _T_14722; // @[Mux.scala 46:16:@11108.4]
  assign _T_14725 = 6'h28 == _T_11317_45; // @[Mux.scala 46:19:@11109.4]
  assign _T_14726 = _T_14725 ? _T_10366_39 : _T_14724; // @[Mux.scala 46:16:@11110.4]
  assign _T_14727 = 6'h27 == _T_11317_45; // @[Mux.scala 46:19:@11111.4]
  assign _T_14728 = _T_14727 ? _T_10366_38 : _T_14726; // @[Mux.scala 46:16:@11112.4]
  assign _T_14729 = 6'h26 == _T_11317_45; // @[Mux.scala 46:19:@11113.4]
  assign _T_14730 = _T_14729 ? _T_10366_37 : _T_14728; // @[Mux.scala 46:16:@11114.4]
  assign _T_14731 = 6'h25 == _T_11317_45; // @[Mux.scala 46:19:@11115.4]
  assign _T_14732 = _T_14731 ? _T_10366_36 : _T_14730; // @[Mux.scala 46:16:@11116.4]
  assign _T_14733 = 6'h24 == _T_11317_45; // @[Mux.scala 46:19:@11117.4]
  assign _T_14734 = _T_14733 ? _T_10366_35 : _T_14732; // @[Mux.scala 46:16:@11118.4]
  assign _T_14735 = 6'h23 == _T_11317_45; // @[Mux.scala 46:19:@11119.4]
  assign _T_14736 = _T_14735 ? _T_10366_34 : _T_14734; // @[Mux.scala 46:16:@11120.4]
  assign _T_14737 = 6'h22 == _T_11317_45; // @[Mux.scala 46:19:@11121.4]
  assign _T_14738 = _T_14737 ? _T_10366_33 : _T_14736; // @[Mux.scala 46:16:@11122.4]
  assign _T_14739 = 6'h21 == _T_11317_45; // @[Mux.scala 46:19:@11123.4]
  assign _T_14740 = _T_14739 ? _T_10366_32 : _T_14738; // @[Mux.scala 46:16:@11124.4]
  assign _T_14741 = 6'h20 == _T_11317_45; // @[Mux.scala 46:19:@11125.4]
  assign _T_14742 = _T_14741 ? _T_10366_31 : _T_14740; // @[Mux.scala 46:16:@11126.4]
  assign _T_14743 = 6'h1f == _T_11317_45; // @[Mux.scala 46:19:@11127.4]
  assign _T_14744 = _T_14743 ? _T_10366_30 : _T_14742; // @[Mux.scala 46:16:@11128.4]
  assign _T_14745 = 6'h1e == _T_11317_45; // @[Mux.scala 46:19:@11129.4]
  assign _T_14746 = _T_14745 ? _T_10366_29 : _T_14744; // @[Mux.scala 46:16:@11130.4]
  assign _T_14747 = 6'h1d == _T_11317_45; // @[Mux.scala 46:19:@11131.4]
  assign _T_14748 = _T_14747 ? _T_10366_28 : _T_14746; // @[Mux.scala 46:16:@11132.4]
  assign _T_14749 = 6'h1c == _T_11317_45; // @[Mux.scala 46:19:@11133.4]
  assign _T_14750 = _T_14749 ? _T_10366_27 : _T_14748; // @[Mux.scala 46:16:@11134.4]
  assign _T_14751 = 6'h1b == _T_11317_45; // @[Mux.scala 46:19:@11135.4]
  assign _T_14752 = _T_14751 ? _T_10366_26 : _T_14750; // @[Mux.scala 46:16:@11136.4]
  assign _T_14753 = 6'h1a == _T_11317_45; // @[Mux.scala 46:19:@11137.4]
  assign _T_14754 = _T_14753 ? _T_10366_25 : _T_14752; // @[Mux.scala 46:16:@11138.4]
  assign _T_14755 = 6'h19 == _T_11317_45; // @[Mux.scala 46:19:@11139.4]
  assign _T_14756 = _T_14755 ? _T_10366_24 : _T_14754; // @[Mux.scala 46:16:@11140.4]
  assign _T_14757 = 6'h18 == _T_11317_45; // @[Mux.scala 46:19:@11141.4]
  assign _T_14758 = _T_14757 ? _T_10366_23 : _T_14756; // @[Mux.scala 46:16:@11142.4]
  assign _T_14759 = 6'h17 == _T_11317_45; // @[Mux.scala 46:19:@11143.4]
  assign _T_14760 = _T_14759 ? _T_10366_22 : _T_14758; // @[Mux.scala 46:16:@11144.4]
  assign _T_14761 = 6'h16 == _T_11317_45; // @[Mux.scala 46:19:@11145.4]
  assign _T_14762 = _T_14761 ? _T_10366_21 : _T_14760; // @[Mux.scala 46:16:@11146.4]
  assign _T_14763 = 6'h15 == _T_11317_45; // @[Mux.scala 46:19:@11147.4]
  assign _T_14764 = _T_14763 ? _T_10366_20 : _T_14762; // @[Mux.scala 46:16:@11148.4]
  assign _T_14765 = 6'h14 == _T_11317_45; // @[Mux.scala 46:19:@11149.4]
  assign _T_14766 = _T_14765 ? _T_10366_19 : _T_14764; // @[Mux.scala 46:16:@11150.4]
  assign _T_14767 = 6'h13 == _T_11317_45; // @[Mux.scala 46:19:@11151.4]
  assign _T_14768 = _T_14767 ? _T_10366_18 : _T_14766; // @[Mux.scala 46:16:@11152.4]
  assign _T_14769 = 6'h12 == _T_11317_45; // @[Mux.scala 46:19:@11153.4]
  assign _T_14770 = _T_14769 ? _T_10366_17 : _T_14768; // @[Mux.scala 46:16:@11154.4]
  assign _T_14771 = 6'h11 == _T_11317_45; // @[Mux.scala 46:19:@11155.4]
  assign _T_14772 = _T_14771 ? _T_10366_16 : _T_14770; // @[Mux.scala 46:16:@11156.4]
  assign _T_14773 = 6'h10 == _T_11317_45; // @[Mux.scala 46:19:@11157.4]
  assign _T_14774 = _T_14773 ? _T_10366_15 : _T_14772; // @[Mux.scala 46:16:@11158.4]
  assign _T_14775 = 6'hf == _T_11317_45; // @[Mux.scala 46:19:@11159.4]
  assign _T_14776 = _T_14775 ? _T_10366_14 : _T_14774; // @[Mux.scala 46:16:@11160.4]
  assign _T_14777 = 6'he == _T_11317_45; // @[Mux.scala 46:19:@11161.4]
  assign _T_14778 = _T_14777 ? _T_10366_13 : _T_14776; // @[Mux.scala 46:16:@11162.4]
  assign _T_14779 = 6'hd == _T_11317_45; // @[Mux.scala 46:19:@11163.4]
  assign _T_14780 = _T_14779 ? _T_10366_12 : _T_14778; // @[Mux.scala 46:16:@11164.4]
  assign _T_14781 = 6'hc == _T_11317_45; // @[Mux.scala 46:19:@11165.4]
  assign _T_14782 = _T_14781 ? _T_10366_11 : _T_14780; // @[Mux.scala 46:16:@11166.4]
  assign _T_14783 = 6'hb == _T_11317_45; // @[Mux.scala 46:19:@11167.4]
  assign _T_14784 = _T_14783 ? _T_10366_10 : _T_14782; // @[Mux.scala 46:16:@11168.4]
  assign _T_14785 = 6'ha == _T_11317_45; // @[Mux.scala 46:19:@11169.4]
  assign _T_14786 = _T_14785 ? _T_10366_9 : _T_14784; // @[Mux.scala 46:16:@11170.4]
  assign _T_14787 = 6'h9 == _T_11317_45; // @[Mux.scala 46:19:@11171.4]
  assign _T_14788 = _T_14787 ? _T_10366_8 : _T_14786; // @[Mux.scala 46:16:@11172.4]
  assign _T_14789 = 6'h8 == _T_11317_45; // @[Mux.scala 46:19:@11173.4]
  assign _T_14790 = _T_14789 ? _T_10366_7 : _T_14788; // @[Mux.scala 46:16:@11174.4]
  assign _T_14791 = 6'h7 == _T_11317_45; // @[Mux.scala 46:19:@11175.4]
  assign _T_14792 = _T_14791 ? _T_10366_6 : _T_14790; // @[Mux.scala 46:16:@11176.4]
  assign _T_14793 = 6'h6 == _T_11317_45; // @[Mux.scala 46:19:@11177.4]
  assign _T_14794 = _T_14793 ? _T_10366_5 : _T_14792; // @[Mux.scala 46:16:@11178.4]
  assign _T_14795 = 6'h5 == _T_11317_45; // @[Mux.scala 46:19:@11179.4]
  assign _T_14796 = _T_14795 ? _T_10366_4 : _T_14794; // @[Mux.scala 46:16:@11180.4]
  assign _T_14797 = 6'h4 == _T_11317_45; // @[Mux.scala 46:19:@11181.4]
  assign _T_14798 = _T_14797 ? _T_10366_3 : _T_14796; // @[Mux.scala 46:16:@11182.4]
  assign _T_14799 = 6'h3 == _T_11317_45; // @[Mux.scala 46:19:@11183.4]
  assign _T_14800 = _T_14799 ? _T_10366_2 : _T_14798; // @[Mux.scala 46:16:@11184.4]
  assign _T_14801 = 6'h2 == _T_11317_45; // @[Mux.scala 46:19:@11185.4]
  assign _T_14802 = _T_14801 ? _T_10366_1 : _T_14800; // @[Mux.scala 46:16:@11186.4]
  assign _T_14803 = 6'h1 == _T_11317_45; // @[Mux.scala 46:19:@11187.4]
  assign _T_14804 = _T_14803 ? _T_10366_0 : _T_14802; // @[Mux.scala 46:16:@11188.4]
  assign _T_14853 = 6'h2f == _T_11317_46; // @[Mux.scala 46:19:@11190.4]
  assign _T_14854 = _T_14853 ? _T_10366_46 : 8'h0; // @[Mux.scala 46:16:@11191.4]
  assign _T_14855 = 6'h2e == _T_11317_46; // @[Mux.scala 46:19:@11192.4]
  assign _T_14856 = _T_14855 ? _T_10366_45 : _T_14854; // @[Mux.scala 46:16:@11193.4]
  assign _T_14857 = 6'h2d == _T_11317_46; // @[Mux.scala 46:19:@11194.4]
  assign _T_14858 = _T_14857 ? _T_10366_44 : _T_14856; // @[Mux.scala 46:16:@11195.4]
  assign _T_14859 = 6'h2c == _T_11317_46; // @[Mux.scala 46:19:@11196.4]
  assign _T_14860 = _T_14859 ? _T_10366_43 : _T_14858; // @[Mux.scala 46:16:@11197.4]
  assign _T_14861 = 6'h2b == _T_11317_46; // @[Mux.scala 46:19:@11198.4]
  assign _T_14862 = _T_14861 ? _T_10366_42 : _T_14860; // @[Mux.scala 46:16:@11199.4]
  assign _T_14863 = 6'h2a == _T_11317_46; // @[Mux.scala 46:19:@11200.4]
  assign _T_14864 = _T_14863 ? _T_10366_41 : _T_14862; // @[Mux.scala 46:16:@11201.4]
  assign _T_14865 = 6'h29 == _T_11317_46; // @[Mux.scala 46:19:@11202.4]
  assign _T_14866 = _T_14865 ? _T_10366_40 : _T_14864; // @[Mux.scala 46:16:@11203.4]
  assign _T_14867 = 6'h28 == _T_11317_46; // @[Mux.scala 46:19:@11204.4]
  assign _T_14868 = _T_14867 ? _T_10366_39 : _T_14866; // @[Mux.scala 46:16:@11205.4]
  assign _T_14869 = 6'h27 == _T_11317_46; // @[Mux.scala 46:19:@11206.4]
  assign _T_14870 = _T_14869 ? _T_10366_38 : _T_14868; // @[Mux.scala 46:16:@11207.4]
  assign _T_14871 = 6'h26 == _T_11317_46; // @[Mux.scala 46:19:@11208.4]
  assign _T_14872 = _T_14871 ? _T_10366_37 : _T_14870; // @[Mux.scala 46:16:@11209.4]
  assign _T_14873 = 6'h25 == _T_11317_46; // @[Mux.scala 46:19:@11210.4]
  assign _T_14874 = _T_14873 ? _T_10366_36 : _T_14872; // @[Mux.scala 46:16:@11211.4]
  assign _T_14875 = 6'h24 == _T_11317_46; // @[Mux.scala 46:19:@11212.4]
  assign _T_14876 = _T_14875 ? _T_10366_35 : _T_14874; // @[Mux.scala 46:16:@11213.4]
  assign _T_14877 = 6'h23 == _T_11317_46; // @[Mux.scala 46:19:@11214.4]
  assign _T_14878 = _T_14877 ? _T_10366_34 : _T_14876; // @[Mux.scala 46:16:@11215.4]
  assign _T_14879 = 6'h22 == _T_11317_46; // @[Mux.scala 46:19:@11216.4]
  assign _T_14880 = _T_14879 ? _T_10366_33 : _T_14878; // @[Mux.scala 46:16:@11217.4]
  assign _T_14881 = 6'h21 == _T_11317_46; // @[Mux.scala 46:19:@11218.4]
  assign _T_14882 = _T_14881 ? _T_10366_32 : _T_14880; // @[Mux.scala 46:16:@11219.4]
  assign _T_14883 = 6'h20 == _T_11317_46; // @[Mux.scala 46:19:@11220.4]
  assign _T_14884 = _T_14883 ? _T_10366_31 : _T_14882; // @[Mux.scala 46:16:@11221.4]
  assign _T_14885 = 6'h1f == _T_11317_46; // @[Mux.scala 46:19:@11222.4]
  assign _T_14886 = _T_14885 ? _T_10366_30 : _T_14884; // @[Mux.scala 46:16:@11223.4]
  assign _T_14887 = 6'h1e == _T_11317_46; // @[Mux.scala 46:19:@11224.4]
  assign _T_14888 = _T_14887 ? _T_10366_29 : _T_14886; // @[Mux.scala 46:16:@11225.4]
  assign _T_14889 = 6'h1d == _T_11317_46; // @[Mux.scala 46:19:@11226.4]
  assign _T_14890 = _T_14889 ? _T_10366_28 : _T_14888; // @[Mux.scala 46:16:@11227.4]
  assign _T_14891 = 6'h1c == _T_11317_46; // @[Mux.scala 46:19:@11228.4]
  assign _T_14892 = _T_14891 ? _T_10366_27 : _T_14890; // @[Mux.scala 46:16:@11229.4]
  assign _T_14893 = 6'h1b == _T_11317_46; // @[Mux.scala 46:19:@11230.4]
  assign _T_14894 = _T_14893 ? _T_10366_26 : _T_14892; // @[Mux.scala 46:16:@11231.4]
  assign _T_14895 = 6'h1a == _T_11317_46; // @[Mux.scala 46:19:@11232.4]
  assign _T_14896 = _T_14895 ? _T_10366_25 : _T_14894; // @[Mux.scala 46:16:@11233.4]
  assign _T_14897 = 6'h19 == _T_11317_46; // @[Mux.scala 46:19:@11234.4]
  assign _T_14898 = _T_14897 ? _T_10366_24 : _T_14896; // @[Mux.scala 46:16:@11235.4]
  assign _T_14899 = 6'h18 == _T_11317_46; // @[Mux.scala 46:19:@11236.4]
  assign _T_14900 = _T_14899 ? _T_10366_23 : _T_14898; // @[Mux.scala 46:16:@11237.4]
  assign _T_14901 = 6'h17 == _T_11317_46; // @[Mux.scala 46:19:@11238.4]
  assign _T_14902 = _T_14901 ? _T_10366_22 : _T_14900; // @[Mux.scala 46:16:@11239.4]
  assign _T_14903 = 6'h16 == _T_11317_46; // @[Mux.scala 46:19:@11240.4]
  assign _T_14904 = _T_14903 ? _T_10366_21 : _T_14902; // @[Mux.scala 46:16:@11241.4]
  assign _T_14905 = 6'h15 == _T_11317_46; // @[Mux.scala 46:19:@11242.4]
  assign _T_14906 = _T_14905 ? _T_10366_20 : _T_14904; // @[Mux.scala 46:16:@11243.4]
  assign _T_14907 = 6'h14 == _T_11317_46; // @[Mux.scala 46:19:@11244.4]
  assign _T_14908 = _T_14907 ? _T_10366_19 : _T_14906; // @[Mux.scala 46:16:@11245.4]
  assign _T_14909 = 6'h13 == _T_11317_46; // @[Mux.scala 46:19:@11246.4]
  assign _T_14910 = _T_14909 ? _T_10366_18 : _T_14908; // @[Mux.scala 46:16:@11247.4]
  assign _T_14911 = 6'h12 == _T_11317_46; // @[Mux.scala 46:19:@11248.4]
  assign _T_14912 = _T_14911 ? _T_10366_17 : _T_14910; // @[Mux.scala 46:16:@11249.4]
  assign _T_14913 = 6'h11 == _T_11317_46; // @[Mux.scala 46:19:@11250.4]
  assign _T_14914 = _T_14913 ? _T_10366_16 : _T_14912; // @[Mux.scala 46:16:@11251.4]
  assign _T_14915 = 6'h10 == _T_11317_46; // @[Mux.scala 46:19:@11252.4]
  assign _T_14916 = _T_14915 ? _T_10366_15 : _T_14914; // @[Mux.scala 46:16:@11253.4]
  assign _T_14917 = 6'hf == _T_11317_46; // @[Mux.scala 46:19:@11254.4]
  assign _T_14918 = _T_14917 ? _T_10366_14 : _T_14916; // @[Mux.scala 46:16:@11255.4]
  assign _T_14919 = 6'he == _T_11317_46; // @[Mux.scala 46:19:@11256.4]
  assign _T_14920 = _T_14919 ? _T_10366_13 : _T_14918; // @[Mux.scala 46:16:@11257.4]
  assign _T_14921 = 6'hd == _T_11317_46; // @[Mux.scala 46:19:@11258.4]
  assign _T_14922 = _T_14921 ? _T_10366_12 : _T_14920; // @[Mux.scala 46:16:@11259.4]
  assign _T_14923 = 6'hc == _T_11317_46; // @[Mux.scala 46:19:@11260.4]
  assign _T_14924 = _T_14923 ? _T_10366_11 : _T_14922; // @[Mux.scala 46:16:@11261.4]
  assign _T_14925 = 6'hb == _T_11317_46; // @[Mux.scala 46:19:@11262.4]
  assign _T_14926 = _T_14925 ? _T_10366_10 : _T_14924; // @[Mux.scala 46:16:@11263.4]
  assign _T_14927 = 6'ha == _T_11317_46; // @[Mux.scala 46:19:@11264.4]
  assign _T_14928 = _T_14927 ? _T_10366_9 : _T_14926; // @[Mux.scala 46:16:@11265.4]
  assign _T_14929 = 6'h9 == _T_11317_46; // @[Mux.scala 46:19:@11266.4]
  assign _T_14930 = _T_14929 ? _T_10366_8 : _T_14928; // @[Mux.scala 46:16:@11267.4]
  assign _T_14931 = 6'h8 == _T_11317_46; // @[Mux.scala 46:19:@11268.4]
  assign _T_14932 = _T_14931 ? _T_10366_7 : _T_14930; // @[Mux.scala 46:16:@11269.4]
  assign _T_14933 = 6'h7 == _T_11317_46; // @[Mux.scala 46:19:@11270.4]
  assign _T_14934 = _T_14933 ? _T_10366_6 : _T_14932; // @[Mux.scala 46:16:@11271.4]
  assign _T_14935 = 6'h6 == _T_11317_46; // @[Mux.scala 46:19:@11272.4]
  assign _T_14936 = _T_14935 ? _T_10366_5 : _T_14934; // @[Mux.scala 46:16:@11273.4]
  assign _T_14937 = 6'h5 == _T_11317_46; // @[Mux.scala 46:19:@11274.4]
  assign _T_14938 = _T_14937 ? _T_10366_4 : _T_14936; // @[Mux.scala 46:16:@11275.4]
  assign _T_14939 = 6'h4 == _T_11317_46; // @[Mux.scala 46:19:@11276.4]
  assign _T_14940 = _T_14939 ? _T_10366_3 : _T_14938; // @[Mux.scala 46:16:@11277.4]
  assign _T_14941 = 6'h3 == _T_11317_46; // @[Mux.scala 46:19:@11278.4]
  assign _T_14942 = _T_14941 ? _T_10366_2 : _T_14940; // @[Mux.scala 46:16:@11279.4]
  assign _T_14943 = 6'h2 == _T_11317_46; // @[Mux.scala 46:19:@11280.4]
  assign _T_14944 = _T_14943 ? _T_10366_1 : _T_14942; // @[Mux.scala 46:16:@11281.4]
  assign _T_14945 = 6'h1 == _T_11317_46; // @[Mux.scala 46:19:@11282.4]
  assign _T_14946 = _T_14945 ? _T_10366_0 : _T_14944; // @[Mux.scala 46:16:@11283.4]
  assign _T_14996 = 6'h30 == _T_11317_47; // @[Mux.scala 46:19:@11285.4]
  assign _T_14997 = _T_14996 ? _T_10366_47 : 8'h0; // @[Mux.scala 46:16:@11286.4]
  assign _T_14998 = 6'h2f == _T_11317_47; // @[Mux.scala 46:19:@11287.4]
  assign _T_14999 = _T_14998 ? _T_10366_46 : _T_14997; // @[Mux.scala 46:16:@11288.4]
  assign _T_15000 = 6'h2e == _T_11317_47; // @[Mux.scala 46:19:@11289.4]
  assign _T_15001 = _T_15000 ? _T_10366_45 : _T_14999; // @[Mux.scala 46:16:@11290.4]
  assign _T_15002 = 6'h2d == _T_11317_47; // @[Mux.scala 46:19:@11291.4]
  assign _T_15003 = _T_15002 ? _T_10366_44 : _T_15001; // @[Mux.scala 46:16:@11292.4]
  assign _T_15004 = 6'h2c == _T_11317_47; // @[Mux.scala 46:19:@11293.4]
  assign _T_15005 = _T_15004 ? _T_10366_43 : _T_15003; // @[Mux.scala 46:16:@11294.4]
  assign _T_15006 = 6'h2b == _T_11317_47; // @[Mux.scala 46:19:@11295.4]
  assign _T_15007 = _T_15006 ? _T_10366_42 : _T_15005; // @[Mux.scala 46:16:@11296.4]
  assign _T_15008 = 6'h2a == _T_11317_47; // @[Mux.scala 46:19:@11297.4]
  assign _T_15009 = _T_15008 ? _T_10366_41 : _T_15007; // @[Mux.scala 46:16:@11298.4]
  assign _T_15010 = 6'h29 == _T_11317_47; // @[Mux.scala 46:19:@11299.4]
  assign _T_15011 = _T_15010 ? _T_10366_40 : _T_15009; // @[Mux.scala 46:16:@11300.4]
  assign _T_15012 = 6'h28 == _T_11317_47; // @[Mux.scala 46:19:@11301.4]
  assign _T_15013 = _T_15012 ? _T_10366_39 : _T_15011; // @[Mux.scala 46:16:@11302.4]
  assign _T_15014 = 6'h27 == _T_11317_47; // @[Mux.scala 46:19:@11303.4]
  assign _T_15015 = _T_15014 ? _T_10366_38 : _T_15013; // @[Mux.scala 46:16:@11304.4]
  assign _T_15016 = 6'h26 == _T_11317_47; // @[Mux.scala 46:19:@11305.4]
  assign _T_15017 = _T_15016 ? _T_10366_37 : _T_15015; // @[Mux.scala 46:16:@11306.4]
  assign _T_15018 = 6'h25 == _T_11317_47; // @[Mux.scala 46:19:@11307.4]
  assign _T_15019 = _T_15018 ? _T_10366_36 : _T_15017; // @[Mux.scala 46:16:@11308.4]
  assign _T_15020 = 6'h24 == _T_11317_47; // @[Mux.scala 46:19:@11309.4]
  assign _T_15021 = _T_15020 ? _T_10366_35 : _T_15019; // @[Mux.scala 46:16:@11310.4]
  assign _T_15022 = 6'h23 == _T_11317_47; // @[Mux.scala 46:19:@11311.4]
  assign _T_15023 = _T_15022 ? _T_10366_34 : _T_15021; // @[Mux.scala 46:16:@11312.4]
  assign _T_15024 = 6'h22 == _T_11317_47; // @[Mux.scala 46:19:@11313.4]
  assign _T_15025 = _T_15024 ? _T_10366_33 : _T_15023; // @[Mux.scala 46:16:@11314.4]
  assign _T_15026 = 6'h21 == _T_11317_47; // @[Mux.scala 46:19:@11315.4]
  assign _T_15027 = _T_15026 ? _T_10366_32 : _T_15025; // @[Mux.scala 46:16:@11316.4]
  assign _T_15028 = 6'h20 == _T_11317_47; // @[Mux.scala 46:19:@11317.4]
  assign _T_15029 = _T_15028 ? _T_10366_31 : _T_15027; // @[Mux.scala 46:16:@11318.4]
  assign _T_15030 = 6'h1f == _T_11317_47; // @[Mux.scala 46:19:@11319.4]
  assign _T_15031 = _T_15030 ? _T_10366_30 : _T_15029; // @[Mux.scala 46:16:@11320.4]
  assign _T_15032 = 6'h1e == _T_11317_47; // @[Mux.scala 46:19:@11321.4]
  assign _T_15033 = _T_15032 ? _T_10366_29 : _T_15031; // @[Mux.scala 46:16:@11322.4]
  assign _T_15034 = 6'h1d == _T_11317_47; // @[Mux.scala 46:19:@11323.4]
  assign _T_15035 = _T_15034 ? _T_10366_28 : _T_15033; // @[Mux.scala 46:16:@11324.4]
  assign _T_15036 = 6'h1c == _T_11317_47; // @[Mux.scala 46:19:@11325.4]
  assign _T_15037 = _T_15036 ? _T_10366_27 : _T_15035; // @[Mux.scala 46:16:@11326.4]
  assign _T_15038 = 6'h1b == _T_11317_47; // @[Mux.scala 46:19:@11327.4]
  assign _T_15039 = _T_15038 ? _T_10366_26 : _T_15037; // @[Mux.scala 46:16:@11328.4]
  assign _T_15040 = 6'h1a == _T_11317_47; // @[Mux.scala 46:19:@11329.4]
  assign _T_15041 = _T_15040 ? _T_10366_25 : _T_15039; // @[Mux.scala 46:16:@11330.4]
  assign _T_15042 = 6'h19 == _T_11317_47; // @[Mux.scala 46:19:@11331.4]
  assign _T_15043 = _T_15042 ? _T_10366_24 : _T_15041; // @[Mux.scala 46:16:@11332.4]
  assign _T_15044 = 6'h18 == _T_11317_47; // @[Mux.scala 46:19:@11333.4]
  assign _T_15045 = _T_15044 ? _T_10366_23 : _T_15043; // @[Mux.scala 46:16:@11334.4]
  assign _T_15046 = 6'h17 == _T_11317_47; // @[Mux.scala 46:19:@11335.4]
  assign _T_15047 = _T_15046 ? _T_10366_22 : _T_15045; // @[Mux.scala 46:16:@11336.4]
  assign _T_15048 = 6'h16 == _T_11317_47; // @[Mux.scala 46:19:@11337.4]
  assign _T_15049 = _T_15048 ? _T_10366_21 : _T_15047; // @[Mux.scala 46:16:@11338.4]
  assign _T_15050 = 6'h15 == _T_11317_47; // @[Mux.scala 46:19:@11339.4]
  assign _T_15051 = _T_15050 ? _T_10366_20 : _T_15049; // @[Mux.scala 46:16:@11340.4]
  assign _T_15052 = 6'h14 == _T_11317_47; // @[Mux.scala 46:19:@11341.4]
  assign _T_15053 = _T_15052 ? _T_10366_19 : _T_15051; // @[Mux.scala 46:16:@11342.4]
  assign _T_15054 = 6'h13 == _T_11317_47; // @[Mux.scala 46:19:@11343.4]
  assign _T_15055 = _T_15054 ? _T_10366_18 : _T_15053; // @[Mux.scala 46:16:@11344.4]
  assign _T_15056 = 6'h12 == _T_11317_47; // @[Mux.scala 46:19:@11345.4]
  assign _T_15057 = _T_15056 ? _T_10366_17 : _T_15055; // @[Mux.scala 46:16:@11346.4]
  assign _T_15058 = 6'h11 == _T_11317_47; // @[Mux.scala 46:19:@11347.4]
  assign _T_15059 = _T_15058 ? _T_10366_16 : _T_15057; // @[Mux.scala 46:16:@11348.4]
  assign _T_15060 = 6'h10 == _T_11317_47; // @[Mux.scala 46:19:@11349.4]
  assign _T_15061 = _T_15060 ? _T_10366_15 : _T_15059; // @[Mux.scala 46:16:@11350.4]
  assign _T_15062 = 6'hf == _T_11317_47; // @[Mux.scala 46:19:@11351.4]
  assign _T_15063 = _T_15062 ? _T_10366_14 : _T_15061; // @[Mux.scala 46:16:@11352.4]
  assign _T_15064 = 6'he == _T_11317_47; // @[Mux.scala 46:19:@11353.4]
  assign _T_15065 = _T_15064 ? _T_10366_13 : _T_15063; // @[Mux.scala 46:16:@11354.4]
  assign _T_15066 = 6'hd == _T_11317_47; // @[Mux.scala 46:19:@11355.4]
  assign _T_15067 = _T_15066 ? _T_10366_12 : _T_15065; // @[Mux.scala 46:16:@11356.4]
  assign _T_15068 = 6'hc == _T_11317_47; // @[Mux.scala 46:19:@11357.4]
  assign _T_15069 = _T_15068 ? _T_10366_11 : _T_15067; // @[Mux.scala 46:16:@11358.4]
  assign _T_15070 = 6'hb == _T_11317_47; // @[Mux.scala 46:19:@11359.4]
  assign _T_15071 = _T_15070 ? _T_10366_10 : _T_15069; // @[Mux.scala 46:16:@11360.4]
  assign _T_15072 = 6'ha == _T_11317_47; // @[Mux.scala 46:19:@11361.4]
  assign _T_15073 = _T_15072 ? _T_10366_9 : _T_15071; // @[Mux.scala 46:16:@11362.4]
  assign _T_15074 = 6'h9 == _T_11317_47; // @[Mux.scala 46:19:@11363.4]
  assign _T_15075 = _T_15074 ? _T_10366_8 : _T_15073; // @[Mux.scala 46:16:@11364.4]
  assign _T_15076 = 6'h8 == _T_11317_47; // @[Mux.scala 46:19:@11365.4]
  assign _T_15077 = _T_15076 ? _T_10366_7 : _T_15075; // @[Mux.scala 46:16:@11366.4]
  assign _T_15078 = 6'h7 == _T_11317_47; // @[Mux.scala 46:19:@11367.4]
  assign _T_15079 = _T_15078 ? _T_10366_6 : _T_15077; // @[Mux.scala 46:16:@11368.4]
  assign _T_15080 = 6'h6 == _T_11317_47; // @[Mux.scala 46:19:@11369.4]
  assign _T_15081 = _T_15080 ? _T_10366_5 : _T_15079; // @[Mux.scala 46:16:@11370.4]
  assign _T_15082 = 6'h5 == _T_11317_47; // @[Mux.scala 46:19:@11371.4]
  assign _T_15083 = _T_15082 ? _T_10366_4 : _T_15081; // @[Mux.scala 46:16:@11372.4]
  assign _T_15084 = 6'h4 == _T_11317_47; // @[Mux.scala 46:19:@11373.4]
  assign _T_15085 = _T_15084 ? _T_10366_3 : _T_15083; // @[Mux.scala 46:16:@11374.4]
  assign _T_15086 = 6'h3 == _T_11317_47; // @[Mux.scala 46:19:@11375.4]
  assign _T_15087 = _T_15086 ? _T_10366_2 : _T_15085; // @[Mux.scala 46:16:@11376.4]
  assign _T_15088 = 6'h2 == _T_11317_47; // @[Mux.scala 46:19:@11377.4]
  assign _T_15089 = _T_15088 ? _T_10366_1 : _T_15087; // @[Mux.scala 46:16:@11378.4]
  assign _T_15090 = 6'h1 == _T_11317_47; // @[Mux.scala 46:19:@11379.4]
  assign _T_15091 = _T_15090 ? _T_10366_0 : _T_15089; // @[Mux.scala 46:16:@11380.4]
  assign _T_15142 = 6'h31 == _T_11317_48; // @[Mux.scala 46:19:@11382.4]
  assign _T_15143 = _T_15142 ? _T_10366_48 : 8'h0; // @[Mux.scala 46:16:@11383.4]
  assign _T_15144 = 6'h30 == _T_11317_48; // @[Mux.scala 46:19:@11384.4]
  assign _T_15145 = _T_15144 ? _T_10366_47 : _T_15143; // @[Mux.scala 46:16:@11385.4]
  assign _T_15146 = 6'h2f == _T_11317_48; // @[Mux.scala 46:19:@11386.4]
  assign _T_15147 = _T_15146 ? _T_10366_46 : _T_15145; // @[Mux.scala 46:16:@11387.4]
  assign _T_15148 = 6'h2e == _T_11317_48; // @[Mux.scala 46:19:@11388.4]
  assign _T_15149 = _T_15148 ? _T_10366_45 : _T_15147; // @[Mux.scala 46:16:@11389.4]
  assign _T_15150 = 6'h2d == _T_11317_48; // @[Mux.scala 46:19:@11390.4]
  assign _T_15151 = _T_15150 ? _T_10366_44 : _T_15149; // @[Mux.scala 46:16:@11391.4]
  assign _T_15152 = 6'h2c == _T_11317_48; // @[Mux.scala 46:19:@11392.4]
  assign _T_15153 = _T_15152 ? _T_10366_43 : _T_15151; // @[Mux.scala 46:16:@11393.4]
  assign _T_15154 = 6'h2b == _T_11317_48; // @[Mux.scala 46:19:@11394.4]
  assign _T_15155 = _T_15154 ? _T_10366_42 : _T_15153; // @[Mux.scala 46:16:@11395.4]
  assign _T_15156 = 6'h2a == _T_11317_48; // @[Mux.scala 46:19:@11396.4]
  assign _T_15157 = _T_15156 ? _T_10366_41 : _T_15155; // @[Mux.scala 46:16:@11397.4]
  assign _T_15158 = 6'h29 == _T_11317_48; // @[Mux.scala 46:19:@11398.4]
  assign _T_15159 = _T_15158 ? _T_10366_40 : _T_15157; // @[Mux.scala 46:16:@11399.4]
  assign _T_15160 = 6'h28 == _T_11317_48; // @[Mux.scala 46:19:@11400.4]
  assign _T_15161 = _T_15160 ? _T_10366_39 : _T_15159; // @[Mux.scala 46:16:@11401.4]
  assign _T_15162 = 6'h27 == _T_11317_48; // @[Mux.scala 46:19:@11402.4]
  assign _T_15163 = _T_15162 ? _T_10366_38 : _T_15161; // @[Mux.scala 46:16:@11403.4]
  assign _T_15164 = 6'h26 == _T_11317_48; // @[Mux.scala 46:19:@11404.4]
  assign _T_15165 = _T_15164 ? _T_10366_37 : _T_15163; // @[Mux.scala 46:16:@11405.4]
  assign _T_15166 = 6'h25 == _T_11317_48; // @[Mux.scala 46:19:@11406.4]
  assign _T_15167 = _T_15166 ? _T_10366_36 : _T_15165; // @[Mux.scala 46:16:@11407.4]
  assign _T_15168 = 6'h24 == _T_11317_48; // @[Mux.scala 46:19:@11408.4]
  assign _T_15169 = _T_15168 ? _T_10366_35 : _T_15167; // @[Mux.scala 46:16:@11409.4]
  assign _T_15170 = 6'h23 == _T_11317_48; // @[Mux.scala 46:19:@11410.4]
  assign _T_15171 = _T_15170 ? _T_10366_34 : _T_15169; // @[Mux.scala 46:16:@11411.4]
  assign _T_15172 = 6'h22 == _T_11317_48; // @[Mux.scala 46:19:@11412.4]
  assign _T_15173 = _T_15172 ? _T_10366_33 : _T_15171; // @[Mux.scala 46:16:@11413.4]
  assign _T_15174 = 6'h21 == _T_11317_48; // @[Mux.scala 46:19:@11414.4]
  assign _T_15175 = _T_15174 ? _T_10366_32 : _T_15173; // @[Mux.scala 46:16:@11415.4]
  assign _T_15176 = 6'h20 == _T_11317_48; // @[Mux.scala 46:19:@11416.4]
  assign _T_15177 = _T_15176 ? _T_10366_31 : _T_15175; // @[Mux.scala 46:16:@11417.4]
  assign _T_15178 = 6'h1f == _T_11317_48; // @[Mux.scala 46:19:@11418.4]
  assign _T_15179 = _T_15178 ? _T_10366_30 : _T_15177; // @[Mux.scala 46:16:@11419.4]
  assign _T_15180 = 6'h1e == _T_11317_48; // @[Mux.scala 46:19:@11420.4]
  assign _T_15181 = _T_15180 ? _T_10366_29 : _T_15179; // @[Mux.scala 46:16:@11421.4]
  assign _T_15182 = 6'h1d == _T_11317_48; // @[Mux.scala 46:19:@11422.4]
  assign _T_15183 = _T_15182 ? _T_10366_28 : _T_15181; // @[Mux.scala 46:16:@11423.4]
  assign _T_15184 = 6'h1c == _T_11317_48; // @[Mux.scala 46:19:@11424.4]
  assign _T_15185 = _T_15184 ? _T_10366_27 : _T_15183; // @[Mux.scala 46:16:@11425.4]
  assign _T_15186 = 6'h1b == _T_11317_48; // @[Mux.scala 46:19:@11426.4]
  assign _T_15187 = _T_15186 ? _T_10366_26 : _T_15185; // @[Mux.scala 46:16:@11427.4]
  assign _T_15188 = 6'h1a == _T_11317_48; // @[Mux.scala 46:19:@11428.4]
  assign _T_15189 = _T_15188 ? _T_10366_25 : _T_15187; // @[Mux.scala 46:16:@11429.4]
  assign _T_15190 = 6'h19 == _T_11317_48; // @[Mux.scala 46:19:@11430.4]
  assign _T_15191 = _T_15190 ? _T_10366_24 : _T_15189; // @[Mux.scala 46:16:@11431.4]
  assign _T_15192 = 6'h18 == _T_11317_48; // @[Mux.scala 46:19:@11432.4]
  assign _T_15193 = _T_15192 ? _T_10366_23 : _T_15191; // @[Mux.scala 46:16:@11433.4]
  assign _T_15194 = 6'h17 == _T_11317_48; // @[Mux.scala 46:19:@11434.4]
  assign _T_15195 = _T_15194 ? _T_10366_22 : _T_15193; // @[Mux.scala 46:16:@11435.4]
  assign _T_15196 = 6'h16 == _T_11317_48; // @[Mux.scala 46:19:@11436.4]
  assign _T_15197 = _T_15196 ? _T_10366_21 : _T_15195; // @[Mux.scala 46:16:@11437.4]
  assign _T_15198 = 6'h15 == _T_11317_48; // @[Mux.scala 46:19:@11438.4]
  assign _T_15199 = _T_15198 ? _T_10366_20 : _T_15197; // @[Mux.scala 46:16:@11439.4]
  assign _T_15200 = 6'h14 == _T_11317_48; // @[Mux.scala 46:19:@11440.4]
  assign _T_15201 = _T_15200 ? _T_10366_19 : _T_15199; // @[Mux.scala 46:16:@11441.4]
  assign _T_15202 = 6'h13 == _T_11317_48; // @[Mux.scala 46:19:@11442.4]
  assign _T_15203 = _T_15202 ? _T_10366_18 : _T_15201; // @[Mux.scala 46:16:@11443.4]
  assign _T_15204 = 6'h12 == _T_11317_48; // @[Mux.scala 46:19:@11444.4]
  assign _T_15205 = _T_15204 ? _T_10366_17 : _T_15203; // @[Mux.scala 46:16:@11445.4]
  assign _T_15206 = 6'h11 == _T_11317_48; // @[Mux.scala 46:19:@11446.4]
  assign _T_15207 = _T_15206 ? _T_10366_16 : _T_15205; // @[Mux.scala 46:16:@11447.4]
  assign _T_15208 = 6'h10 == _T_11317_48; // @[Mux.scala 46:19:@11448.4]
  assign _T_15209 = _T_15208 ? _T_10366_15 : _T_15207; // @[Mux.scala 46:16:@11449.4]
  assign _T_15210 = 6'hf == _T_11317_48; // @[Mux.scala 46:19:@11450.4]
  assign _T_15211 = _T_15210 ? _T_10366_14 : _T_15209; // @[Mux.scala 46:16:@11451.4]
  assign _T_15212 = 6'he == _T_11317_48; // @[Mux.scala 46:19:@11452.4]
  assign _T_15213 = _T_15212 ? _T_10366_13 : _T_15211; // @[Mux.scala 46:16:@11453.4]
  assign _T_15214 = 6'hd == _T_11317_48; // @[Mux.scala 46:19:@11454.4]
  assign _T_15215 = _T_15214 ? _T_10366_12 : _T_15213; // @[Mux.scala 46:16:@11455.4]
  assign _T_15216 = 6'hc == _T_11317_48; // @[Mux.scala 46:19:@11456.4]
  assign _T_15217 = _T_15216 ? _T_10366_11 : _T_15215; // @[Mux.scala 46:16:@11457.4]
  assign _T_15218 = 6'hb == _T_11317_48; // @[Mux.scala 46:19:@11458.4]
  assign _T_15219 = _T_15218 ? _T_10366_10 : _T_15217; // @[Mux.scala 46:16:@11459.4]
  assign _T_15220 = 6'ha == _T_11317_48; // @[Mux.scala 46:19:@11460.4]
  assign _T_15221 = _T_15220 ? _T_10366_9 : _T_15219; // @[Mux.scala 46:16:@11461.4]
  assign _T_15222 = 6'h9 == _T_11317_48; // @[Mux.scala 46:19:@11462.4]
  assign _T_15223 = _T_15222 ? _T_10366_8 : _T_15221; // @[Mux.scala 46:16:@11463.4]
  assign _T_15224 = 6'h8 == _T_11317_48; // @[Mux.scala 46:19:@11464.4]
  assign _T_15225 = _T_15224 ? _T_10366_7 : _T_15223; // @[Mux.scala 46:16:@11465.4]
  assign _T_15226 = 6'h7 == _T_11317_48; // @[Mux.scala 46:19:@11466.4]
  assign _T_15227 = _T_15226 ? _T_10366_6 : _T_15225; // @[Mux.scala 46:16:@11467.4]
  assign _T_15228 = 6'h6 == _T_11317_48; // @[Mux.scala 46:19:@11468.4]
  assign _T_15229 = _T_15228 ? _T_10366_5 : _T_15227; // @[Mux.scala 46:16:@11469.4]
  assign _T_15230 = 6'h5 == _T_11317_48; // @[Mux.scala 46:19:@11470.4]
  assign _T_15231 = _T_15230 ? _T_10366_4 : _T_15229; // @[Mux.scala 46:16:@11471.4]
  assign _T_15232 = 6'h4 == _T_11317_48; // @[Mux.scala 46:19:@11472.4]
  assign _T_15233 = _T_15232 ? _T_10366_3 : _T_15231; // @[Mux.scala 46:16:@11473.4]
  assign _T_15234 = 6'h3 == _T_11317_48; // @[Mux.scala 46:19:@11474.4]
  assign _T_15235 = _T_15234 ? _T_10366_2 : _T_15233; // @[Mux.scala 46:16:@11475.4]
  assign _T_15236 = 6'h2 == _T_11317_48; // @[Mux.scala 46:19:@11476.4]
  assign _T_15237 = _T_15236 ? _T_10366_1 : _T_15235; // @[Mux.scala 46:16:@11477.4]
  assign _T_15238 = 6'h1 == _T_11317_48; // @[Mux.scala 46:19:@11478.4]
  assign _T_15239 = _T_15238 ? _T_10366_0 : _T_15237; // @[Mux.scala 46:16:@11479.4]
  assign _T_15291 = 6'h32 == _T_11317_49; // @[Mux.scala 46:19:@11481.4]
  assign _T_15292 = _T_15291 ? _T_10366_49 : 8'h0; // @[Mux.scala 46:16:@11482.4]
  assign _T_15293 = 6'h31 == _T_11317_49; // @[Mux.scala 46:19:@11483.4]
  assign _T_15294 = _T_15293 ? _T_10366_48 : _T_15292; // @[Mux.scala 46:16:@11484.4]
  assign _T_15295 = 6'h30 == _T_11317_49; // @[Mux.scala 46:19:@11485.4]
  assign _T_15296 = _T_15295 ? _T_10366_47 : _T_15294; // @[Mux.scala 46:16:@11486.4]
  assign _T_15297 = 6'h2f == _T_11317_49; // @[Mux.scala 46:19:@11487.4]
  assign _T_15298 = _T_15297 ? _T_10366_46 : _T_15296; // @[Mux.scala 46:16:@11488.4]
  assign _T_15299 = 6'h2e == _T_11317_49; // @[Mux.scala 46:19:@11489.4]
  assign _T_15300 = _T_15299 ? _T_10366_45 : _T_15298; // @[Mux.scala 46:16:@11490.4]
  assign _T_15301 = 6'h2d == _T_11317_49; // @[Mux.scala 46:19:@11491.4]
  assign _T_15302 = _T_15301 ? _T_10366_44 : _T_15300; // @[Mux.scala 46:16:@11492.4]
  assign _T_15303 = 6'h2c == _T_11317_49; // @[Mux.scala 46:19:@11493.4]
  assign _T_15304 = _T_15303 ? _T_10366_43 : _T_15302; // @[Mux.scala 46:16:@11494.4]
  assign _T_15305 = 6'h2b == _T_11317_49; // @[Mux.scala 46:19:@11495.4]
  assign _T_15306 = _T_15305 ? _T_10366_42 : _T_15304; // @[Mux.scala 46:16:@11496.4]
  assign _T_15307 = 6'h2a == _T_11317_49; // @[Mux.scala 46:19:@11497.4]
  assign _T_15308 = _T_15307 ? _T_10366_41 : _T_15306; // @[Mux.scala 46:16:@11498.4]
  assign _T_15309 = 6'h29 == _T_11317_49; // @[Mux.scala 46:19:@11499.4]
  assign _T_15310 = _T_15309 ? _T_10366_40 : _T_15308; // @[Mux.scala 46:16:@11500.4]
  assign _T_15311 = 6'h28 == _T_11317_49; // @[Mux.scala 46:19:@11501.4]
  assign _T_15312 = _T_15311 ? _T_10366_39 : _T_15310; // @[Mux.scala 46:16:@11502.4]
  assign _T_15313 = 6'h27 == _T_11317_49; // @[Mux.scala 46:19:@11503.4]
  assign _T_15314 = _T_15313 ? _T_10366_38 : _T_15312; // @[Mux.scala 46:16:@11504.4]
  assign _T_15315 = 6'h26 == _T_11317_49; // @[Mux.scala 46:19:@11505.4]
  assign _T_15316 = _T_15315 ? _T_10366_37 : _T_15314; // @[Mux.scala 46:16:@11506.4]
  assign _T_15317 = 6'h25 == _T_11317_49; // @[Mux.scala 46:19:@11507.4]
  assign _T_15318 = _T_15317 ? _T_10366_36 : _T_15316; // @[Mux.scala 46:16:@11508.4]
  assign _T_15319 = 6'h24 == _T_11317_49; // @[Mux.scala 46:19:@11509.4]
  assign _T_15320 = _T_15319 ? _T_10366_35 : _T_15318; // @[Mux.scala 46:16:@11510.4]
  assign _T_15321 = 6'h23 == _T_11317_49; // @[Mux.scala 46:19:@11511.4]
  assign _T_15322 = _T_15321 ? _T_10366_34 : _T_15320; // @[Mux.scala 46:16:@11512.4]
  assign _T_15323 = 6'h22 == _T_11317_49; // @[Mux.scala 46:19:@11513.4]
  assign _T_15324 = _T_15323 ? _T_10366_33 : _T_15322; // @[Mux.scala 46:16:@11514.4]
  assign _T_15325 = 6'h21 == _T_11317_49; // @[Mux.scala 46:19:@11515.4]
  assign _T_15326 = _T_15325 ? _T_10366_32 : _T_15324; // @[Mux.scala 46:16:@11516.4]
  assign _T_15327 = 6'h20 == _T_11317_49; // @[Mux.scala 46:19:@11517.4]
  assign _T_15328 = _T_15327 ? _T_10366_31 : _T_15326; // @[Mux.scala 46:16:@11518.4]
  assign _T_15329 = 6'h1f == _T_11317_49; // @[Mux.scala 46:19:@11519.4]
  assign _T_15330 = _T_15329 ? _T_10366_30 : _T_15328; // @[Mux.scala 46:16:@11520.4]
  assign _T_15331 = 6'h1e == _T_11317_49; // @[Mux.scala 46:19:@11521.4]
  assign _T_15332 = _T_15331 ? _T_10366_29 : _T_15330; // @[Mux.scala 46:16:@11522.4]
  assign _T_15333 = 6'h1d == _T_11317_49; // @[Mux.scala 46:19:@11523.4]
  assign _T_15334 = _T_15333 ? _T_10366_28 : _T_15332; // @[Mux.scala 46:16:@11524.4]
  assign _T_15335 = 6'h1c == _T_11317_49; // @[Mux.scala 46:19:@11525.4]
  assign _T_15336 = _T_15335 ? _T_10366_27 : _T_15334; // @[Mux.scala 46:16:@11526.4]
  assign _T_15337 = 6'h1b == _T_11317_49; // @[Mux.scala 46:19:@11527.4]
  assign _T_15338 = _T_15337 ? _T_10366_26 : _T_15336; // @[Mux.scala 46:16:@11528.4]
  assign _T_15339 = 6'h1a == _T_11317_49; // @[Mux.scala 46:19:@11529.4]
  assign _T_15340 = _T_15339 ? _T_10366_25 : _T_15338; // @[Mux.scala 46:16:@11530.4]
  assign _T_15341 = 6'h19 == _T_11317_49; // @[Mux.scala 46:19:@11531.4]
  assign _T_15342 = _T_15341 ? _T_10366_24 : _T_15340; // @[Mux.scala 46:16:@11532.4]
  assign _T_15343 = 6'h18 == _T_11317_49; // @[Mux.scala 46:19:@11533.4]
  assign _T_15344 = _T_15343 ? _T_10366_23 : _T_15342; // @[Mux.scala 46:16:@11534.4]
  assign _T_15345 = 6'h17 == _T_11317_49; // @[Mux.scala 46:19:@11535.4]
  assign _T_15346 = _T_15345 ? _T_10366_22 : _T_15344; // @[Mux.scala 46:16:@11536.4]
  assign _T_15347 = 6'h16 == _T_11317_49; // @[Mux.scala 46:19:@11537.4]
  assign _T_15348 = _T_15347 ? _T_10366_21 : _T_15346; // @[Mux.scala 46:16:@11538.4]
  assign _T_15349 = 6'h15 == _T_11317_49; // @[Mux.scala 46:19:@11539.4]
  assign _T_15350 = _T_15349 ? _T_10366_20 : _T_15348; // @[Mux.scala 46:16:@11540.4]
  assign _T_15351 = 6'h14 == _T_11317_49; // @[Mux.scala 46:19:@11541.4]
  assign _T_15352 = _T_15351 ? _T_10366_19 : _T_15350; // @[Mux.scala 46:16:@11542.4]
  assign _T_15353 = 6'h13 == _T_11317_49; // @[Mux.scala 46:19:@11543.4]
  assign _T_15354 = _T_15353 ? _T_10366_18 : _T_15352; // @[Mux.scala 46:16:@11544.4]
  assign _T_15355 = 6'h12 == _T_11317_49; // @[Mux.scala 46:19:@11545.4]
  assign _T_15356 = _T_15355 ? _T_10366_17 : _T_15354; // @[Mux.scala 46:16:@11546.4]
  assign _T_15357 = 6'h11 == _T_11317_49; // @[Mux.scala 46:19:@11547.4]
  assign _T_15358 = _T_15357 ? _T_10366_16 : _T_15356; // @[Mux.scala 46:16:@11548.4]
  assign _T_15359 = 6'h10 == _T_11317_49; // @[Mux.scala 46:19:@11549.4]
  assign _T_15360 = _T_15359 ? _T_10366_15 : _T_15358; // @[Mux.scala 46:16:@11550.4]
  assign _T_15361 = 6'hf == _T_11317_49; // @[Mux.scala 46:19:@11551.4]
  assign _T_15362 = _T_15361 ? _T_10366_14 : _T_15360; // @[Mux.scala 46:16:@11552.4]
  assign _T_15363 = 6'he == _T_11317_49; // @[Mux.scala 46:19:@11553.4]
  assign _T_15364 = _T_15363 ? _T_10366_13 : _T_15362; // @[Mux.scala 46:16:@11554.4]
  assign _T_15365 = 6'hd == _T_11317_49; // @[Mux.scala 46:19:@11555.4]
  assign _T_15366 = _T_15365 ? _T_10366_12 : _T_15364; // @[Mux.scala 46:16:@11556.4]
  assign _T_15367 = 6'hc == _T_11317_49; // @[Mux.scala 46:19:@11557.4]
  assign _T_15368 = _T_15367 ? _T_10366_11 : _T_15366; // @[Mux.scala 46:16:@11558.4]
  assign _T_15369 = 6'hb == _T_11317_49; // @[Mux.scala 46:19:@11559.4]
  assign _T_15370 = _T_15369 ? _T_10366_10 : _T_15368; // @[Mux.scala 46:16:@11560.4]
  assign _T_15371 = 6'ha == _T_11317_49; // @[Mux.scala 46:19:@11561.4]
  assign _T_15372 = _T_15371 ? _T_10366_9 : _T_15370; // @[Mux.scala 46:16:@11562.4]
  assign _T_15373 = 6'h9 == _T_11317_49; // @[Mux.scala 46:19:@11563.4]
  assign _T_15374 = _T_15373 ? _T_10366_8 : _T_15372; // @[Mux.scala 46:16:@11564.4]
  assign _T_15375 = 6'h8 == _T_11317_49; // @[Mux.scala 46:19:@11565.4]
  assign _T_15376 = _T_15375 ? _T_10366_7 : _T_15374; // @[Mux.scala 46:16:@11566.4]
  assign _T_15377 = 6'h7 == _T_11317_49; // @[Mux.scala 46:19:@11567.4]
  assign _T_15378 = _T_15377 ? _T_10366_6 : _T_15376; // @[Mux.scala 46:16:@11568.4]
  assign _T_15379 = 6'h6 == _T_11317_49; // @[Mux.scala 46:19:@11569.4]
  assign _T_15380 = _T_15379 ? _T_10366_5 : _T_15378; // @[Mux.scala 46:16:@11570.4]
  assign _T_15381 = 6'h5 == _T_11317_49; // @[Mux.scala 46:19:@11571.4]
  assign _T_15382 = _T_15381 ? _T_10366_4 : _T_15380; // @[Mux.scala 46:16:@11572.4]
  assign _T_15383 = 6'h4 == _T_11317_49; // @[Mux.scala 46:19:@11573.4]
  assign _T_15384 = _T_15383 ? _T_10366_3 : _T_15382; // @[Mux.scala 46:16:@11574.4]
  assign _T_15385 = 6'h3 == _T_11317_49; // @[Mux.scala 46:19:@11575.4]
  assign _T_15386 = _T_15385 ? _T_10366_2 : _T_15384; // @[Mux.scala 46:16:@11576.4]
  assign _T_15387 = 6'h2 == _T_11317_49; // @[Mux.scala 46:19:@11577.4]
  assign _T_15388 = _T_15387 ? _T_10366_1 : _T_15386; // @[Mux.scala 46:16:@11578.4]
  assign _T_15389 = 6'h1 == _T_11317_49; // @[Mux.scala 46:19:@11579.4]
  assign _T_15390 = _T_15389 ? _T_10366_0 : _T_15388; // @[Mux.scala 46:16:@11580.4]
  assign _T_15443 = 6'h33 == _T_11317_50; // @[Mux.scala 46:19:@11582.4]
  assign _T_15444 = _T_15443 ? _T_10366_50 : 8'h0; // @[Mux.scala 46:16:@11583.4]
  assign _T_15445 = 6'h32 == _T_11317_50; // @[Mux.scala 46:19:@11584.4]
  assign _T_15446 = _T_15445 ? _T_10366_49 : _T_15444; // @[Mux.scala 46:16:@11585.4]
  assign _T_15447 = 6'h31 == _T_11317_50; // @[Mux.scala 46:19:@11586.4]
  assign _T_15448 = _T_15447 ? _T_10366_48 : _T_15446; // @[Mux.scala 46:16:@11587.4]
  assign _T_15449 = 6'h30 == _T_11317_50; // @[Mux.scala 46:19:@11588.4]
  assign _T_15450 = _T_15449 ? _T_10366_47 : _T_15448; // @[Mux.scala 46:16:@11589.4]
  assign _T_15451 = 6'h2f == _T_11317_50; // @[Mux.scala 46:19:@11590.4]
  assign _T_15452 = _T_15451 ? _T_10366_46 : _T_15450; // @[Mux.scala 46:16:@11591.4]
  assign _T_15453 = 6'h2e == _T_11317_50; // @[Mux.scala 46:19:@11592.4]
  assign _T_15454 = _T_15453 ? _T_10366_45 : _T_15452; // @[Mux.scala 46:16:@11593.4]
  assign _T_15455 = 6'h2d == _T_11317_50; // @[Mux.scala 46:19:@11594.4]
  assign _T_15456 = _T_15455 ? _T_10366_44 : _T_15454; // @[Mux.scala 46:16:@11595.4]
  assign _T_15457 = 6'h2c == _T_11317_50; // @[Mux.scala 46:19:@11596.4]
  assign _T_15458 = _T_15457 ? _T_10366_43 : _T_15456; // @[Mux.scala 46:16:@11597.4]
  assign _T_15459 = 6'h2b == _T_11317_50; // @[Mux.scala 46:19:@11598.4]
  assign _T_15460 = _T_15459 ? _T_10366_42 : _T_15458; // @[Mux.scala 46:16:@11599.4]
  assign _T_15461 = 6'h2a == _T_11317_50; // @[Mux.scala 46:19:@11600.4]
  assign _T_15462 = _T_15461 ? _T_10366_41 : _T_15460; // @[Mux.scala 46:16:@11601.4]
  assign _T_15463 = 6'h29 == _T_11317_50; // @[Mux.scala 46:19:@11602.4]
  assign _T_15464 = _T_15463 ? _T_10366_40 : _T_15462; // @[Mux.scala 46:16:@11603.4]
  assign _T_15465 = 6'h28 == _T_11317_50; // @[Mux.scala 46:19:@11604.4]
  assign _T_15466 = _T_15465 ? _T_10366_39 : _T_15464; // @[Mux.scala 46:16:@11605.4]
  assign _T_15467 = 6'h27 == _T_11317_50; // @[Mux.scala 46:19:@11606.4]
  assign _T_15468 = _T_15467 ? _T_10366_38 : _T_15466; // @[Mux.scala 46:16:@11607.4]
  assign _T_15469 = 6'h26 == _T_11317_50; // @[Mux.scala 46:19:@11608.4]
  assign _T_15470 = _T_15469 ? _T_10366_37 : _T_15468; // @[Mux.scala 46:16:@11609.4]
  assign _T_15471 = 6'h25 == _T_11317_50; // @[Mux.scala 46:19:@11610.4]
  assign _T_15472 = _T_15471 ? _T_10366_36 : _T_15470; // @[Mux.scala 46:16:@11611.4]
  assign _T_15473 = 6'h24 == _T_11317_50; // @[Mux.scala 46:19:@11612.4]
  assign _T_15474 = _T_15473 ? _T_10366_35 : _T_15472; // @[Mux.scala 46:16:@11613.4]
  assign _T_15475 = 6'h23 == _T_11317_50; // @[Mux.scala 46:19:@11614.4]
  assign _T_15476 = _T_15475 ? _T_10366_34 : _T_15474; // @[Mux.scala 46:16:@11615.4]
  assign _T_15477 = 6'h22 == _T_11317_50; // @[Mux.scala 46:19:@11616.4]
  assign _T_15478 = _T_15477 ? _T_10366_33 : _T_15476; // @[Mux.scala 46:16:@11617.4]
  assign _T_15479 = 6'h21 == _T_11317_50; // @[Mux.scala 46:19:@11618.4]
  assign _T_15480 = _T_15479 ? _T_10366_32 : _T_15478; // @[Mux.scala 46:16:@11619.4]
  assign _T_15481 = 6'h20 == _T_11317_50; // @[Mux.scala 46:19:@11620.4]
  assign _T_15482 = _T_15481 ? _T_10366_31 : _T_15480; // @[Mux.scala 46:16:@11621.4]
  assign _T_15483 = 6'h1f == _T_11317_50; // @[Mux.scala 46:19:@11622.4]
  assign _T_15484 = _T_15483 ? _T_10366_30 : _T_15482; // @[Mux.scala 46:16:@11623.4]
  assign _T_15485 = 6'h1e == _T_11317_50; // @[Mux.scala 46:19:@11624.4]
  assign _T_15486 = _T_15485 ? _T_10366_29 : _T_15484; // @[Mux.scala 46:16:@11625.4]
  assign _T_15487 = 6'h1d == _T_11317_50; // @[Mux.scala 46:19:@11626.4]
  assign _T_15488 = _T_15487 ? _T_10366_28 : _T_15486; // @[Mux.scala 46:16:@11627.4]
  assign _T_15489 = 6'h1c == _T_11317_50; // @[Mux.scala 46:19:@11628.4]
  assign _T_15490 = _T_15489 ? _T_10366_27 : _T_15488; // @[Mux.scala 46:16:@11629.4]
  assign _T_15491 = 6'h1b == _T_11317_50; // @[Mux.scala 46:19:@11630.4]
  assign _T_15492 = _T_15491 ? _T_10366_26 : _T_15490; // @[Mux.scala 46:16:@11631.4]
  assign _T_15493 = 6'h1a == _T_11317_50; // @[Mux.scala 46:19:@11632.4]
  assign _T_15494 = _T_15493 ? _T_10366_25 : _T_15492; // @[Mux.scala 46:16:@11633.4]
  assign _T_15495 = 6'h19 == _T_11317_50; // @[Mux.scala 46:19:@11634.4]
  assign _T_15496 = _T_15495 ? _T_10366_24 : _T_15494; // @[Mux.scala 46:16:@11635.4]
  assign _T_15497 = 6'h18 == _T_11317_50; // @[Mux.scala 46:19:@11636.4]
  assign _T_15498 = _T_15497 ? _T_10366_23 : _T_15496; // @[Mux.scala 46:16:@11637.4]
  assign _T_15499 = 6'h17 == _T_11317_50; // @[Mux.scala 46:19:@11638.4]
  assign _T_15500 = _T_15499 ? _T_10366_22 : _T_15498; // @[Mux.scala 46:16:@11639.4]
  assign _T_15501 = 6'h16 == _T_11317_50; // @[Mux.scala 46:19:@11640.4]
  assign _T_15502 = _T_15501 ? _T_10366_21 : _T_15500; // @[Mux.scala 46:16:@11641.4]
  assign _T_15503 = 6'h15 == _T_11317_50; // @[Mux.scala 46:19:@11642.4]
  assign _T_15504 = _T_15503 ? _T_10366_20 : _T_15502; // @[Mux.scala 46:16:@11643.4]
  assign _T_15505 = 6'h14 == _T_11317_50; // @[Mux.scala 46:19:@11644.4]
  assign _T_15506 = _T_15505 ? _T_10366_19 : _T_15504; // @[Mux.scala 46:16:@11645.4]
  assign _T_15507 = 6'h13 == _T_11317_50; // @[Mux.scala 46:19:@11646.4]
  assign _T_15508 = _T_15507 ? _T_10366_18 : _T_15506; // @[Mux.scala 46:16:@11647.4]
  assign _T_15509 = 6'h12 == _T_11317_50; // @[Mux.scala 46:19:@11648.4]
  assign _T_15510 = _T_15509 ? _T_10366_17 : _T_15508; // @[Mux.scala 46:16:@11649.4]
  assign _T_15511 = 6'h11 == _T_11317_50; // @[Mux.scala 46:19:@11650.4]
  assign _T_15512 = _T_15511 ? _T_10366_16 : _T_15510; // @[Mux.scala 46:16:@11651.4]
  assign _T_15513 = 6'h10 == _T_11317_50; // @[Mux.scala 46:19:@11652.4]
  assign _T_15514 = _T_15513 ? _T_10366_15 : _T_15512; // @[Mux.scala 46:16:@11653.4]
  assign _T_15515 = 6'hf == _T_11317_50; // @[Mux.scala 46:19:@11654.4]
  assign _T_15516 = _T_15515 ? _T_10366_14 : _T_15514; // @[Mux.scala 46:16:@11655.4]
  assign _T_15517 = 6'he == _T_11317_50; // @[Mux.scala 46:19:@11656.4]
  assign _T_15518 = _T_15517 ? _T_10366_13 : _T_15516; // @[Mux.scala 46:16:@11657.4]
  assign _T_15519 = 6'hd == _T_11317_50; // @[Mux.scala 46:19:@11658.4]
  assign _T_15520 = _T_15519 ? _T_10366_12 : _T_15518; // @[Mux.scala 46:16:@11659.4]
  assign _T_15521 = 6'hc == _T_11317_50; // @[Mux.scala 46:19:@11660.4]
  assign _T_15522 = _T_15521 ? _T_10366_11 : _T_15520; // @[Mux.scala 46:16:@11661.4]
  assign _T_15523 = 6'hb == _T_11317_50; // @[Mux.scala 46:19:@11662.4]
  assign _T_15524 = _T_15523 ? _T_10366_10 : _T_15522; // @[Mux.scala 46:16:@11663.4]
  assign _T_15525 = 6'ha == _T_11317_50; // @[Mux.scala 46:19:@11664.4]
  assign _T_15526 = _T_15525 ? _T_10366_9 : _T_15524; // @[Mux.scala 46:16:@11665.4]
  assign _T_15527 = 6'h9 == _T_11317_50; // @[Mux.scala 46:19:@11666.4]
  assign _T_15528 = _T_15527 ? _T_10366_8 : _T_15526; // @[Mux.scala 46:16:@11667.4]
  assign _T_15529 = 6'h8 == _T_11317_50; // @[Mux.scala 46:19:@11668.4]
  assign _T_15530 = _T_15529 ? _T_10366_7 : _T_15528; // @[Mux.scala 46:16:@11669.4]
  assign _T_15531 = 6'h7 == _T_11317_50; // @[Mux.scala 46:19:@11670.4]
  assign _T_15532 = _T_15531 ? _T_10366_6 : _T_15530; // @[Mux.scala 46:16:@11671.4]
  assign _T_15533 = 6'h6 == _T_11317_50; // @[Mux.scala 46:19:@11672.4]
  assign _T_15534 = _T_15533 ? _T_10366_5 : _T_15532; // @[Mux.scala 46:16:@11673.4]
  assign _T_15535 = 6'h5 == _T_11317_50; // @[Mux.scala 46:19:@11674.4]
  assign _T_15536 = _T_15535 ? _T_10366_4 : _T_15534; // @[Mux.scala 46:16:@11675.4]
  assign _T_15537 = 6'h4 == _T_11317_50; // @[Mux.scala 46:19:@11676.4]
  assign _T_15538 = _T_15537 ? _T_10366_3 : _T_15536; // @[Mux.scala 46:16:@11677.4]
  assign _T_15539 = 6'h3 == _T_11317_50; // @[Mux.scala 46:19:@11678.4]
  assign _T_15540 = _T_15539 ? _T_10366_2 : _T_15538; // @[Mux.scala 46:16:@11679.4]
  assign _T_15541 = 6'h2 == _T_11317_50; // @[Mux.scala 46:19:@11680.4]
  assign _T_15542 = _T_15541 ? _T_10366_1 : _T_15540; // @[Mux.scala 46:16:@11681.4]
  assign _T_15543 = 6'h1 == _T_11317_50; // @[Mux.scala 46:19:@11682.4]
  assign _T_15544 = _T_15543 ? _T_10366_0 : _T_15542; // @[Mux.scala 46:16:@11683.4]
  assign _T_15598 = 6'h34 == _T_11317_51; // @[Mux.scala 46:19:@11685.4]
  assign _T_15599 = _T_15598 ? _T_10366_51 : 8'h0; // @[Mux.scala 46:16:@11686.4]
  assign _T_15600 = 6'h33 == _T_11317_51; // @[Mux.scala 46:19:@11687.4]
  assign _T_15601 = _T_15600 ? _T_10366_50 : _T_15599; // @[Mux.scala 46:16:@11688.4]
  assign _T_15602 = 6'h32 == _T_11317_51; // @[Mux.scala 46:19:@11689.4]
  assign _T_15603 = _T_15602 ? _T_10366_49 : _T_15601; // @[Mux.scala 46:16:@11690.4]
  assign _T_15604 = 6'h31 == _T_11317_51; // @[Mux.scala 46:19:@11691.4]
  assign _T_15605 = _T_15604 ? _T_10366_48 : _T_15603; // @[Mux.scala 46:16:@11692.4]
  assign _T_15606 = 6'h30 == _T_11317_51; // @[Mux.scala 46:19:@11693.4]
  assign _T_15607 = _T_15606 ? _T_10366_47 : _T_15605; // @[Mux.scala 46:16:@11694.4]
  assign _T_15608 = 6'h2f == _T_11317_51; // @[Mux.scala 46:19:@11695.4]
  assign _T_15609 = _T_15608 ? _T_10366_46 : _T_15607; // @[Mux.scala 46:16:@11696.4]
  assign _T_15610 = 6'h2e == _T_11317_51; // @[Mux.scala 46:19:@11697.4]
  assign _T_15611 = _T_15610 ? _T_10366_45 : _T_15609; // @[Mux.scala 46:16:@11698.4]
  assign _T_15612 = 6'h2d == _T_11317_51; // @[Mux.scala 46:19:@11699.4]
  assign _T_15613 = _T_15612 ? _T_10366_44 : _T_15611; // @[Mux.scala 46:16:@11700.4]
  assign _T_15614 = 6'h2c == _T_11317_51; // @[Mux.scala 46:19:@11701.4]
  assign _T_15615 = _T_15614 ? _T_10366_43 : _T_15613; // @[Mux.scala 46:16:@11702.4]
  assign _T_15616 = 6'h2b == _T_11317_51; // @[Mux.scala 46:19:@11703.4]
  assign _T_15617 = _T_15616 ? _T_10366_42 : _T_15615; // @[Mux.scala 46:16:@11704.4]
  assign _T_15618 = 6'h2a == _T_11317_51; // @[Mux.scala 46:19:@11705.4]
  assign _T_15619 = _T_15618 ? _T_10366_41 : _T_15617; // @[Mux.scala 46:16:@11706.4]
  assign _T_15620 = 6'h29 == _T_11317_51; // @[Mux.scala 46:19:@11707.4]
  assign _T_15621 = _T_15620 ? _T_10366_40 : _T_15619; // @[Mux.scala 46:16:@11708.4]
  assign _T_15622 = 6'h28 == _T_11317_51; // @[Mux.scala 46:19:@11709.4]
  assign _T_15623 = _T_15622 ? _T_10366_39 : _T_15621; // @[Mux.scala 46:16:@11710.4]
  assign _T_15624 = 6'h27 == _T_11317_51; // @[Mux.scala 46:19:@11711.4]
  assign _T_15625 = _T_15624 ? _T_10366_38 : _T_15623; // @[Mux.scala 46:16:@11712.4]
  assign _T_15626 = 6'h26 == _T_11317_51; // @[Mux.scala 46:19:@11713.4]
  assign _T_15627 = _T_15626 ? _T_10366_37 : _T_15625; // @[Mux.scala 46:16:@11714.4]
  assign _T_15628 = 6'h25 == _T_11317_51; // @[Mux.scala 46:19:@11715.4]
  assign _T_15629 = _T_15628 ? _T_10366_36 : _T_15627; // @[Mux.scala 46:16:@11716.4]
  assign _T_15630 = 6'h24 == _T_11317_51; // @[Mux.scala 46:19:@11717.4]
  assign _T_15631 = _T_15630 ? _T_10366_35 : _T_15629; // @[Mux.scala 46:16:@11718.4]
  assign _T_15632 = 6'h23 == _T_11317_51; // @[Mux.scala 46:19:@11719.4]
  assign _T_15633 = _T_15632 ? _T_10366_34 : _T_15631; // @[Mux.scala 46:16:@11720.4]
  assign _T_15634 = 6'h22 == _T_11317_51; // @[Mux.scala 46:19:@11721.4]
  assign _T_15635 = _T_15634 ? _T_10366_33 : _T_15633; // @[Mux.scala 46:16:@11722.4]
  assign _T_15636 = 6'h21 == _T_11317_51; // @[Mux.scala 46:19:@11723.4]
  assign _T_15637 = _T_15636 ? _T_10366_32 : _T_15635; // @[Mux.scala 46:16:@11724.4]
  assign _T_15638 = 6'h20 == _T_11317_51; // @[Mux.scala 46:19:@11725.4]
  assign _T_15639 = _T_15638 ? _T_10366_31 : _T_15637; // @[Mux.scala 46:16:@11726.4]
  assign _T_15640 = 6'h1f == _T_11317_51; // @[Mux.scala 46:19:@11727.4]
  assign _T_15641 = _T_15640 ? _T_10366_30 : _T_15639; // @[Mux.scala 46:16:@11728.4]
  assign _T_15642 = 6'h1e == _T_11317_51; // @[Mux.scala 46:19:@11729.4]
  assign _T_15643 = _T_15642 ? _T_10366_29 : _T_15641; // @[Mux.scala 46:16:@11730.4]
  assign _T_15644 = 6'h1d == _T_11317_51; // @[Mux.scala 46:19:@11731.4]
  assign _T_15645 = _T_15644 ? _T_10366_28 : _T_15643; // @[Mux.scala 46:16:@11732.4]
  assign _T_15646 = 6'h1c == _T_11317_51; // @[Mux.scala 46:19:@11733.4]
  assign _T_15647 = _T_15646 ? _T_10366_27 : _T_15645; // @[Mux.scala 46:16:@11734.4]
  assign _T_15648 = 6'h1b == _T_11317_51; // @[Mux.scala 46:19:@11735.4]
  assign _T_15649 = _T_15648 ? _T_10366_26 : _T_15647; // @[Mux.scala 46:16:@11736.4]
  assign _T_15650 = 6'h1a == _T_11317_51; // @[Mux.scala 46:19:@11737.4]
  assign _T_15651 = _T_15650 ? _T_10366_25 : _T_15649; // @[Mux.scala 46:16:@11738.4]
  assign _T_15652 = 6'h19 == _T_11317_51; // @[Mux.scala 46:19:@11739.4]
  assign _T_15653 = _T_15652 ? _T_10366_24 : _T_15651; // @[Mux.scala 46:16:@11740.4]
  assign _T_15654 = 6'h18 == _T_11317_51; // @[Mux.scala 46:19:@11741.4]
  assign _T_15655 = _T_15654 ? _T_10366_23 : _T_15653; // @[Mux.scala 46:16:@11742.4]
  assign _T_15656 = 6'h17 == _T_11317_51; // @[Mux.scala 46:19:@11743.4]
  assign _T_15657 = _T_15656 ? _T_10366_22 : _T_15655; // @[Mux.scala 46:16:@11744.4]
  assign _T_15658 = 6'h16 == _T_11317_51; // @[Mux.scala 46:19:@11745.4]
  assign _T_15659 = _T_15658 ? _T_10366_21 : _T_15657; // @[Mux.scala 46:16:@11746.4]
  assign _T_15660 = 6'h15 == _T_11317_51; // @[Mux.scala 46:19:@11747.4]
  assign _T_15661 = _T_15660 ? _T_10366_20 : _T_15659; // @[Mux.scala 46:16:@11748.4]
  assign _T_15662 = 6'h14 == _T_11317_51; // @[Mux.scala 46:19:@11749.4]
  assign _T_15663 = _T_15662 ? _T_10366_19 : _T_15661; // @[Mux.scala 46:16:@11750.4]
  assign _T_15664 = 6'h13 == _T_11317_51; // @[Mux.scala 46:19:@11751.4]
  assign _T_15665 = _T_15664 ? _T_10366_18 : _T_15663; // @[Mux.scala 46:16:@11752.4]
  assign _T_15666 = 6'h12 == _T_11317_51; // @[Mux.scala 46:19:@11753.4]
  assign _T_15667 = _T_15666 ? _T_10366_17 : _T_15665; // @[Mux.scala 46:16:@11754.4]
  assign _T_15668 = 6'h11 == _T_11317_51; // @[Mux.scala 46:19:@11755.4]
  assign _T_15669 = _T_15668 ? _T_10366_16 : _T_15667; // @[Mux.scala 46:16:@11756.4]
  assign _T_15670 = 6'h10 == _T_11317_51; // @[Mux.scala 46:19:@11757.4]
  assign _T_15671 = _T_15670 ? _T_10366_15 : _T_15669; // @[Mux.scala 46:16:@11758.4]
  assign _T_15672 = 6'hf == _T_11317_51; // @[Mux.scala 46:19:@11759.4]
  assign _T_15673 = _T_15672 ? _T_10366_14 : _T_15671; // @[Mux.scala 46:16:@11760.4]
  assign _T_15674 = 6'he == _T_11317_51; // @[Mux.scala 46:19:@11761.4]
  assign _T_15675 = _T_15674 ? _T_10366_13 : _T_15673; // @[Mux.scala 46:16:@11762.4]
  assign _T_15676 = 6'hd == _T_11317_51; // @[Mux.scala 46:19:@11763.4]
  assign _T_15677 = _T_15676 ? _T_10366_12 : _T_15675; // @[Mux.scala 46:16:@11764.4]
  assign _T_15678 = 6'hc == _T_11317_51; // @[Mux.scala 46:19:@11765.4]
  assign _T_15679 = _T_15678 ? _T_10366_11 : _T_15677; // @[Mux.scala 46:16:@11766.4]
  assign _T_15680 = 6'hb == _T_11317_51; // @[Mux.scala 46:19:@11767.4]
  assign _T_15681 = _T_15680 ? _T_10366_10 : _T_15679; // @[Mux.scala 46:16:@11768.4]
  assign _T_15682 = 6'ha == _T_11317_51; // @[Mux.scala 46:19:@11769.4]
  assign _T_15683 = _T_15682 ? _T_10366_9 : _T_15681; // @[Mux.scala 46:16:@11770.4]
  assign _T_15684 = 6'h9 == _T_11317_51; // @[Mux.scala 46:19:@11771.4]
  assign _T_15685 = _T_15684 ? _T_10366_8 : _T_15683; // @[Mux.scala 46:16:@11772.4]
  assign _T_15686 = 6'h8 == _T_11317_51; // @[Mux.scala 46:19:@11773.4]
  assign _T_15687 = _T_15686 ? _T_10366_7 : _T_15685; // @[Mux.scala 46:16:@11774.4]
  assign _T_15688 = 6'h7 == _T_11317_51; // @[Mux.scala 46:19:@11775.4]
  assign _T_15689 = _T_15688 ? _T_10366_6 : _T_15687; // @[Mux.scala 46:16:@11776.4]
  assign _T_15690 = 6'h6 == _T_11317_51; // @[Mux.scala 46:19:@11777.4]
  assign _T_15691 = _T_15690 ? _T_10366_5 : _T_15689; // @[Mux.scala 46:16:@11778.4]
  assign _T_15692 = 6'h5 == _T_11317_51; // @[Mux.scala 46:19:@11779.4]
  assign _T_15693 = _T_15692 ? _T_10366_4 : _T_15691; // @[Mux.scala 46:16:@11780.4]
  assign _T_15694 = 6'h4 == _T_11317_51; // @[Mux.scala 46:19:@11781.4]
  assign _T_15695 = _T_15694 ? _T_10366_3 : _T_15693; // @[Mux.scala 46:16:@11782.4]
  assign _T_15696 = 6'h3 == _T_11317_51; // @[Mux.scala 46:19:@11783.4]
  assign _T_15697 = _T_15696 ? _T_10366_2 : _T_15695; // @[Mux.scala 46:16:@11784.4]
  assign _T_15698 = 6'h2 == _T_11317_51; // @[Mux.scala 46:19:@11785.4]
  assign _T_15699 = _T_15698 ? _T_10366_1 : _T_15697; // @[Mux.scala 46:16:@11786.4]
  assign _T_15700 = 6'h1 == _T_11317_51; // @[Mux.scala 46:19:@11787.4]
  assign _T_15701 = _T_15700 ? _T_10366_0 : _T_15699; // @[Mux.scala 46:16:@11788.4]
  assign _T_15756 = 6'h35 == _T_11317_52; // @[Mux.scala 46:19:@11790.4]
  assign _T_15757 = _T_15756 ? _T_10366_52 : 8'h0; // @[Mux.scala 46:16:@11791.4]
  assign _T_15758 = 6'h34 == _T_11317_52; // @[Mux.scala 46:19:@11792.4]
  assign _T_15759 = _T_15758 ? _T_10366_51 : _T_15757; // @[Mux.scala 46:16:@11793.4]
  assign _T_15760 = 6'h33 == _T_11317_52; // @[Mux.scala 46:19:@11794.4]
  assign _T_15761 = _T_15760 ? _T_10366_50 : _T_15759; // @[Mux.scala 46:16:@11795.4]
  assign _T_15762 = 6'h32 == _T_11317_52; // @[Mux.scala 46:19:@11796.4]
  assign _T_15763 = _T_15762 ? _T_10366_49 : _T_15761; // @[Mux.scala 46:16:@11797.4]
  assign _T_15764 = 6'h31 == _T_11317_52; // @[Mux.scala 46:19:@11798.4]
  assign _T_15765 = _T_15764 ? _T_10366_48 : _T_15763; // @[Mux.scala 46:16:@11799.4]
  assign _T_15766 = 6'h30 == _T_11317_52; // @[Mux.scala 46:19:@11800.4]
  assign _T_15767 = _T_15766 ? _T_10366_47 : _T_15765; // @[Mux.scala 46:16:@11801.4]
  assign _T_15768 = 6'h2f == _T_11317_52; // @[Mux.scala 46:19:@11802.4]
  assign _T_15769 = _T_15768 ? _T_10366_46 : _T_15767; // @[Mux.scala 46:16:@11803.4]
  assign _T_15770 = 6'h2e == _T_11317_52; // @[Mux.scala 46:19:@11804.4]
  assign _T_15771 = _T_15770 ? _T_10366_45 : _T_15769; // @[Mux.scala 46:16:@11805.4]
  assign _T_15772 = 6'h2d == _T_11317_52; // @[Mux.scala 46:19:@11806.4]
  assign _T_15773 = _T_15772 ? _T_10366_44 : _T_15771; // @[Mux.scala 46:16:@11807.4]
  assign _T_15774 = 6'h2c == _T_11317_52; // @[Mux.scala 46:19:@11808.4]
  assign _T_15775 = _T_15774 ? _T_10366_43 : _T_15773; // @[Mux.scala 46:16:@11809.4]
  assign _T_15776 = 6'h2b == _T_11317_52; // @[Mux.scala 46:19:@11810.4]
  assign _T_15777 = _T_15776 ? _T_10366_42 : _T_15775; // @[Mux.scala 46:16:@11811.4]
  assign _T_15778 = 6'h2a == _T_11317_52; // @[Mux.scala 46:19:@11812.4]
  assign _T_15779 = _T_15778 ? _T_10366_41 : _T_15777; // @[Mux.scala 46:16:@11813.4]
  assign _T_15780 = 6'h29 == _T_11317_52; // @[Mux.scala 46:19:@11814.4]
  assign _T_15781 = _T_15780 ? _T_10366_40 : _T_15779; // @[Mux.scala 46:16:@11815.4]
  assign _T_15782 = 6'h28 == _T_11317_52; // @[Mux.scala 46:19:@11816.4]
  assign _T_15783 = _T_15782 ? _T_10366_39 : _T_15781; // @[Mux.scala 46:16:@11817.4]
  assign _T_15784 = 6'h27 == _T_11317_52; // @[Mux.scala 46:19:@11818.4]
  assign _T_15785 = _T_15784 ? _T_10366_38 : _T_15783; // @[Mux.scala 46:16:@11819.4]
  assign _T_15786 = 6'h26 == _T_11317_52; // @[Mux.scala 46:19:@11820.4]
  assign _T_15787 = _T_15786 ? _T_10366_37 : _T_15785; // @[Mux.scala 46:16:@11821.4]
  assign _T_15788 = 6'h25 == _T_11317_52; // @[Mux.scala 46:19:@11822.4]
  assign _T_15789 = _T_15788 ? _T_10366_36 : _T_15787; // @[Mux.scala 46:16:@11823.4]
  assign _T_15790 = 6'h24 == _T_11317_52; // @[Mux.scala 46:19:@11824.4]
  assign _T_15791 = _T_15790 ? _T_10366_35 : _T_15789; // @[Mux.scala 46:16:@11825.4]
  assign _T_15792 = 6'h23 == _T_11317_52; // @[Mux.scala 46:19:@11826.4]
  assign _T_15793 = _T_15792 ? _T_10366_34 : _T_15791; // @[Mux.scala 46:16:@11827.4]
  assign _T_15794 = 6'h22 == _T_11317_52; // @[Mux.scala 46:19:@11828.4]
  assign _T_15795 = _T_15794 ? _T_10366_33 : _T_15793; // @[Mux.scala 46:16:@11829.4]
  assign _T_15796 = 6'h21 == _T_11317_52; // @[Mux.scala 46:19:@11830.4]
  assign _T_15797 = _T_15796 ? _T_10366_32 : _T_15795; // @[Mux.scala 46:16:@11831.4]
  assign _T_15798 = 6'h20 == _T_11317_52; // @[Mux.scala 46:19:@11832.4]
  assign _T_15799 = _T_15798 ? _T_10366_31 : _T_15797; // @[Mux.scala 46:16:@11833.4]
  assign _T_15800 = 6'h1f == _T_11317_52; // @[Mux.scala 46:19:@11834.4]
  assign _T_15801 = _T_15800 ? _T_10366_30 : _T_15799; // @[Mux.scala 46:16:@11835.4]
  assign _T_15802 = 6'h1e == _T_11317_52; // @[Mux.scala 46:19:@11836.4]
  assign _T_15803 = _T_15802 ? _T_10366_29 : _T_15801; // @[Mux.scala 46:16:@11837.4]
  assign _T_15804 = 6'h1d == _T_11317_52; // @[Mux.scala 46:19:@11838.4]
  assign _T_15805 = _T_15804 ? _T_10366_28 : _T_15803; // @[Mux.scala 46:16:@11839.4]
  assign _T_15806 = 6'h1c == _T_11317_52; // @[Mux.scala 46:19:@11840.4]
  assign _T_15807 = _T_15806 ? _T_10366_27 : _T_15805; // @[Mux.scala 46:16:@11841.4]
  assign _T_15808 = 6'h1b == _T_11317_52; // @[Mux.scala 46:19:@11842.4]
  assign _T_15809 = _T_15808 ? _T_10366_26 : _T_15807; // @[Mux.scala 46:16:@11843.4]
  assign _T_15810 = 6'h1a == _T_11317_52; // @[Mux.scala 46:19:@11844.4]
  assign _T_15811 = _T_15810 ? _T_10366_25 : _T_15809; // @[Mux.scala 46:16:@11845.4]
  assign _T_15812 = 6'h19 == _T_11317_52; // @[Mux.scala 46:19:@11846.4]
  assign _T_15813 = _T_15812 ? _T_10366_24 : _T_15811; // @[Mux.scala 46:16:@11847.4]
  assign _T_15814 = 6'h18 == _T_11317_52; // @[Mux.scala 46:19:@11848.4]
  assign _T_15815 = _T_15814 ? _T_10366_23 : _T_15813; // @[Mux.scala 46:16:@11849.4]
  assign _T_15816 = 6'h17 == _T_11317_52; // @[Mux.scala 46:19:@11850.4]
  assign _T_15817 = _T_15816 ? _T_10366_22 : _T_15815; // @[Mux.scala 46:16:@11851.4]
  assign _T_15818 = 6'h16 == _T_11317_52; // @[Mux.scala 46:19:@11852.4]
  assign _T_15819 = _T_15818 ? _T_10366_21 : _T_15817; // @[Mux.scala 46:16:@11853.4]
  assign _T_15820 = 6'h15 == _T_11317_52; // @[Mux.scala 46:19:@11854.4]
  assign _T_15821 = _T_15820 ? _T_10366_20 : _T_15819; // @[Mux.scala 46:16:@11855.4]
  assign _T_15822 = 6'h14 == _T_11317_52; // @[Mux.scala 46:19:@11856.4]
  assign _T_15823 = _T_15822 ? _T_10366_19 : _T_15821; // @[Mux.scala 46:16:@11857.4]
  assign _T_15824 = 6'h13 == _T_11317_52; // @[Mux.scala 46:19:@11858.4]
  assign _T_15825 = _T_15824 ? _T_10366_18 : _T_15823; // @[Mux.scala 46:16:@11859.4]
  assign _T_15826 = 6'h12 == _T_11317_52; // @[Mux.scala 46:19:@11860.4]
  assign _T_15827 = _T_15826 ? _T_10366_17 : _T_15825; // @[Mux.scala 46:16:@11861.4]
  assign _T_15828 = 6'h11 == _T_11317_52; // @[Mux.scala 46:19:@11862.4]
  assign _T_15829 = _T_15828 ? _T_10366_16 : _T_15827; // @[Mux.scala 46:16:@11863.4]
  assign _T_15830 = 6'h10 == _T_11317_52; // @[Mux.scala 46:19:@11864.4]
  assign _T_15831 = _T_15830 ? _T_10366_15 : _T_15829; // @[Mux.scala 46:16:@11865.4]
  assign _T_15832 = 6'hf == _T_11317_52; // @[Mux.scala 46:19:@11866.4]
  assign _T_15833 = _T_15832 ? _T_10366_14 : _T_15831; // @[Mux.scala 46:16:@11867.4]
  assign _T_15834 = 6'he == _T_11317_52; // @[Mux.scala 46:19:@11868.4]
  assign _T_15835 = _T_15834 ? _T_10366_13 : _T_15833; // @[Mux.scala 46:16:@11869.4]
  assign _T_15836 = 6'hd == _T_11317_52; // @[Mux.scala 46:19:@11870.4]
  assign _T_15837 = _T_15836 ? _T_10366_12 : _T_15835; // @[Mux.scala 46:16:@11871.4]
  assign _T_15838 = 6'hc == _T_11317_52; // @[Mux.scala 46:19:@11872.4]
  assign _T_15839 = _T_15838 ? _T_10366_11 : _T_15837; // @[Mux.scala 46:16:@11873.4]
  assign _T_15840 = 6'hb == _T_11317_52; // @[Mux.scala 46:19:@11874.4]
  assign _T_15841 = _T_15840 ? _T_10366_10 : _T_15839; // @[Mux.scala 46:16:@11875.4]
  assign _T_15842 = 6'ha == _T_11317_52; // @[Mux.scala 46:19:@11876.4]
  assign _T_15843 = _T_15842 ? _T_10366_9 : _T_15841; // @[Mux.scala 46:16:@11877.4]
  assign _T_15844 = 6'h9 == _T_11317_52; // @[Mux.scala 46:19:@11878.4]
  assign _T_15845 = _T_15844 ? _T_10366_8 : _T_15843; // @[Mux.scala 46:16:@11879.4]
  assign _T_15846 = 6'h8 == _T_11317_52; // @[Mux.scala 46:19:@11880.4]
  assign _T_15847 = _T_15846 ? _T_10366_7 : _T_15845; // @[Mux.scala 46:16:@11881.4]
  assign _T_15848 = 6'h7 == _T_11317_52; // @[Mux.scala 46:19:@11882.4]
  assign _T_15849 = _T_15848 ? _T_10366_6 : _T_15847; // @[Mux.scala 46:16:@11883.4]
  assign _T_15850 = 6'h6 == _T_11317_52; // @[Mux.scala 46:19:@11884.4]
  assign _T_15851 = _T_15850 ? _T_10366_5 : _T_15849; // @[Mux.scala 46:16:@11885.4]
  assign _T_15852 = 6'h5 == _T_11317_52; // @[Mux.scala 46:19:@11886.4]
  assign _T_15853 = _T_15852 ? _T_10366_4 : _T_15851; // @[Mux.scala 46:16:@11887.4]
  assign _T_15854 = 6'h4 == _T_11317_52; // @[Mux.scala 46:19:@11888.4]
  assign _T_15855 = _T_15854 ? _T_10366_3 : _T_15853; // @[Mux.scala 46:16:@11889.4]
  assign _T_15856 = 6'h3 == _T_11317_52; // @[Mux.scala 46:19:@11890.4]
  assign _T_15857 = _T_15856 ? _T_10366_2 : _T_15855; // @[Mux.scala 46:16:@11891.4]
  assign _T_15858 = 6'h2 == _T_11317_52; // @[Mux.scala 46:19:@11892.4]
  assign _T_15859 = _T_15858 ? _T_10366_1 : _T_15857; // @[Mux.scala 46:16:@11893.4]
  assign _T_15860 = 6'h1 == _T_11317_52; // @[Mux.scala 46:19:@11894.4]
  assign _T_15861 = _T_15860 ? _T_10366_0 : _T_15859; // @[Mux.scala 46:16:@11895.4]
  assign _T_15917 = 6'h36 == _T_11317_53; // @[Mux.scala 46:19:@11897.4]
  assign _T_15918 = _T_15917 ? _T_10366_53 : 8'h0; // @[Mux.scala 46:16:@11898.4]
  assign _T_15919 = 6'h35 == _T_11317_53; // @[Mux.scala 46:19:@11899.4]
  assign _T_15920 = _T_15919 ? _T_10366_52 : _T_15918; // @[Mux.scala 46:16:@11900.4]
  assign _T_15921 = 6'h34 == _T_11317_53; // @[Mux.scala 46:19:@11901.4]
  assign _T_15922 = _T_15921 ? _T_10366_51 : _T_15920; // @[Mux.scala 46:16:@11902.4]
  assign _T_15923 = 6'h33 == _T_11317_53; // @[Mux.scala 46:19:@11903.4]
  assign _T_15924 = _T_15923 ? _T_10366_50 : _T_15922; // @[Mux.scala 46:16:@11904.4]
  assign _T_15925 = 6'h32 == _T_11317_53; // @[Mux.scala 46:19:@11905.4]
  assign _T_15926 = _T_15925 ? _T_10366_49 : _T_15924; // @[Mux.scala 46:16:@11906.4]
  assign _T_15927 = 6'h31 == _T_11317_53; // @[Mux.scala 46:19:@11907.4]
  assign _T_15928 = _T_15927 ? _T_10366_48 : _T_15926; // @[Mux.scala 46:16:@11908.4]
  assign _T_15929 = 6'h30 == _T_11317_53; // @[Mux.scala 46:19:@11909.4]
  assign _T_15930 = _T_15929 ? _T_10366_47 : _T_15928; // @[Mux.scala 46:16:@11910.4]
  assign _T_15931 = 6'h2f == _T_11317_53; // @[Mux.scala 46:19:@11911.4]
  assign _T_15932 = _T_15931 ? _T_10366_46 : _T_15930; // @[Mux.scala 46:16:@11912.4]
  assign _T_15933 = 6'h2e == _T_11317_53; // @[Mux.scala 46:19:@11913.4]
  assign _T_15934 = _T_15933 ? _T_10366_45 : _T_15932; // @[Mux.scala 46:16:@11914.4]
  assign _T_15935 = 6'h2d == _T_11317_53; // @[Mux.scala 46:19:@11915.4]
  assign _T_15936 = _T_15935 ? _T_10366_44 : _T_15934; // @[Mux.scala 46:16:@11916.4]
  assign _T_15937 = 6'h2c == _T_11317_53; // @[Mux.scala 46:19:@11917.4]
  assign _T_15938 = _T_15937 ? _T_10366_43 : _T_15936; // @[Mux.scala 46:16:@11918.4]
  assign _T_15939 = 6'h2b == _T_11317_53; // @[Mux.scala 46:19:@11919.4]
  assign _T_15940 = _T_15939 ? _T_10366_42 : _T_15938; // @[Mux.scala 46:16:@11920.4]
  assign _T_15941 = 6'h2a == _T_11317_53; // @[Mux.scala 46:19:@11921.4]
  assign _T_15942 = _T_15941 ? _T_10366_41 : _T_15940; // @[Mux.scala 46:16:@11922.4]
  assign _T_15943 = 6'h29 == _T_11317_53; // @[Mux.scala 46:19:@11923.4]
  assign _T_15944 = _T_15943 ? _T_10366_40 : _T_15942; // @[Mux.scala 46:16:@11924.4]
  assign _T_15945 = 6'h28 == _T_11317_53; // @[Mux.scala 46:19:@11925.4]
  assign _T_15946 = _T_15945 ? _T_10366_39 : _T_15944; // @[Mux.scala 46:16:@11926.4]
  assign _T_15947 = 6'h27 == _T_11317_53; // @[Mux.scala 46:19:@11927.4]
  assign _T_15948 = _T_15947 ? _T_10366_38 : _T_15946; // @[Mux.scala 46:16:@11928.4]
  assign _T_15949 = 6'h26 == _T_11317_53; // @[Mux.scala 46:19:@11929.4]
  assign _T_15950 = _T_15949 ? _T_10366_37 : _T_15948; // @[Mux.scala 46:16:@11930.4]
  assign _T_15951 = 6'h25 == _T_11317_53; // @[Mux.scala 46:19:@11931.4]
  assign _T_15952 = _T_15951 ? _T_10366_36 : _T_15950; // @[Mux.scala 46:16:@11932.4]
  assign _T_15953 = 6'h24 == _T_11317_53; // @[Mux.scala 46:19:@11933.4]
  assign _T_15954 = _T_15953 ? _T_10366_35 : _T_15952; // @[Mux.scala 46:16:@11934.4]
  assign _T_15955 = 6'h23 == _T_11317_53; // @[Mux.scala 46:19:@11935.4]
  assign _T_15956 = _T_15955 ? _T_10366_34 : _T_15954; // @[Mux.scala 46:16:@11936.4]
  assign _T_15957 = 6'h22 == _T_11317_53; // @[Mux.scala 46:19:@11937.4]
  assign _T_15958 = _T_15957 ? _T_10366_33 : _T_15956; // @[Mux.scala 46:16:@11938.4]
  assign _T_15959 = 6'h21 == _T_11317_53; // @[Mux.scala 46:19:@11939.4]
  assign _T_15960 = _T_15959 ? _T_10366_32 : _T_15958; // @[Mux.scala 46:16:@11940.4]
  assign _T_15961 = 6'h20 == _T_11317_53; // @[Mux.scala 46:19:@11941.4]
  assign _T_15962 = _T_15961 ? _T_10366_31 : _T_15960; // @[Mux.scala 46:16:@11942.4]
  assign _T_15963 = 6'h1f == _T_11317_53; // @[Mux.scala 46:19:@11943.4]
  assign _T_15964 = _T_15963 ? _T_10366_30 : _T_15962; // @[Mux.scala 46:16:@11944.4]
  assign _T_15965 = 6'h1e == _T_11317_53; // @[Mux.scala 46:19:@11945.4]
  assign _T_15966 = _T_15965 ? _T_10366_29 : _T_15964; // @[Mux.scala 46:16:@11946.4]
  assign _T_15967 = 6'h1d == _T_11317_53; // @[Mux.scala 46:19:@11947.4]
  assign _T_15968 = _T_15967 ? _T_10366_28 : _T_15966; // @[Mux.scala 46:16:@11948.4]
  assign _T_15969 = 6'h1c == _T_11317_53; // @[Mux.scala 46:19:@11949.4]
  assign _T_15970 = _T_15969 ? _T_10366_27 : _T_15968; // @[Mux.scala 46:16:@11950.4]
  assign _T_15971 = 6'h1b == _T_11317_53; // @[Mux.scala 46:19:@11951.4]
  assign _T_15972 = _T_15971 ? _T_10366_26 : _T_15970; // @[Mux.scala 46:16:@11952.4]
  assign _T_15973 = 6'h1a == _T_11317_53; // @[Mux.scala 46:19:@11953.4]
  assign _T_15974 = _T_15973 ? _T_10366_25 : _T_15972; // @[Mux.scala 46:16:@11954.4]
  assign _T_15975 = 6'h19 == _T_11317_53; // @[Mux.scala 46:19:@11955.4]
  assign _T_15976 = _T_15975 ? _T_10366_24 : _T_15974; // @[Mux.scala 46:16:@11956.4]
  assign _T_15977 = 6'h18 == _T_11317_53; // @[Mux.scala 46:19:@11957.4]
  assign _T_15978 = _T_15977 ? _T_10366_23 : _T_15976; // @[Mux.scala 46:16:@11958.4]
  assign _T_15979 = 6'h17 == _T_11317_53; // @[Mux.scala 46:19:@11959.4]
  assign _T_15980 = _T_15979 ? _T_10366_22 : _T_15978; // @[Mux.scala 46:16:@11960.4]
  assign _T_15981 = 6'h16 == _T_11317_53; // @[Mux.scala 46:19:@11961.4]
  assign _T_15982 = _T_15981 ? _T_10366_21 : _T_15980; // @[Mux.scala 46:16:@11962.4]
  assign _T_15983 = 6'h15 == _T_11317_53; // @[Mux.scala 46:19:@11963.4]
  assign _T_15984 = _T_15983 ? _T_10366_20 : _T_15982; // @[Mux.scala 46:16:@11964.4]
  assign _T_15985 = 6'h14 == _T_11317_53; // @[Mux.scala 46:19:@11965.4]
  assign _T_15986 = _T_15985 ? _T_10366_19 : _T_15984; // @[Mux.scala 46:16:@11966.4]
  assign _T_15987 = 6'h13 == _T_11317_53; // @[Mux.scala 46:19:@11967.4]
  assign _T_15988 = _T_15987 ? _T_10366_18 : _T_15986; // @[Mux.scala 46:16:@11968.4]
  assign _T_15989 = 6'h12 == _T_11317_53; // @[Mux.scala 46:19:@11969.4]
  assign _T_15990 = _T_15989 ? _T_10366_17 : _T_15988; // @[Mux.scala 46:16:@11970.4]
  assign _T_15991 = 6'h11 == _T_11317_53; // @[Mux.scala 46:19:@11971.4]
  assign _T_15992 = _T_15991 ? _T_10366_16 : _T_15990; // @[Mux.scala 46:16:@11972.4]
  assign _T_15993 = 6'h10 == _T_11317_53; // @[Mux.scala 46:19:@11973.4]
  assign _T_15994 = _T_15993 ? _T_10366_15 : _T_15992; // @[Mux.scala 46:16:@11974.4]
  assign _T_15995 = 6'hf == _T_11317_53; // @[Mux.scala 46:19:@11975.4]
  assign _T_15996 = _T_15995 ? _T_10366_14 : _T_15994; // @[Mux.scala 46:16:@11976.4]
  assign _T_15997 = 6'he == _T_11317_53; // @[Mux.scala 46:19:@11977.4]
  assign _T_15998 = _T_15997 ? _T_10366_13 : _T_15996; // @[Mux.scala 46:16:@11978.4]
  assign _T_15999 = 6'hd == _T_11317_53; // @[Mux.scala 46:19:@11979.4]
  assign _T_16000 = _T_15999 ? _T_10366_12 : _T_15998; // @[Mux.scala 46:16:@11980.4]
  assign _T_16001 = 6'hc == _T_11317_53; // @[Mux.scala 46:19:@11981.4]
  assign _T_16002 = _T_16001 ? _T_10366_11 : _T_16000; // @[Mux.scala 46:16:@11982.4]
  assign _T_16003 = 6'hb == _T_11317_53; // @[Mux.scala 46:19:@11983.4]
  assign _T_16004 = _T_16003 ? _T_10366_10 : _T_16002; // @[Mux.scala 46:16:@11984.4]
  assign _T_16005 = 6'ha == _T_11317_53; // @[Mux.scala 46:19:@11985.4]
  assign _T_16006 = _T_16005 ? _T_10366_9 : _T_16004; // @[Mux.scala 46:16:@11986.4]
  assign _T_16007 = 6'h9 == _T_11317_53; // @[Mux.scala 46:19:@11987.4]
  assign _T_16008 = _T_16007 ? _T_10366_8 : _T_16006; // @[Mux.scala 46:16:@11988.4]
  assign _T_16009 = 6'h8 == _T_11317_53; // @[Mux.scala 46:19:@11989.4]
  assign _T_16010 = _T_16009 ? _T_10366_7 : _T_16008; // @[Mux.scala 46:16:@11990.4]
  assign _T_16011 = 6'h7 == _T_11317_53; // @[Mux.scala 46:19:@11991.4]
  assign _T_16012 = _T_16011 ? _T_10366_6 : _T_16010; // @[Mux.scala 46:16:@11992.4]
  assign _T_16013 = 6'h6 == _T_11317_53; // @[Mux.scala 46:19:@11993.4]
  assign _T_16014 = _T_16013 ? _T_10366_5 : _T_16012; // @[Mux.scala 46:16:@11994.4]
  assign _T_16015 = 6'h5 == _T_11317_53; // @[Mux.scala 46:19:@11995.4]
  assign _T_16016 = _T_16015 ? _T_10366_4 : _T_16014; // @[Mux.scala 46:16:@11996.4]
  assign _T_16017 = 6'h4 == _T_11317_53; // @[Mux.scala 46:19:@11997.4]
  assign _T_16018 = _T_16017 ? _T_10366_3 : _T_16016; // @[Mux.scala 46:16:@11998.4]
  assign _T_16019 = 6'h3 == _T_11317_53; // @[Mux.scala 46:19:@11999.4]
  assign _T_16020 = _T_16019 ? _T_10366_2 : _T_16018; // @[Mux.scala 46:16:@12000.4]
  assign _T_16021 = 6'h2 == _T_11317_53; // @[Mux.scala 46:19:@12001.4]
  assign _T_16022 = _T_16021 ? _T_10366_1 : _T_16020; // @[Mux.scala 46:16:@12002.4]
  assign _T_16023 = 6'h1 == _T_11317_53; // @[Mux.scala 46:19:@12003.4]
  assign _T_16024 = _T_16023 ? _T_10366_0 : _T_16022; // @[Mux.scala 46:16:@12004.4]
  assign _T_16081 = 6'h37 == _T_11317_54; // @[Mux.scala 46:19:@12006.4]
  assign _T_16082 = _T_16081 ? _T_10366_54 : 8'h0; // @[Mux.scala 46:16:@12007.4]
  assign _T_16083 = 6'h36 == _T_11317_54; // @[Mux.scala 46:19:@12008.4]
  assign _T_16084 = _T_16083 ? _T_10366_53 : _T_16082; // @[Mux.scala 46:16:@12009.4]
  assign _T_16085 = 6'h35 == _T_11317_54; // @[Mux.scala 46:19:@12010.4]
  assign _T_16086 = _T_16085 ? _T_10366_52 : _T_16084; // @[Mux.scala 46:16:@12011.4]
  assign _T_16087 = 6'h34 == _T_11317_54; // @[Mux.scala 46:19:@12012.4]
  assign _T_16088 = _T_16087 ? _T_10366_51 : _T_16086; // @[Mux.scala 46:16:@12013.4]
  assign _T_16089 = 6'h33 == _T_11317_54; // @[Mux.scala 46:19:@12014.4]
  assign _T_16090 = _T_16089 ? _T_10366_50 : _T_16088; // @[Mux.scala 46:16:@12015.4]
  assign _T_16091 = 6'h32 == _T_11317_54; // @[Mux.scala 46:19:@12016.4]
  assign _T_16092 = _T_16091 ? _T_10366_49 : _T_16090; // @[Mux.scala 46:16:@12017.4]
  assign _T_16093 = 6'h31 == _T_11317_54; // @[Mux.scala 46:19:@12018.4]
  assign _T_16094 = _T_16093 ? _T_10366_48 : _T_16092; // @[Mux.scala 46:16:@12019.4]
  assign _T_16095 = 6'h30 == _T_11317_54; // @[Mux.scala 46:19:@12020.4]
  assign _T_16096 = _T_16095 ? _T_10366_47 : _T_16094; // @[Mux.scala 46:16:@12021.4]
  assign _T_16097 = 6'h2f == _T_11317_54; // @[Mux.scala 46:19:@12022.4]
  assign _T_16098 = _T_16097 ? _T_10366_46 : _T_16096; // @[Mux.scala 46:16:@12023.4]
  assign _T_16099 = 6'h2e == _T_11317_54; // @[Mux.scala 46:19:@12024.4]
  assign _T_16100 = _T_16099 ? _T_10366_45 : _T_16098; // @[Mux.scala 46:16:@12025.4]
  assign _T_16101 = 6'h2d == _T_11317_54; // @[Mux.scala 46:19:@12026.4]
  assign _T_16102 = _T_16101 ? _T_10366_44 : _T_16100; // @[Mux.scala 46:16:@12027.4]
  assign _T_16103 = 6'h2c == _T_11317_54; // @[Mux.scala 46:19:@12028.4]
  assign _T_16104 = _T_16103 ? _T_10366_43 : _T_16102; // @[Mux.scala 46:16:@12029.4]
  assign _T_16105 = 6'h2b == _T_11317_54; // @[Mux.scala 46:19:@12030.4]
  assign _T_16106 = _T_16105 ? _T_10366_42 : _T_16104; // @[Mux.scala 46:16:@12031.4]
  assign _T_16107 = 6'h2a == _T_11317_54; // @[Mux.scala 46:19:@12032.4]
  assign _T_16108 = _T_16107 ? _T_10366_41 : _T_16106; // @[Mux.scala 46:16:@12033.4]
  assign _T_16109 = 6'h29 == _T_11317_54; // @[Mux.scala 46:19:@12034.4]
  assign _T_16110 = _T_16109 ? _T_10366_40 : _T_16108; // @[Mux.scala 46:16:@12035.4]
  assign _T_16111 = 6'h28 == _T_11317_54; // @[Mux.scala 46:19:@12036.4]
  assign _T_16112 = _T_16111 ? _T_10366_39 : _T_16110; // @[Mux.scala 46:16:@12037.4]
  assign _T_16113 = 6'h27 == _T_11317_54; // @[Mux.scala 46:19:@12038.4]
  assign _T_16114 = _T_16113 ? _T_10366_38 : _T_16112; // @[Mux.scala 46:16:@12039.4]
  assign _T_16115 = 6'h26 == _T_11317_54; // @[Mux.scala 46:19:@12040.4]
  assign _T_16116 = _T_16115 ? _T_10366_37 : _T_16114; // @[Mux.scala 46:16:@12041.4]
  assign _T_16117 = 6'h25 == _T_11317_54; // @[Mux.scala 46:19:@12042.4]
  assign _T_16118 = _T_16117 ? _T_10366_36 : _T_16116; // @[Mux.scala 46:16:@12043.4]
  assign _T_16119 = 6'h24 == _T_11317_54; // @[Mux.scala 46:19:@12044.4]
  assign _T_16120 = _T_16119 ? _T_10366_35 : _T_16118; // @[Mux.scala 46:16:@12045.4]
  assign _T_16121 = 6'h23 == _T_11317_54; // @[Mux.scala 46:19:@12046.4]
  assign _T_16122 = _T_16121 ? _T_10366_34 : _T_16120; // @[Mux.scala 46:16:@12047.4]
  assign _T_16123 = 6'h22 == _T_11317_54; // @[Mux.scala 46:19:@12048.4]
  assign _T_16124 = _T_16123 ? _T_10366_33 : _T_16122; // @[Mux.scala 46:16:@12049.4]
  assign _T_16125 = 6'h21 == _T_11317_54; // @[Mux.scala 46:19:@12050.4]
  assign _T_16126 = _T_16125 ? _T_10366_32 : _T_16124; // @[Mux.scala 46:16:@12051.4]
  assign _T_16127 = 6'h20 == _T_11317_54; // @[Mux.scala 46:19:@12052.4]
  assign _T_16128 = _T_16127 ? _T_10366_31 : _T_16126; // @[Mux.scala 46:16:@12053.4]
  assign _T_16129 = 6'h1f == _T_11317_54; // @[Mux.scala 46:19:@12054.4]
  assign _T_16130 = _T_16129 ? _T_10366_30 : _T_16128; // @[Mux.scala 46:16:@12055.4]
  assign _T_16131 = 6'h1e == _T_11317_54; // @[Mux.scala 46:19:@12056.4]
  assign _T_16132 = _T_16131 ? _T_10366_29 : _T_16130; // @[Mux.scala 46:16:@12057.4]
  assign _T_16133 = 6'h1d == _T_11317_54; // @[Mux.scala 46:19:@12058.4]
  assign _T_16134 = _T_16133 ? _T_10366_28 : _T_16132; // @[Mux.scala 46:16:@12059.4]
  assign _T_16135 = 6'h1c == _T_11317_54; // @[Mux.scala 46:19:@12060.4]
  assign _T_16136 = _T_16135 ? _T_10366_27 : _T_16134; // @[Mux.scala 46:16:@12061.4]
  assign _T_16137 = 6'h1b == _T_11317_54; // @[Mux.scala 46:19:@12062.4]
  assign _T_16138 = _T_16137 ? _T_10366_26 : _T_16136; // @[Mux.scala 46:16:@12063.4]
  assign _T_16139 = 6'h1a == _T_11317_54; // @[Mux.scala 46:19:@12064.4]
  assign _T_16140 = _T_16139 ? _T_10366_25 : _T_16138; // @[Mux.scala 46:16:@12065.4]
  assign _T_16141 = 6'h19 == _T_11317_54; // @[Mux.scala 46:19:@12066.4]
  assign _T_16142 = _T_16141 ? _T_10366_24 : _T_16140; // @[Mux.scala 46:16:@12067.4]
  assign _T_16143 = 6'h18 == _T_11317_54; // @[Mux.scala 46:19:@12068.4]
  assign _T_16144 = _T_16143 ? _T_10366_23 : _T_16142; // @[Mux.scala 46:16:@12069.4]
  assign _T_16145 = 6'h17 == _T_11317_54; // @[Mux.scala 46:19:@12070.4]
  assign _T_16146 = _T_16145 ? _T_10366_22 : _T_16144; // @[Mux.scala 46:16:@12071.4]
  assign _T_16147 = 6'h16 == _T_11317_54; // @[Mux.scala 46:19:@12072.4]
  assign _T_16148 = _T_16147 ? _T_10366_21 : _T_16146; // @[Mux.scala 46:16:@12073.4]
  assign _T_16149 = 6'h15 == _T_11317_54; // @[Mux.scala 46:19:@12074.4]
  assign _T_16150 = _T_16149 ? _T_10366_20 : _T_16148; // @[Mux.scala 46:16:@12075.4]
  assign _T_16151 = 6'h14 == _T_11317_54; // @[Mux.scala 46:19:@12076.4]
  assign _T_16152 = _T_16151 ? _T_10366_19 : _T_16150; // @[Mux.scala 46:16:@12077.4]
  assign _T_16153 = 6'h13 == _T_11317_54; // @[Mux.scala 46:19:@12078.4]
  assign _T_16154 = _T_16153 ? _T_10366_18 : _T_16152; // @[Mux.scala 46:16:@12079.4]
  assign _T_16155 = 6'h12 == _T_11317_54; // @[Mux.scala 46:19:@12080.4]
  assign _T_16156 = _T_16155 ? _T_10366_17 : _T_16154; // @[Mux.scala 46:16:@12081.4]
  assign _T_16157 = 6'h11 == _T_11317_54; // @[Mux.scala 46:19:@12082.4]
  assign _T_16158 = _T_16157 ? _T_10366_16 : _T_16156; // @[Mux.scala 46:16:@12083.4]
  assign _T_16159 = 6'h10 == _T_11317_54; // @[Mux.scala 46:19:@12084.4]
  assign _T_16160 = _T_16159 ? _T_10366_15 : _T_16158; // @[Mux.scala 46:16:@12085.4]
  assign _T_16161 = 6'hf == _T_11317_54; // @[Mux.scala 46:19:@12086.4]
  assign _T_16162 = _T_16161 ? _T_10366_14 : _T_16160; // @[Mux.scala 46:16:@12087.4]
  assign _T_16163 = 6'he == _T_11317_54; // @[Mux.scala 46:19:@12088.4]
  assign _T_16164 = _T_16163 ? _T_10366_13 : _T_16162; // @[Mux.scala 46:16:@12089.4]
  assign _T_16165 = 6'hd == _T_11317_54; // @[Mux.scala 46:19:@12090.4]
  assign _T_16166 = _T_16165 ? _T_10366_12 : _T_16164; // @[Mux.scala 46:16:@12091.4]
  assign _T_16167 = 6'hc == _T_11317_54; // @[Mux.scala 46:19:@12092.4]
  assign _T_16168 = _T_16167 ? _T_10366_11 : _T_16166; // @[Mux.scala 46:16:@12093.4]
  assign _T_16169 = 6'hb == _T_11317_54; // @[Mux.scala 46:19:@12094.4]
  assign _T_16170 = _T_16169 ? _T_10366_10 : _T_16168; // @[Mux.scala 46:16:@12095.4]
  assign _T_16171 = 6'ha == _T_11317_54; // @[Mux.scala 46:19:@12096.4]
  assign _T_16172 = _T_16171 ? _T_10366_9 : _T_16170; // @[Mux.scala 46:16:@12097.4]
  assign _T_16173 = 6'h9 == _T_11317_54; // @[Mux.scala 46:19:@12098.4]
  assign _T_16174 = _T_16173 ? _T_10366_8 : _T_16172; // @[Mux.scala 46:16:@12099.4]
  assign _T_16175 = 6'h8 == _T_11317_54; // @[Mux.scala 46:19:@12100.4]
  assign _T_16176 = _T_16175 ? _T_10366_7 : _T_16174; // @[Mux.scala 46:16:@12101.4]
  assign _T_16177 = 6'h7 == _T_11317_54; // @[Mux.scala 46:19:@12102.4]
  assign _T_16178 = _T_16177 ? _T_10366_6 : _T_16176; // @[Mux.scala 46:16:@12103.4]
  assign _T_16179 = 6'h6 == _T_11317_54; // @[Mux.scala 46:19:@12104.4]
  assign _T_16180 = _T_16179 ? _T_10366_5 : _T_16178; // @[Mux.scala 46:16:@12105.4]
  assign _T_16181 = 6'h5 == _T_11317_54; // @[Mux.scala 46:19:@12106.4]
  assign _T_16182 = _T_16181 ? _T_10366_4 : _T_16180; // @[Mux.scala 46:16:@12107.4]
  assign _T_16183 = 6'h4 == _T_11317_54; // @[Mux.scala 46:19:@12108.4]
  assign _T_16184 = _T_16183 ? _T_10366_3 : _T_16182; // @[Mux.scala 46:16:@12109.4]
  assign _T_16185 = 6'h3 == _T_11317_54; // @[Mux.scala 46:19:@12110.4]
  assign _T_16186 = _T_16185 ? _T_10366_2 : _T_16184; // @[Mux.scala 46:16:@12111.4]
  assign _T_16187 = 6'h2 == _T_11317_54; // @[Mux.scala 46:19:@12112.4]
  assign _T_16188 = _T_16187 ? _T_10366_1 : _T_16186; // @[Mux.scala 46:16:@12113.4]
  assign _T_16189 = 6'h1 == _T_11317_54; // @[Mux.scala 46:19:@12114.4]
  assign _T_16190 = _T_16189 ? _T_10366_0 : _T_16188; // @[Mux.scala 46:16:@12115.4]
  assign _T_16248 = 6'h38 == _T_11317_55; // @[Mux.scala 46:19:@12117.4]
  assign _T_16249 = _T_16248 ? _T_10366_55 : 8'h0; // @[Mux.scala 46:16:@12118.4]
  assign _T_16250 = 6'h37 == _T_11317_55; // @[Mux.scala 46:19:@12119.4]
  assign _T_16251 = _T_16250 ? _T_10366_54 : _T_16249; // @[Mux.scala 46:16:@12120.4]
  assign _T_16252 = 6'h36 == _T_11317_55; // @[Mux.scala 46:19:@12121.4]
  assign _T_16253 = _T_16252 ? _T_10366_53 : _T_16251; // @[Mux.scala 46:16:@12122.4]
  assign _T_16254 = 6'h35 == _T_11317_55; // @[Mux.scala 46:19:@12123.4]
  assign _T_16255 = _T_16254 ? _T_10366_52 : _T_16253; // @[Mux.scala 46:16:@12124.4]
  assign _T_16256 = 6'h34 == _T_11317_55; // @[Mux.scala 46:19:@12125.4]
  assign _T_16257 = _T_16256 ? _T_10366_51 : _T_16255; // @[Mux.scala 46:16:@12126.4]
  assign _T_16258 = 6'h33 == _T_11317_55; // @[Mux.scala 46:19:@12127.4]
  assign _T_16259 = _T_16258 ? _T_10366_50 : _T_16257; // @[Mux.scala 46:16:@12128.4]
  assign _T_16260 = 6'h32 == _T_11317_55; // @[Mux.scala 46:19:@12129.4]
  assign _T_16261 = _T_16260 ? _T_10366_49 : _T_16259; // @[Mux.scala 46:16:@12130.4]
  assign _T_16262 = 6'h31 == _T_11317_55; // @[Mux.scala 46:19:@12131.4]
  assign _T_16263 = _T_16262 ? _T_10366_48 : _T_16261; // @[Mux.scala 46:16:@12132.4]
  assign _T_16264 = 6'h30 == _T_11317_55; // @[Mux.scala 46:19:@12133.4]
  assign _T_16265 = _T_16264 ? _T_10366_47 : _T_16263; // @[Mux.scala 46:16:@12134.4]
  assign _T_16266 = 6'h2f == _T_11317_55; // @[Mux.scala 46:19:@12135.4]
  assign _T_16267 = _T_16266 ? _T_10366_46 : _T_16265; // @[Mux.scala 46:16:@12136.4]
  assign _T_16268 = 6'h2e == _T_11317_55; // @[Mux.scala 46:19:@12137.4]
  assign _T_16269 = _T_16268 ? _T_10366_45 : _T_16267; // @[Mux.scala 46:16:@12138.4]
  assign _T_16270 = 6'h2d == _T_11317_55; // @[Mux.scala 46:19:@12139.4]
  assign _T_16271 = _T_16270 ? _T_10366_44 : _T_16269; // @[Mux.scala 46:16:@12140.4]
  assign _T_16272 = 6'h2c == _T_11317_55; // @[Mux.scala 46:19:@12141.4]
  assign _T_16273 = _T_16272 ? _T_10366_43 : _T_16271; // @[Mux.scala 46:16:@12142.4]
  assign _T_16274 = 6'h2b == _T_11317_55; // @[Mux.scala 46:19:@12143.4]
  assign _T_16275 = _T_16274 ? _T_10366_42 : _T_16273; // @[Mux.scala 46:16:@12144.4]
  assign _T_16276 = 6'h2a == _T_11317_55; // @[Mux.scala 46:19:@12145.4]
  assign _T_16277 = _T_16276 ? _T_10366_41 : _T_16275; // @[Mux.scala 46:16:@12146.4]
  assign _T_16278 = 6'h29 == _T_11317_55; // @[Mux.scala 46:19:@12147.4]
  assign _T_16279 = _T_16278 ? _T_10366_40 : _T_16277; // @[Mux.scala 46:16:@12148.4]
  assign _T_16280 = 6'h28 == _T_11317_55; // @[Mux.scala 46:19:@12149.4]
  assign _T_16281 = _T_16280 ? _T_10366_39 : _T_16279; // @[Mux.scala 46:16:@12150.4]
  assign _T_16282 = 6'h27 == _T_11317_55; // @[Mux.scala 46:19:@12151.4]
  assign _T_16283 = _T_16282 ? _T_10366_38 : _T_16281; // @[Mux.scala 46:16:@12152.4]
  assign _T_16284 = 6'h26 == _T_11317_55; // @[Mux.scala 46:19:@12153.4]
  assign _T_16285 = _T_16284 ? _T_10366_37 : _T_16283; // @[Mux.scala 46:16:@12154.4]
  assign _T_16286 = 6'h25 == _T_11317_55; // @[Mux.scala 46:19:@12155.4]
  assign _T_16287 = _T_16286 ? _T_10366_36 : _T_16285; // @[Mux.scala 46:16:@12156.4]
  assign _T_16288 = 6'h24 == _T_11317_55; // @[Mux.scala 46:19:@12157.4]
  assign _T_16289 = _T_16288 ? _T_10366_35 : _T_16287; // @[Mux.scala 46:16:@12158.4]
  assign _T_16290 = 6'h23 == _T_11317_55; // @[Mux.scala 46:19:@12159.4]
  assign _T_16291 = _T_16290 ? _T_10366_34 : _T_16289; // @[Mux.scala 46:16:@12160.4]
  assign _T_16292 = 6'h22 == _T_11317_55; // @[Mux.scala 46:19:@12161.4]
  assign _T_16293 = _T_16292 ? _T_10366_33 : _T_16291; // @[Mux.scala 46:16:@12162.4]
  assign _T_16294 = 6'h21 == _T_11317_55; // @[Mux.scala 46:19:@12163.4]
  assign _T_16295 = _T_16294 ? _T_10366_32 : _T_16293; // @[Mux.scala 46:16:@12164.4]
  assign _T_16296 = 6'h20 == _T_11317_55; // @[Mux.scala 46:19:@12165.4]
  assign _T_16297 = _T_16296 ? _T_10366_31 : _T_16295; // @[Mux.scala 46:16:@12166.4]
  assign _T_16298 = 6'h1f == _T_11317_55; // @[Mux.scala 46:19:@12167.4]
  assign _T_16299 = _T_16298 ? _T_10366_30 : _T_16297; // @[Mux.scala 46:16:@12168.4]
  assign _T_16300 = 6'h1e == _T_11317_55; // @[Mux.scala 46:19:@12169.4]
  assign _T_16301 = _T_16300 ? _T_10366_29 : _T_16299; // @[Mux.scala 46:16:@12170.4]
  assign _T_16302 = 6'h1d == _T_11317_55; // @[Mux.scala 46:19:@12171.4]
  assign _T_16303 = _T_16302 ? _T_10366_28 : _T_16301; // @[Mux.scala 46:16:@12172.4]
  assign _T_16304 = 6'h1c == _T_11317_55; // @[Mux.scala 46:19:@12173.4]
  assign _T_16305 = _T_16304 ? _T_10366_27 : _T_16303; // @[Mux.scala 46:16:@12174.4]
  assign _T_16306 = 6'h1b == _T_11317_55; // @[Mux.scala 46:19:@12175.4]
  assign _T_16307 = _T_16306 ? _T_10366_26 : _T_16305; // @[Mux.scala 46:16:@12176.4]
  assign _T_16308 = 6'h1a == _T_11317_55; // @[Mux.scala 46:19:@12177.4]
  assign _T_16309 = _T_16308 ? _T_10366_25 : _T_16307; // @[Mux.scala 46:16:@12178.4]
  assign _T_16310 = 6'h19 == _T_11317_55; // @[Mux.scala 46:19:@12179.4]
  assign _T_16311 = _T_16310 ? _T_10366_24 : _T_16309; // @[Mux.scala 46:16:@12180.4]
  assign _T_16312 = 6'h18 == _T_11317_55; // @[Mux.scala 46:19:@12181.4]
  assign _T_16313 = _T_16312 ? _T_10366_23 : _T_16311; // @[Mux.scala 46:16:@12182.4]
  assign _T_16314 = 6'h17 == _T_11317_55; // @[Mux.scala 46:19:@12183.4]
  assign _T_16315 = _T_16314 ? _T_10366_22 : _T_16313; // @[Mux.scala 46:16:@12184.4]
  assign _T_16316 = 6'h16 == _T_11317_55; // @[Mux.scala 46:19:@12185.4]
  assign _T_16317 = _T_16316 ? _T_10366_21 : _T_16315; // @[Mux.scala 46:16:@12186.4]
  assign _T_16318 = 6'h15 == _T_11317_55; // @[Mux.scala 46:19:@12187.4]
  assign _T_16319 = _T_16318 ? _T_10366_20 : _T_16317; // @[Mux.scala 46:16:@12188.4]
  assign _T_16320 = 6'h14 == _T_11317_55; // @[Mux.scala 46:19:@12189.4]
  assign _T_16321 = _T_16320 ? _T_10366_19 : _T_16319; // @[Mux.scala 46:16:@12190.4]
  assign _T_16322 = 6'h13 == _T_11317_55; // @[Mux.scala 46:19:@12191.4]
  assign _T_16323 = _T_16322 ? _T_10366_18 : _T_16321; // @[Mux.scala 46:16:@12192.4]
  assign _T_16324 = 6'h12 == _T_11317_55; // @[Mux.scala 46:19:@12193.4]
  assign _T_16325 = _T_16324 ? _T_10366_17 : _T_16323; // @[Mux.scala 46:16:@12194.4]
  assign _T_16326 = 6'h11 == _T_11317_55; // @[Mux.scala 46:19:@12195.4]
  assign _T_16327 = _T_16326 ? _T_10366_16 : _T_16325; // @[Mux.scala 46:16:@12196.4]
  assign _T_16328 = 6'h10 == _T_11317_55; // @[Mux.scala 46:19:@12197.4]
  assign _T_16329 = _T_16328 ? _T_10366_15 : _T_16327; // @[Mux.scala 46:16:@12198.4]
  assign _T_16330 = 6'hf == _T_11317_55; // @[Mux.scala 46:19:@12199.4]
  assign _T_16331 = _T_16330 ? _T_10366_14 : _T_16329; // @[Mux.scala 46:16:@12200.4]
  assign _T_16332 = 6'he == _T_11317_55; // @[Mux.scala 46:19:@12201.4]
  assign _T_16333 = _T_16332 ? _T_10366_13 : _T_16331; // @[Mux.scala 46:16:@12202.4]
  assign _T_16334 = 6'hd == _T_11317_55; // @[Mux.scala 46:19:@12203.4]
  assign _T_16335 = _T_16334 ? _T_10366_12 : _T_16333; // @[Mux.scala 46:16:@12204.4]
  assign _T_16336 = 6'hc == _T_11317_55; // @[Mux.scala 46:19:@12205.4]
  assign _T_16337 = _T_16336 ? _T_10366_11 : _T_16335; // @[Mux.scala 46:16:@12206.4]
  assign _T_16338 = 6'hb == _T_11317_55; // @[Mux.scala 46:19:@12207.4]
  assign _T_16339 = _T_16338 ? _T_10366_10 : _T_16337; // @[Mux.scala 46:16:@12208.4]
  assign _T_16340 = 6'ha == _T_11317_55; // @[Mux.scala 46:19:@12209.4]
  assign _T_16341 = _T_16340 ? _T_10366_9 : _T_16339; // @[Mux.scala 46:16:@12210.4]
  assign _T_16342 = 6'h9 == _T_11317_55; // @[Mux.scala 46:19:@12211.4]
  assign _T_16343 = _T_16342 ? _T_10366_8 : _T_16341; // @[Mux.scala 46:16:@12212.4]
  assign _T_16344 = 6'h8 == _T_11317_55; // @[Mux.scala 46:19:@12213.4]
  assign _T_16345 = _T_16344 ? _T_10366_7 : _T_16343; // @[Mux.scala 46:16:@12214.4]
  assign _T_16346 = 6'h7 == _T_11317_55; // @[Mux.scala 46:19:@12215.4]
  assign _T_16347 = _T_16346 ? _T_10366_6 : _T_16345; // @[Mux.scala 46:16:@12216.4]
  assign _T_16348 = 6'h6 == _T_11317_55; // @[Mux.scala 46:19:@12217.4]
  assign _T_16349 = _T_16348 ? _T_10366_5 : _T_16347; // @[Mux.scala 46:16:@12218.4]
  assign _T_16350 = 6'h5 == _T_11317_55; // @[Mux.scala 46:19:@12219.4]
  assign _T_16351 = _T_16350 ? _T_10366_4 : _T_16349; // @[Mux.scala 46:16:@12220.4]
  assign _T_16352 = 6'h4 == _T_11317_55; // @[Mux.scala 46:19:@12221.4]
  assign _T_16353 = _T_16352 ? _T_10366_3 : _T_16351; // @[Mux.scala 46:16:@12222.4]
  assign _T_16354 = 6'h3 == _T_11317_55; // @[Mux.scala 46:19:@12223.4]
  assign _T_16355 = _T_16354 ? _T_10366_2 : _T_16353; // @[Mux.scala 46:16:@12224.4]
  assign _T_16356 = 6'h2 == _T_11317_55; // @[Mux.scala 46:19:@12225.4]
  assign _T_16357 = _T_16356 ? _T_10366_1 : _T_16355; // @[Mux.scala 46:16:@12226.4]
  assign _T_16358 = 6'h1 == _T_11317_55; // @[Mux.scala 46:19:@12227.4]
  assign _T_16359 = _T_16358 ? _T_10366_0 : _T_16357; // @[Mux.scala 46:16:@12228.4]
  assign _T_16418 = 6'h39 == _T_11317_56; // @[Mux.scala 46:19:@12230.4]
  assign _T_16419 = _T_16418 ? _T_10366_56 : 8'h0; // @[Mux.scala 46:16:@12231.4]
  assign _T_16420 = 6'h38 == _T_11317_56; // @[Mux.scala 46:19:@12232.4]
  assign _T_16421 = _T_16420 ? _T_10366_55 : _T_16419; // @[Mux.scala 46:16:@12233.4]
  assign _T_16422 = 6'h37 == _T_11317_56; // @[Mux.scala 46:19:@12234.4]
  assign _T_16423 = _T_16422 ? _T_10366_54 : _T_16421; // @[Mux.scala 46:16:@12235.4]
  assign _T_16424 = 6'h36 == _T_11317_56; // @[Mux.scala 46:19:@12236.4]
  assign _T_16425 = _T_16424 ? _T_10366_53 : _T_16423; // @[Mux.scala 46:16:@12237.4]
  assign _T_16426 = 6'h35 == _T_11317_56; // @[Mux.scala 46:19:@12238.4]
  assign _T_16427 = _T_16426 ? _T_10366_52 : _T_16425; // @[Mux.scala 46:16:@12239.4]
  assign _T_16428 = 6'h34 == _T_11317_56; // @[Mux.scala 46:19:@12240.4]
  assign _T_16429 = _T_16428 ? _T_10366_51 : _T_16427; // @[Mux.scala 46:16:@12241.4]
  assign _T_16430 = 6'h33 == _T_11317_56; // @[Mux.scala 46:19:@12242.4]
  assign _T_16431 = _T_16430 ? _T_10366_50 : _T_16429; // @[Mux.scala 46:16:@12243.4]
  assign _T_16432 = 6'h32 == _T_11317_56; // @[Mux.scala 46:19:@12244.4]
  assign _T_16433 = _T_16432 ? _T_10366_49 : _T_16431; // @[Mux.scala 46:16:@12245.4]
  assign _T_16434 = 6'h31 == _T_11317_56; // @[Mux.scala 46:19:@12246.4]
  assign _T_16435 = _T_16434 ? _T_10366_48 : _T_16433; // @[Mux.scala 46:16:@12247.4]
  assign _T_16436 = 6'h30 == _T_11317_56; // @[Mux.scala 46:19:@12248.4]
  assign _T_16437 = _T_16436 ? _T_10366_47 : _T_16435; // @[Mux.scala 46:16:@12249.4]
  assign _T_16438 = 6'h2f == _T_11317_56; // @[Mux.scala 46:19:@12250.4]
  assign _T_16439 = _T_16438 ? _T_10366_46 : _T_16437; // @[Mux.scala 46:16:@12251.4]
  assign _T_16440 = 6'h2e == _T_11317_56; // @[Mux.scala 46:19:@12252.4]
  assign _T_16441 = _T_16440 ? _T_10366_45 : _T_16439; // @[Mux.scala 46:16:@12253.4]
  assign _T_16442 = 6'h2d == _T_11317_56; // @[Mux.scala 46:19:@12254.4]
  assign _T_16443 = _T_16442 ? _T_10366_44 : _T_16441; // @[Mux.scala 46:16:@12255.4]
  assign _T_16444 = 6'h2c == _T_11317_56; // @[Mux.scala 46:19:@12256.4]
  assign _T_16445 = _T_16444 ? _T_10366_43 : _T_16443; // @[Mux.scala 46:16:@12257.4]
  assign _T_16446 = 6'h2b == _T_11317_56; // @[Mux.scala 46:19:@12258.4]
  assign _T_16447 = _T_16446 ? _T_10366_42 : _T_16445; // @[Mux.scala 46:16:@12259.4]
  assign _T_16448 = 6'h2a == _T_11317_56; // @[Mux.scala 46:19:@12260.4]
  assign _T_16449 = _T_16448 ? _T_10366_41 : _T_16447; // @[Mux.scala 46:16:@12261.4]
  assign _T_16450 = 6'h29 == _T_11317_56; // @[Mux.scala 46:19:@12262.4]
  assign _T_16451 = _T_16450 ? _T_10366_40 : _T_16449; // @[Mux.scala 46:16:@12263.4]
  assign _T_16452 = 6'h28 == _T_11317_56; // @[Mux.scala 46:19:@12264.4]
  assign _T_16453 = _T_16452 ? _T_10366_39 : _T_16451; // @[Mux.scala 46:16:@12265.4]
  assign _T_16454 = 6'h27 == _T_11317_56; // @[Mux.scala 46:19:@12266.4]
  assign _T_16455 = _T_16454 ? _T_10366_38 : _T_16453; // @[Mux.scala 46:16:@12267.4]
  assign _T_16456 = 6'h26 == _T_11317_56; // @[Mux.scala 46:19:@12268.4]
  assign _T_16457 = _T_16456 ? _T_10366_37 : _T_16455; // @[Mux.scala 46:16:@12269.4]
  assign _T_16458 = 6'h25 == _T_11317_56; // @[Mux.scala 46:19:@12270.4]
  assign _T_16459 = _T_16458 ? _T_10366_36 : _T_16457; // @[Mux.scala 46:16:@12271.4]
  assign _T_16460 = 6'h24 == _T_11317_56; // @[Mux.scala 46:19:@12272.4]
  assign _T_16461 = _T_16460 ? _T_10366_35 : _T_16459; // @[Mux.scala 46:16:@12273.4]
  assign _T_16462 = 6'h23 == _T_11317_56; // @[Mux.scala 46:19:@12274.4]
  assign _T_16463 = _T_16462 ? _T_10366_34 : _T_16461; // @[Mux.scala 46:16:@12275.4]
  assign _T_16464 = 6'h22 == _T_11317_56; // @[Mux.scala 46:19:@12276.4]
  assign _T_16465 = _T_16464 ? _T_10366_33 : _T_16463; // @[Mux.scala 46:16:@12277.4]
  assign _T_16466 = 6'h21 == _T_11317_56; // @[Mux.scala 46:19:@12278.4]
  assign _T_16467 = _T_16466 ? _T_10366_32 : _T_16465; // @[Mux.scala 46:16:@12279.4]
  assign _T_16468 = 6'h20 == _T_11317_56; // @[Mux.scala 46:19:@12280.4]
  assign _T_16469 = _T_16468 ? _T_10366_31 : _T_16467; // @[Mux.scala 46:16:@12281.4]
  assign _T_16470 = 6'h1f == _T_11317_56; // @[Mux.scala 46:19:@12282.4]
  assign _T_16471 = _T_16470 ? _T_10366_30 : _T_16469; // @[Mux.scala 46:16:@12283.4]
  assign _T_16472 = 6'h1e == _T_11317_56; // @[Mux.scala 46:19:@12284.4]
  assign _T_16473 = _T_16472 ? _T_10366_29 : _T_16471; // @[Mux.scala 46:16:@12285.4]
  assign _T_16474 = 6'h1d == _T_11317_56; // @[Mux.scala 46:19:@12286.4]
  assign _T_16475 = _T_16474 ? _T_10366_28 : _T_16473; // @[Mux.scala 46:16:@12287.4]
  assign _T_16476 = 6'h1c == _T_11317_56; // @[Mux.scala 46:19:@12288.4]
  assign _T_16477 = _T_16476 ? _T_10366_27 : _T_16475; // @[Mux.scala 46:16:@12289.4]
  assign _T_16478 = 6'h1b == _T_11317_56; // @[Mux.scala 46:19:@12290.4]
  assign _T_16479 = _T_16478 ? _T_10366_26 : _T_16477; // @[Mux.scala 46:16:@12291.4]
  assign _T_16480 = 6'h1a == _T_11317_56; // @[Mux.scala 46:19:@12292.4]
  assign _T_16481 = _T_16480 ? _T_10366_25 : _T_16479; // @[Mux.scala 46:16:@12293.4]
  assign _T_16482 = 6'h19 == _T_11317_56; // @[Mux.scala 46:19:@12294.4]
  assign _T_16483 = _T_16482 ? _T_10366_24 : _T_16481; // @[Mux.scala 46:16:@12295.4]
  assign _T_16484 = 6'h18 == _T_11317_56; // @[Mux.scala 46:19:@12296.4]
  assign _T_16485 = _T_16484 ? _T_10366_23 : _T_16483; // @[Mux.scala 46:16:@12297.4]
  assign _T_16486 = 6'h17 == _T_11317_56; // @[Mux.scala 46:19:@12298.4]
  assign _T_16487 = _T_16486 ? _T_10366_22 : _T_16485; // @[Mux.scala 46:16:@12299.4]
  assign _T_16488 = 6'h16 == _T_11317_56; // @[Mux.scala 46:19:@12300.4]
  assign _T_16489 = _T_16488 ? _T_10366_21 : _T_16487; // @[Mux.scala 46:16:@12301.4]
  assign _T_16490 = 6'h15 == _T_11317_56; // @[Mux.scala 46:19:@12302.4]
  assign _T_16491 = _T_16490 ? _T_10366_20 : _T_16489; // @[Mux.scala 46:16:@12303.4]
  assign _T_16492 = 6'h14 == _T_11317_56; // @[Mux.scala 46:19:@12304.4]
  assign _T_16493 = _T_16492 ? _T_10366_19 : _T_16491; // @[Mux.scala 46:16:@12305.4]
  assign _T_16494 = 6'h13 == _T_11317_56; // @[Mux.scala 46:19:@12306.4]
  assign _T_16495 = _T_16494 ? _T_10366_18 : _T_16493; // @[Mux.scala 46:16:@12307.4]
  assign _T_16496 = 6'h12 == _T_11317_56; // @[Mux.scala 46:19:@12308.4]
  assign _T_16497 = _T_16496 ? _T_10366_17 : _T_16495; // @[Mux.scala 46:16:@12309.4]
  assign _T_16498 = 6'h11 == _T_11317_56; // @[Mux.scala 46:19:@12310.4]
  assign _T_16499 = _T_16498 ? _T_10366_16 : _T_16497; // @[Mux.scala 46:16:@12311.4]
  assign _T_16500 = 6'h10 == _T_11317_56; // @[Mux.scala 46:19:@12312.4]
  assign _T_16501 = _T_16500 ? _T_10366_15 : _T_16499; // @[Mux.scala 46:16:@12313.4]
  assign _T_16502 = 6'hf == _T_11317_56; // @[Mux.scala 46:19:@12314.4]
  assign _T_16503 = _T_16502 ? _T_10366_14 : _T_16501; // @[Mux.scala 46:16:@12315.4]
  assign _T_16504 = 6'he == _T_11317_56; // @[Mux.scala 46:19:@12316.4]
  assign _T_16505 = _T_16504 ? _T_10366_13 : _T_16503; // @[Mux.scala 46:16:@12317.4]
  assign _T_16506 = 6'hd == _T_11317_56; // @[Mux.scala 46:19:@12318.4]
  assign _T_16507 = _T_16506 ? _T_10366_12 : _T_16505; // @[Mux.scala 46:16:@12319.4]
  assign _T_16508 = 6'hc == _T_11317_56; // @[Mux.scala 46:19:@12320.4]
  assign _T_16509 = _T_16508 ? _T_10366_11 : _T_16507; // @[Mux.scala 46:16:@12321.4]
  assign _T_16510 = 6'hb == _T_11317_56; // @[Mux.scala 46:19:@12322.4]
  assign _T_16511 = _T_16510 ? _T_10366_10 : _T_16509; // @[Mux.scala 46:16:@12323.4]
  assign _T_16512 = 6'ha == _T_11317_56; // @[Mux.scala 46:19:@12324.4]
  assign _T_16513 = _T_16512 ? _T_10366_9 : _T_16511; // @[Mux.scala 46:16:@12325.4]
  assign _T_16514 = 6'h9 == _T_11317_56; // @[Mux.scala 46:19:@12326.4]
  assign _T_16515 = _T_16514 ? _T_10366_8 : _T_16513; // @[Mux.scala 46:16:@12327.4]
  assign _T_16516 = 6'h8 == _T_11317_56; // @[Mux.scala 46:19:@12328.4]
  assign _T_16517 = _T_16516 ? _T_10366_7 : _T_16515; // @[Mux.scala 46:16:@12329.4]
  assign _T_16518 = 6'h7 == _T_11317_56; // @[Mux.scala 46:19:@12330.4]
  assign _T_16519 = _T_16518 ? _T_10366_6 : _T_16517; // @[Mux.scala 46:16:@12331.4]
  assign _T_16520 = 6'h6 == _T_11317_56; // @[Mux.scala 46:19:@12332.4]
  assign _T_16521 = _T_16520 ? _T_10366_5 : _T_16519; // @[Mux.scala 46:16:@12333.4]
  assign _T_16522 = 6'h5 == _T_11317_56; // @[Mux.scala 46:19:@12334.4]
  assign _T_16523 = _T_16522 ? _T_10366_4 : _T_16521; // @[Mux.scala 46:16:@12335.4]
  assign _T_16524 = 6'h4 == _T_11317_56; // @[Mux.scala 46:19:@12336.4]
  assign _T_16525 = _T_16524 ? _T_10366_3 : _T_16523; // @[Mux.scala 46:16:@12337.4]
  assign _T_16526 = 6'h3 == _T_11317_56; // @[Mux.scala 46:19:@12338.4]
  assign _T_16527 = _T_16526 ? _T_10366_2 : _T_16525; // @[Mux.scala 46:16:@12339.4]
  assign _T_16528 = 6'h2 == _T_11317_56; // @[Mux.scala 46:19:@12340.4]
  assign _T_16529 = _T_16528 ? _T_10366_1 : _T_16527; // @[Mux.scala 46:16:@12341.4]
  assign _T_16530 = 6'h1 == _T_11317_56; // @[Mux.scala 46:19:@12342.4]
  assign _T_16531 = _T_16530 ? _T_10366_0 : _T_16529; // @[Mux.scala 46:16:@12343.4]
  assign _T_16591 = 6'h3a == _T_11317_57; // @[Mux.scala 46:19:@12345.4]
  assign _T_16592 = _T_16591 ? _T_10366_57 : 8'h0; // @[Mux.scala 46:16:@12346.4]
  assign _T_16593 = 6'h39 == _T_11317_57; // @[Mux.scala 46:19:@12347.4]
  assign _T_16594 = _T_16593 ? _T_10366_56 : _T_16592; // @[Mux.scala 46:16:@12348.4]
  assign _T_16595 = 6'h38 == _T_11317_57; // @[Mux.scala 46:19:@12349.4]
  assign _T_16596 = _T_16595 ? _T_10366_55 : _T_16594; // @[Mux.scala 46:16:@12350.4]
  assign _T_16597 = 6'h37 == _T_11317_57; // @[Mux.scala 46:19:@12351.4]
  assign _T_16598 = _T_16597 ? _T_10366_54 : _T_16596; // @[Mux.scala 46:16:@12352.4]
  assign _T_16599 = 6'h36 == _T_11317_57; // @[Mux.scala 46:19:@12353.4]
  assign _T_16600 = _T_16599 ? _T_10366_53 : _T_16598; // @[Mux.scala 46:16:@12354.4]
  assign _T_16601 = 6'h35 == _T_11317_57; // @[Mux.scala 46:19:@12355.4]
  assign _T_16602 = _T_16601 ? _T_10366_52 : _T_16600; // @[Mux.scala 46:16:@12356.4]
  assign _T_16603 = 6'h34 == _T_11317_57; // @[Mux.scala 46:19:@12357.4]
  assign _T_16604 = _T_16603 ? _T_10366_51 : _T_16602; // @[Mux.scala 46:16:@12358.4]
  assign _T_16605 = 6'h33 == _T_11317_57; // @[Mux.scala 46:19:@12359.4]
  assign _T_16606 = _T_16605 ? _T_10366_50 : _T_16604; // @[Mux.scala 46:16:@12360.4]
  assign _T_16607 = 6'h32 == _T_11317_57; // @[Mux.scala 46:19:@12361.4]
  assign _T_16608 = _T_16607 ? _T_10366_49 : _T_16606; // @[Mux.scala 46:16:@12362.4]
  assign _T_16609 = 6'h31 == _T_11317_57; // @[Mux.scala 46:19:@12363.4]
  assign _T_16610 = _T_16609 ? _T_10366_48 : _T_16608; // @[Mux.scala 46:16:@12364.4]
  assign _T_16611 = 6'h30 == _T_11317_57; // @[Mux.scala 46:19:@12365.4]
  assign _T_16612 = _T_16611 ? _T_10366_47 : _T_16610; // @[Mux.scala 46:16:@12366.4]
  assign _T_16613 = 6'h2f == _T_11317_57; // @[Mux.scala 46:19:@12367.4]
  assign _T_16614 = _T_16613 ? _T_10366_46 : _T_16612; // @[Mux.scala 46:16:@12368.4]
  assign _T_16615 = 6'h2e == _T_11317_57; // @[Mux.scala 46:19:@12369.4]
  assign _T_16616 = _T_16615 ? _T_10366_45 : _T_16614; // @[Mux.scala 46:16:@12370.4]
  assign _T_16617 = 6'h2d == _T_11317_57; // @[Mux.scala 46:19:@12371.4]
  assign _T_16618 = _T_16617 ? _T_10366_44 : _T_16616; // @[Mux.scala 46:16:@12372.4]
  assign _T_16619 = 6'h2c == _T_11317_57; // @[Mux.scala 46:19:@12373.4]
  assign _T_16620 = _T_16619 ? _T_10366_43 : _T_16618; // @[Mux.scala 46:16:@12374.4]
  assign _T_16621 = 6'h2b == _T_11317_57; // @[Mux.scala 46:19:@12375.4]
  assign _T_16622 = _T_16621 ? _T_10366_42 : _T_16620; // @[Mux.scala 46:16:@12376.4]
  assign _T_16623 = 6'h2a == _T_11317_57; // @[Mux.scala 46:19:@12377.4]
  assign _T_16624 = _T_16623 ? _T_10366_41 : _T_16622; // @[Mux.scala 46:16:@12378.4]
  assign _T_16625 = 6'h29 == _T_11317_57; // @[Mux.scala 46:19:@12379.4]
  assign _T_16626 = _T_16625 ? _T_10366_40 : _T_16624; // @[Mux.scala 46:16:@12380.4]
  assign _T_16627 = 6'h28 == _T_11317_57; // @[Mux.scala 46:19:@12381.4]
  assign _T_16628 = _T_16627 ? _T_10366_39 : _T_16626; // @[Mux.scala 46:16:@12382.4]
  assign _T_16629 = 6'h27 == _T_11317_57; // @[Mux.scala 46:19:@12383.4]
  assign _T_16630 = _T_16629 ? _T_10366_38 : _T_16628; // @[Mux.scala 46:16:@12384.4]
  assign _T_16631 = 6'h26 == _T_11317_57; // @[Mux.scala 46:19:@12385.4]
  assign _T_16632 = _T_16631 ? _T_10366_37 : _T_16630; // @[Mux.scala 46:16:@12386.4]
  assign _T_16633 = 6'h25 == _T_11317_57; // @[Mux.scala 46:19:@12387.4]
  assign _T_16634 = _T_16633 ? _T_10366_36 : _T_16632; // @[Mux.scala 46:16:@12388.4]
  assign _T_16635 = 6'h24 == _T_11317_57; // @[Mux.scala 46:19:@12389.4]
  assign _T_16636 = _T_16635 ? _T_10366_35 : _T_16634; // @[Mux.scala 46:16:@12390.4]
  assign _T_16637 = 6'h23 == _T_11317_57; // @[Mux.scala 46:19:@12391.4]
  assign _T_16638 = _T_16637 ? _T_10366_34 : _T_16636; // @[Mux.scala 46:16:@12392.4]
  assign _T_16639 = 6'h22 == _T_11317_57; // @[Mux.scala 46:19:@12393.4]
  assign _T_16640 = _T_16639 ? _T_10366_33 : _T_16638; // @[Mux.scala 46:16:@12394.4]
  assign _T_16641 = 6'h21 == _T_11317_57; // @[Mux.scala 46:19:@12395.4]
  assign _T_16642 = _T_16641 ? _T_10366_32 : _T_16640; // @[Mux.scala 46:16:@12396.4]
  assign _T_16643 = 6'h20 == _T_11317_57; // @[Mux.scala 46:19:@12397.4]
  assign _T_16644 = _T_16643 ? _T_10366_31 : _T_16642; // @[Mux.scala 46:16:@12398.4]
  assign _T_16645 = 6'h1f == _T_11317_57; // @[Mux.scala 46:19:@12399.4]
  assign _T_16646 = _T_16645 ? _T_10366_30 : _T_16644; // @[Mux.scala 46:16:@12400.4]
  assign _T_16647 = 6'h1e == _T_11317_57; // @[Mux.scala 46:19:@12401.4]
  assign _T_16648 = _T_16647 ? _T_10366_29 : _T_16646; // @[Mux.scala 46:16:@12402.4]
  assign _T_16649 = 6'h1d == _T_11317_57; // @[Mux.scala 46:19:@12403.4]
  assign _T_16650 = _T_16649 ? _T_10366_28 : _T_16648; // @[Mux.scala 46:16:@12404.4]
  assign _T_16651 = 6'h1c == _T_11317_57; // @[Mux.scala 46:19:@12405.4]
  assign _T_16652 = _T_16651 ? _T_10366_27 : _T_16650; // @[Mux.scala 46:16:@12406.4]
  assign _T_16653 = 6'h1b == _T_11317_57; // @[Mux.scala 46:19:@12407.4]
  assign _T_16654 = _T_16653 ? _T_10366_26 : _T_16652; // @[Mux.scala 46:16:@12408.4]
  assign _T_16655 = 6'h1a == _T_11317_57; // @[Mux.scala 46:19:@12409.4]
  assign _T_16656 = _T_16655 ? _T_10366_25 : _T_16654; // @[Mux.scala 46:16:@12410.4]
  assign _T_16657 = 6'h19 == _T_11317_57; // @[Mux.scala 46:19:@12411.4]
  assign _T_16658 = _T_16657 ? _T_10366_24 : _T_16656; // @[Mux.scala 46:16:@12412.4]
  assign _T_16659 = 6'h18 == _T_11317_57; // @[Mux.scala 46:19:@12413.4]
  assign _T_16660 = _T_16659 ? _T_10366_23 : _T_16658; // @[Mux.scala 46:16:@12414.4]
  assign _T_16661 = 6'h17 == _T_11317_57; // @[Mux.scala 46:19:@12415.4]
  assign _T_16662 = _T_16661 ? _T_10366_22 : _T_16660; // @[Mux.scala 46:16:@12416.4]
  assign _T_16663 = 6'h16 == _T_11317_57; // @[Mux.scala 46:19:@12417.4]
  assign _T_16664 = _T_16663 ? _T_10366_21 : _T_16662; // @[Mux.scala 46:16:@12418.4]
  assign _T_16665 = 6'h15 == _T_11317_57; // @[Mux.scala 46:19:@12419.4]
  assign _T_16666 = _T_16665 ? _T_10366_20 : _T_16664; // @[Mux.scala 46:16:@12420.4]
  assign _T_16667 = 6'h14 == _T_11317_57; // @[Mux.scala 46:19:@12421.4]
  assign _T_16668 = _T_16667 ? _T_10366_19 : _T_16666; // @[Mux.scala 46:16:@12422.4]
  assign _T_16669 = 6'h13 == _T_11317_57; // @[Mux.scala 46:19:@12423.4]
  assign _T_16670 = _T_16669 ? _T_10366_18 : _T_16668; // @[Mux.scala 46:16:@12424.4]
  assign _T_16671 = 6'h12 == _T_11317_57; // @[Mux.scala 46:19:@12425.4]
  assign _T_16672 = _T_16671 ? _T_10366_17 : _T_16670; // @[Mux.scala 46:16:@12426.4]
  assign _T_16673 = 6'h11 == _T_11317_57; // @[Mux.scala 46:19:@12427.4]
  assign _T_16674 = _T_16673 ? _T_10366_16 : _T_16672; // @[Mux.scala 46:16:@12428.4]
  assign _T_16675 = 6'h10 == _T_11317_57; // @[Mux.scala 46:19:@12429.4]
  assign _T_16676 = _T_16675 ? _T_10366_15 : _T_16674; // @[Mux.scala 46:16:@12430.4]
  assign _T_16677 = 6'hf == _T_11317_57; // @[Mux.scala 46:19:@12431.4]
  assign _T_16678 = _T_16677 ? _T_10366_14 : _T_16676; // @[Mux.scala 46:16:@12432.4]
  assign _T_16679 = 6'he == _T_11317_57; // @[Mux.scala 46:19:@12433.4]
  assign _T_16680 = _T_16679 ? _T_10366_13 : _T_16678; // @[Mux.scala 46:16:@12434.4]
  assign _T_16681 = 6'hd == _T_11317_57; // @[Mux.scala 46:19:@12435.4]
  assign _T_16682 = _T_16681 ? _T_10366_12 : _T_16680; // @[Mux.scala 46:16:@12436.4]
  assign _T_16683 = 6'hc == _T_11317_57; // @[Mux.scala 46:19:@12437.4]
  assign _T_16684 = _T_16683 ? _T_10366_11 : _T_16682; // @[Mux.scala 46:16:@12438.4]
  assign _T_16685 = 6'hb == _T_11317_57; // @[Mux.scala 46:19:@12439.4]
  assign _T_16686 = _T_16685 ? _T_10366_10 : _T_16684; // @[Mux.scala 46:16:@12440.4]
  assign _T_16687 = 6'ha == _T_11317_57; // @[Mux.scala 46:19:@12441.4]
  assign _T_16688 = _T_16687 ? _T_10366_9 : _T_16686; // @[Mux.scala 46:16:@12442.4]
  assign _T_16689 = 6'h9 == _T_11317_57; // @[Mux.scala 46:19:@12443.4]
  assign _T_16690 = _T_16689 ? _T_10366_8 : _T_16688; // @[Mux.scala 46:16:@12444.4]
  assign _T_16691 = 6'h8 == _T_11317_57; // @[Mux.scala 46:19:@12445.4]
  assign _T_16692 = _T_16691 ? _T_10366_7 : _T_16690; // @[Mux.scala 46:16:@12446.4]
  assign _T_16693 = 6'h7 == _T_11317_57; // @[Mux.scala 46:19:@12447.4]
  assign _T_16694 = _T_16693 ? _T_10366_6 : _T_16692; // @[Mux.scala 46:16:@12448.4]
  assign _T_16695 = 6'h6 == _T_11317_57; // @[Mux.scala 46:19:@12449.4]
  assign _T_16696 = _T_16695 ? _T_10366_5 : _T_16694; // @[Mux.scala 46:16:@12450.4]
  assign _T_16697 = 6'h5 == _T_11317_57; // @[Mux.scala 46:19:@12451.4]
  assign _T_16698 = _T_16697 ? _T_10366_4 : _T_16696; // @[Mux.scala 46:16:@12452.4]
  assign _T_16699 = 6'h4 == _T_11317_57; // @[Mux.scala 46:19:@12453.4]
  assign _T_16700 = _T_16699 ? _T_10366_3 : _T_16698; // @[Mux.scala 46:16:@12454.4]
  assign _T_16701 = 6'h3 == _T_11317_57; // @[Mux.scala 46:19:@12455.4]
  assign _T_16702 = _T_16701 ? _T_10366_2 : _T_16700; // @[Mux.scala 46:16:@12456.4]
  assign _T_16703 = 6'h2 == _T_11317_57; // @[Mux.scala 46:19:@12457.4]
  assign _T_16704 = _T_16703 ? _T_10366_1 : _T_16702; // @[Mux.scala 46:16:@12458.4]
  assign _T_16705 = 6'h1 == _T_11317_57; // @[Mux.scala 46:19:@12459.4]
  assign _T_16706 = _T_16705 ? _T_10366_0 : _T_16704; // @[Mux.scala 46:16:@12460.4]
  assign _T_16767 = 6'h3b == _T_11317_58; // @[Mux.scala 46:19:@12462.4]
  assign _T_16768 = _T_16767 ? _T_10366_58 : 8'h0; // @[Mux.scala 46:16:@12463.4]
  assign _T_16769 = 6'h3a == _T_11317_58; // @[Mux.scala 46:19:@12464.4]
  assign _T_16770 = _T_16769 ? _T_10366_57 : _T_16768; // @[Mux.scala 46:16:@12465.4]
  assign _T_16771 = 6'h39 == _T_11317_58; // @[Mux.scala 46:19:@12466.4]
  assign _T_16772 = _T_16771 ? _T_10366_56 : _T_16770; // @[Mux.scala 46:16:@12467.4]
  assign _T_16773 = 6'h38 == _T_11317_58; // @[Mux.scala 46:19:@12468.4]
  assign _T_16774 = _T_16773 ? _T_10366_55 : _T_16772; // @[Mux.scala 46:16:@12469.4]
  assign _T_16775 = 6'h37 == _T_11317_58; // @[Mux.scala 46:19:@12470.4]
  assign _T_16776 = _T_16775 ? _T_10366_54 : _T_16774; // @[Mux.scala 46:16:@12471.4]
  assign _T_16777 = 6'h36 == _T_11317_58; // @[Mux.scala 46:19:@12472.4]
  assign _T_16778 = _T_16777 ? _T_10366_53 : _T_16776; // @[Mux.scala 46:16:@12473.4]
  assign _T_16779 = 6'h35 == _T_11317_58; // @[Mux.scala 46:19:@12474.4]
  assign _T_16780 = _T_16779 ? _T_10366_52 : _T_16778; // @[Mux.scala 46:16:@12475.4]
  assign _T_16781 = 6'h34 == _T_11317_58; // @[Mux.scala 46:19:@12476.4]
  assign _T_16782 = _T_16781 ? _T_10366_51 : _T_16780; // @[Mux.scala 46:16:@12477.4]
  assign _T_16783 = 6'h33 == _T_11317_58; // @[Mux.scala 46:19:@12478.4]
  assign _T_16784 = _T_16783 ? _T_10366_50 : _T_16782; // @[Mux.scala 46:16:@12479.4]
  assign _T_16785 = 6'h32 == _T_11317_58; // @[Mux.scala 46:19:@12480.4]
  assign _T_16786 = _T_16785 ? _T_10366_49 : _T_16784; // @[Mux.scala 46:16:@12481.4]
  assign _T_16787 = 6'h31 == _T_11317_58; // @[Mux.scala 46:19:@12482.4]
  assign _T_16788 = _T_16787 ? _T_10366_48 : _T_16786; // @[Mux.scala 46:16:@12483.4]
  assign _T_16789 = 6'h30 == _T_11317_58; // @[Mux.scala 46:19:@12484.4]
  assign _T_16790 = _T_16789 ? _T_10366_47 : _T_16788; // @[Mux.scala 46:16:@12485.4]
  assign _T_16791 = 6'h2f == _T_11317_58; // @[Mux.scala 46:19:@12486.4]
  assign _T_16792 = _T_16791 ? _T_10366_46 : _T_16790; // @[Mux.scala 46:16:@12487.4]
  assign _T_16793 = 6'h2e == _T_11317_58; // @[Mux.scala 46:19:@12488.4]
  assign _T_16794 = _T_16793 ? _T_10366_45 : _T_16792; // @[Mux.scala 46:16:@12489.4]
  assign _T_16795 = 6'h2d == _T_11317_58; // @[Mux.scala 46:19:@12490.4]
  assign _T_16796 = _T_16795 ? _T_10366_44 : _T_16794; // @[Mux.scala 46:16:@12491.4]
  assign _T_16797 = 6'h2c == _T_11317_58; // @[Mux.scala 46:19:@12492.4]
  assign _T_16798 = _T_16797 ? _T_10366_43 : _T_16796; // @[Mux.scala 46:16:@12493.4]
  assign _T_16799 = 6'h2b == _T_11317_58; // @[Mux.scala 46:19:@12494.4]
  assign _T_16800 = _T_16799 ? _T_10366_42 : _T_16798; // @[Mux.scala 46:16:@12495.4]
  assign _T_16801 = 6'h2a == _T_11317_58; // @[Mux.scala 46:19:@12496.4]
  assign _T_16802 = _T_16801 ? _T_10366_41 : _T_16800; // @[Mux.scala 46:16:@12497.4]
  assign _T_16803 = 6'h29 == _T_11317_58; // @[Mux.scala 46:19:@12498.4]
  assign _T_16804 = _T_16803 ? _T_10366_40 : _T_16802; // @[Mux.scala 46:16:@12499.4]
  assign _T_16805 = 6'h28 == _T_11317_58; // @[Mux.scala 46:19:@12500.4]
  assign _T_16806 = _T_16805 ? _T_10366_39 : _T_16804; // @[Mux.scala 46:16:@12501.4]
  assign _T_16807 = 6'h27 == _T_11317_58; // @[Mux.scala 46:19:@12502.4]
  assign _T_16808 = _T_16807 ? _T_10366_38 : _T_16806; // @[Mux.scala 46:16:@12503.4]
  assign _T_16809 = 6'h26 == _T_11317_58; // @[Mux.scala 46:19:@12504.4]
  assign _T_16810 = _T_16809 ? _T_10366_37 : _T_16808; // @[Mux.scala 46:16:@12505.4]
  assign _T_16811 = 6'h25 == _T_11317_58; // @[Mux.scala 46:19:@12506.4]
  assign _T_16812 = _T_16811 ? _T_10366_36 : _T_16810; // @[Mux.scala 46:16:@12507.4]
  assign _T_16813 = 6'h24 == _T_11317_58; // @[Mux.scala 46:19:@12508.4]
  assign _T_16814 = _T_16813 ? _T_10366_35 : _T_16812; // @[Mux.scala 46:16:@12509.4]
  assign _T_16815 = 6'h23 == _T_11317_58; // @[Mux.scala 46:19:@12510.4]
  assign _T_16816 = _T_16815 ? _T_10366_34 : _T_16814; // @[Mux.scala 46:16:@12511.4]
  assign _T_16817 = 6'h22 == _T_11317_58; // @[Mux.scala 46:19:@12512.4]
  assign _T_16818 = _T_16817 ? _T_10366_33 : _T_16816; // @[Mux.scala 46:16:@12513.4]
  assign _T_16819 = 6'h21 == _T_11317_58; // @[Mux.scala 46:19:@12514.4]
  assign _T_16820 = _T_16819 ? _T_10366_32 : _T_16818; // @[Mux.scala 46:16:@12515.4]
  assign _T_16821 = 6'h20 == _T_11317_58; // @[Mux.scala 46:19:@12516.4]
  assign _T_16822 = _T_16821 ? _T_10366_31 : _T_16820; // @[Mux.scala 46:16:@12517.4]
  assign _T_16823 = 6'h1f == _T_11317_58; // @[Mux.scala 46:19:@12518.4]
  assign _T_16824 = _T_16823 ? _T_10366_30 : _T_16822; // @[Mux.scala 46:16:@12519.4]
  assign _T_16825 = 6'h1e == _T_11317_58; // @[Mux.scala 46:19:@12520.4]
  assign _T_16826 = _T_16825 ? _T_10366_29 : _T_16824; // @[Mux.scala 46:16:@12521.4]
  assign _T_16827 = 6'h1d == _T_11317_58; // @[Mux.scala 46:19:@12522.4]
  assign _T_16828 = _T_16827 ? _T_10366_28 : _T_16826; // @[Mux.scala 46:16:@12523.4]
  assign _T_16829 = 6'h1c == _T_11317_58; // @[Mux.scala 46:19:@12524.4]
  assign _T_16830 = _T_16829 ? _T_10366_27 : _T_16828; // @[Mux.scala 46:16:@12525.4]
  assign _T_16831 = 6'h1b == _T_11317_58; // @[Mux.scala 46:19:@12526.4]
  assign _T_16832 = _T_16831 ? _T_10366_26 : _T_16830; // @[Mux.scala 46:16:@12527.4]
  assign _T_16833 = 6'h1a == _T_11317_58; // @[Mux.scala 46:19:@12528.4]
  assign _T_16834 = _T_16833 ? _T_10366_25 : _T_16832; // @[Mux.scala 46:16:@12529.4]
  assign _T_16835 = 6'h19 == _T_11317_58; // @[Mux.scala 46:19:@12530.4]
  assign _T_16836 = _T_16835 ? _T_10366_24 : _T_16834; // @[Mux.scala 46:16:@12531.4]
  assign _T_16837 = 6'h18 == _T_11317_58; // @[Mux.scala 46:19:@12532.4]
  assign _T_16838 = _T_16837 ? _T_10366_23 : _T_16836; // @[Mux.scala 46:16:@12533.4]
  assign _T_16839 = 6'h17 == _T_11317_58; // @[Mux.scala 46:19:@12534.4]
  assign _T_16840 = _T_16839 ? _T_10366_22 : _T_16838; // @[Mux.scala 46:16:@12535.4]
  assign _T_16841 = 6'h16 == _T_11317_58; // @[Mux.scala 46:19:@12536.4]
  assign _T_16842 = _T_16841 ? _T_10366_21 : _T_16840; // @[Mux.scala 46:16:@12537.4]
  assign _T_16843 = 6'h15 == _T_11317_58; // @[Mux.scala 46:19:@12538.4]
  assign _T_16844 = _T_16843 ? _T_10366_20 : _T_16842; // @[Mux.scala 46:16:@12539.4]
  assign _T_16845 = 6'h14 == _T_11317_58; // @[Mux.scala 46:19:@12540.4]
  assign _T_16846 = _T_16845 ? _T_10366_19 : _T_16844; // @[Mux.scala 46:16:@12541.4]
  assign _T_16847 = 6'h13 == _T_11317_58; // @[Mux.scala 46:19:@12542.4]
  assign _T_16848 = _T_16847 ? _T_10366_18 : _T_16846; // @[Mux.scala 46:16:@12543.4]
  assign _T_16849 = 6'h12 == _T_11317_58; // @[Mux.scala 46:19:@12544.4]
  assign _T_16850 = _T_16849 ? _T_10366_17 : _T_16848; // @[Mux.scala 46:16:@12545.4]
  assign _T_16851 = 6'h11 == _T_11317_58; // @[Mux.scala 46:19:@12546.4]
  assign _T_16852 = _T_16851 ? _T_10366_16 : _T_16850; // @[Mux.scala 46:16:@12547.4]
  assign _T_16853 = 6'h10 == _T_11317_58; // @[Mux.scala 46:19:@12548.4]
  assign _T_16854 = _T_16853 ? _T_10366_15 : _T_16852; // @[Mux.scala 46:16:@12549.4]
  assign _T_16855 = 6'hf == _T_11317_58; // @[Mux.scala 46:19:@12550.4]
  assign _T_16856 = _T_16855 ? _T_10366_14 : _T_16854; // @[Mux.scala 46:16:@12551.4]
  assign _T_16857 = 6'he == _T_11317_58; // @[Mux.scala 46:19:@12552.4]
  assign _T_16858 = _T_16857 ? _T_10366_13 : _T_16856; // @[Mux.scala 46:16:@12553.4]
  assign _T_16859 = 6'hd == _T_11317_58; // @[Mux.scala 46:19:@12554.4]
  assign _T_16860 = _T_16859 ? _T_10366_12 : _T_16858; // @[Mux.scala 46:16:@12555.4]
  assign _T_16861 = 6'hc == _T_11317_58; // @[Mux.scala 46:19:@12556.4]
  assign _T_16862 = _T_16861 ? _T_10366_11 : _T_16860; // @[Mux.scala 46:16:@12557.4]
  assign _T_16863 = 6'hb == _T_11317_58; // @[Mux.scala 46:19:@12558.4]
  assign _T_16864 = _T_16863 ? _T_10366_10 : _T_16862; // @[Mux.scala 46:16:@12559.4]
  assign _T_16865 = 6'ha == _T_11317_58; // @[Mux.scala 46:19:@12560.4]
  assign _T_16866 = _T_16865 ? _T_10366_9 : _T_16864; // @[Mux.scala 46:16:@12561.4]
  assign _T_16867 = 6'h9 == _T_11317_58; // @[Mux.scala 46:19:@12562.4]
  assign _T_16868 = _T_16867 ? _T_10366_8 : _T_16866; // @[Mux.scala 46:16:@12563.4]
  assign _T_16869 = 6'h8 == _T_11317_58; // @[Mux.scala 46:19:@12564.4]
  assign _T_16870 = _T_16869 ? _T_10366_7 : _T_16868; // @[Mux.scala 46:16:@12565.4]
  assign _T_16871 = 6'h7 == _T_11317_58; // @[Mux.scala 46:19:@12566.4]
  assign _T_16872 = _T_16871 ? _T_10366_6 : _T_16870; // @[Mux.scala 46:16:@12567.4]
  assign _T_16873 = 6'h6 == _T_11317_58; // @[Mux.scala 46:19:@12568.4]
  assign _T_16874 = _T_16873 ? _T_10366_5 : _T_16872; // @[Mux.scala 46:16:@12569.4]
  assign _T_16875 = 6'h5 == _T_11317_58; // @[Mux.scala 46:19:@12570.4]
  assign _T_16876 = _T_16875 ? _T_10366_4 : _T_16874; // @[Mux.scala 46:16:@12571.4]
  assign _T_16877 = 6'h4 == _T_11317_58; // @[Mux.scala 46:19:@12572.4]
  assign _T_16878 = _T_16877 ? _T_10366_3 : _T_16876; // @[Mux.scala 46:16:@12573.4]
  assign _T_16879 = 6'h3 == _T_11317_58; // @[Mux.scala 46:19:@12574.4]
  assign _T_16880 = _T_16879 ? _T_10366_2 : _T_16878; // @[Mux.scala 46:16:@12575.4]
  assign _T_16881 = 6'h2 == _T_11317_58; // @[Mux.scala 46:19:@12576.4]
  assign _T_16882 = _T_16881 ? _T_10366_1 : _T_16880; // @[Mux.scala 46:16:@12577.4]
  assign _T_16883 = 6'h1 == _T_11317_58; // @[Mux.scala 46:19:@12578.4]
  assign _T_16884 = _T_16883 ? _T_10366_0 : _T_16882; // @[Mux.scala 46:16:@12579.4]
  assign _T_16946 = 6'h3c == _T_11317_59; // @[Mux.scala 46:19:@12581.4]
  assign _T_16947 = _T_16946 ? _T_10366_59 : 8'h0; // @[Mux.scala 46:16:@12582.4]
  assign _T_16948 = 6'h3b == _T_11317_59; // @[Mux.scala 46:19:@12583.4]
  assign _T_16949 = _T_16948 ? _T_10366_58 : _T_16947; // @[Mux.scala 46:16:@12584.4]
  assign _T_16950 = 6'h3a == _T_11317_59; // @[Mux.scala 46:19:@12585.4]
  assign _T_16951 = _T_16950 ? _T_10366_57 : _T_16949; // @[Mux.scala 46:16:@12586.4]
  assign _T_16952 = 6'h39 == _T_11317_59; // @[Mux.scala 46:19:@12587.4]
  assign _T_16953 = _T_16952 ? _T_10366_56 : _T_16951; // @[Mux.scala 46:16:@12588.4]
  assign _T_16954 = 6'h38 == _T_11317_59; // @[Mux.scala 46:19:@12589.4]
  assign _T_16955 = _T_16954 ? _T_10366_55 : _T_16953; // @[Mux.scala 46:16:@12590.4]
  assign _T_16956 = 6'h37 == _T_11317_59; // @[Mux.scala 46:19:@12591.4]
  assign _T_16957 = _T_16956 ? _T_10366_54 : _T_16955; // @[Mux.scala 46:16:@12592.4]
  assign _T_16958 = 6'h36 == _T_11317_59; // @[Mux.scala 46:19:@12593.4]
  assign _T_16959 = _T_16958 ? _T_10366_53 : _T_16957; // @[Mux.scala 46:16:@12594.4]
  assign _T_16960 = 6'h35 == _T_11317_59; // @[Mux.scala 46:19:@12595.4]
  assign _T_16961 = _T_16960 ? _T_10366_52 : _T_16959; // @[Mux.scala 46:16:@12596.4]
  assign _T_16962 = 6'h34 == _T_11317_59; // @[Mux.scala 46:19:@12597.4]
  assign _T_16963 = _T_16962 ? _T_10366_51 : _T_16961; // @[Mux.scala 46:16:@12598.4]
  assign _T_16964 = 6'h33 == _T_11317_59; // @[Mux.scala 46:19:@12599.4]
  assign _T_16965 = _T_16964 ? _T_10366_50 : _T_16963; // @[Mux.scala 46:16:@12600.4]
  assign _T_16966 = 6'h32 == _T_11317_59; // @[Mux.scala 46:19:@12601.4]
  assign _T_16967 = _T_16966 ? _T_10366_49 : _T_16965; // @[Mux.scala 46:16:@12602.4]
  assign _T_16968 = 6'h31 == _T_11317_59; // @[Mux.scala 46:19:@12603.4]
  assign _T_16969 = _T_16968 ? _T_10366_48 : _T_16967; // @[Mux.scala 46:16:@12604.4]
  assign _T_16970 = 6'h30 == _T_11317_59; // @[Mux.scala 46:19:@12605.4]
  assign _T_16971 = _T_16970 ? _T_10366_47 : _T_16969; // @[Mux.scala 46:16:@12606.4]
  assign _T_16972 = 6'h2f == _T_11317_59; // @[Mux.scala 46:19:@12607.4]
  assign _T_16973 = _T_16972 ? _T_10366_46 : _T_16971; // @[Mux.scala 46:16:@12608.4]
  assign _T_16974 = 6'h2e == _T_11317_59; // @[Mux.scala 46:19:@12609.4]
  assign _T_16975 = _T_16974 ? _T_10366_45 : _T_16973; // @[Mux.scala 46:16:@12610.4]
  assign _T_16976 = 6'h2d == _T_11317_59; // @[Mux.scala 46:19:@12611.4]
  assign _T_16977 = _T_16976 ? _T_10366_44 : _T_16975; // @[Mux.scala 46:16:@12612.4]
  assign _T_16978 = 6'h2c == _T_11317_59; // @[Mux.scala 46:19:@12613.4]
  assign _T_16979 = _T_16978 ? _T_10366_43 : _T_16977; // @[Mux.scala 46:16:@12614.4]
  assign _T_16980 = 6'h2b == _T_11317_59; // @[Mux.scala 46:19:@12615.4]
  assign _T_16981 = _T_16980 ? _T_10366_42 : _T_16979; // @[Mux.scala 46:16:@12616.4]
  assign _T_16982 = 6'h2a == _T_11317_59; // @[Mux.scala 46:19:@12617.4]
  assign _T_16983 = _T_16982 ? _T_10366_41 : _T_16981; // @[Mux.scala 46:16:@12618.4]
  assign _T_16984 = 6'h29 == _T_11317_59; // @[Mux.scala 46:19:@12619.4]
  assign _T_16985 = _T_16984 ? _T_10366_40 : _T_16983; // @[Mux.scala 46:16:@12620.4]
  assign _T_16986 = 6'h28 == _T_11317_59; // @[Mux.scala 46:19:@12621.4]
  assign _T_16987 = _T_16986 ? _T_10366_39 : _T_16985; // @[Mux.scala 46:16:@12622.4]
  assign _T_16988 = 6'h27 == _T_11317_59; // @[Mux.scala 46:19:@12623.4]
  assign _T_16989 = _T_16988 ? _T_10366_38 : _T_16987; // @[Mux.scala 46:16:@12624.4]
  assign _T_16990 = 6'h26 == _T_11317_59; // @[Mux.scala 46:19:@12625.4]
  assign _T_16991 = _T_16990 ? _T_10366_37 : _T_16989; // @[Mux.scala 46:16:@12626.4]
  assign _T_16992 = 6'h25 == _T_11317_59; // @[Mux.scala 46:19:@12627.4]
  assign _T_16993 = _T_16992 ? _T_10366_36 : _T_16991; // @[Mux.scala 46:16:@12628.4]
  assign _T_16994 = 6'h24 == _T_11317_59; // @[Mux.scala 46:19:@12629.4]
  assign _T_16995 = _T_16994 ? _T_10366_35 : _T_16993; // @[Mux.scala 46:16:@12630.4]
  assign _T_16996 = 6'h23 == _T_11317_59; // @[Mux.scala 46:19:@12631.4]
  assign _T_16997 = _T_16996 ? _T_10366_34 : _T_16995; // @[Mux.scala 46:16:@12632.4]
  assign _T_16998 = 6'h22 == _T_11317_59; // @[Mux.scala 46:19:@12633.4]
  assign _T_16999 = _T_16998 ? _T_10366_33 : _T_16997; // @[Mux.scala 46:16:@12634.4]
  assign _T_17000 = 6'h21 == _T_11317_59; // @[Mux.scala 46:19:@12635.4]
  assign _T_17001 = _T_17000 ? _T_10366_32 : _T_16999; // @[Mux.scala 46:16:@12636.4]
  assign _T_17002 = 6'h20 == _T_11317_59; // @[Mux.scala 46:19:@12637.4]
  assign _T_17003 = _T_17002 ? _T_10366_31 : _T_17001; // @[Mux.scala 46:16:@12638.4]
  assign _T_17004 = 6'h1f == _T_11317_59; // @[Mux.scala 46:19:@12639.4]
  assign _T_17005 = _T_17004 ? _T_10366_30 : _T_17003; // @[Mux.scala 46:16:@12640.4]
  assign _T_17006 = 6'h1e == _T_11317_59; // @[Mux.scala 46:19:@12641.4]
  assign _T_17007 = _T_17006 ? _T_10366_29 : _T_17005; // @[Mux.scala 46:16:@12642.4]
  assign _T_17008 = 6'h1d == _T_11317_59; // @[Mux.scala 46:19:@12643.4]
  assign _T_17009 = _T_17008 ? _T_10366_28 : _T_17007; // @[Mux.scala 46:16:@12644.4]
  assign _T_17010 = 6'h1c == _T_11317_59; // @[Mux.scala 46:19:@12645.4]
  assign _T_17011 = _T_17010 ? _T_10366_27 : _T_17009; // @[Mux.scala 46:16:@12646.4]
  assign _T_17012 = 6'h1b == _T_11317_59; // @[Mux.scala 46:19:@12647.4]
  assign _T_17013 = _T_17012 ? _T_10366_26 : _T_17011; // @[Mux.scala 46:16:@12648.4]
  assign _T_17014 = 6'h1a == _T_11317_59; // @[Mux.scala 46:19:@12649.4]
  assign _T_17015 = _T_17014 ? _T_10366_25 : _T_17013; // @[Mux.scala 46:16:@12650.4]
  assign _T_17016 = 6'h19 == _T_11317_59; // @[Mux.scala 46:19:@12651.4]
  assign _T_17017 = _T_17016 ? _T_10366_24 : _T_17015; // @[Mux.scala 46:16:@12652.4]
  assign _T_17018 = 6'h18 == _T_11317_59; // @[Mux.scala 46:19:@12653.4]
  assign _T_17019 = _T_17018 ? _T_10366_23 : _T_17017; // @[Mux.scala 46:16:@12654.4]
  assign _T_17020 = 6'h17 == _T_11317_59; // @[Mux.scala 46:19:@12655.4]
  assign _T_17021 = _T_17020 ? _T_10366_22 : _T_17019; // @[Mux.scala 46:16:@12656.4]
  assign _T_17022 = 6'h16 == _T_11317_59; // @[Mux.scala 46:19:@12657.4]
  assign _T_17023 = _T_17022 ? _T_10366_21 : _T_17021; // @[Mux.scala 46:16:@12658.4]
  assign _T_17024 = 6'h15 == _T_11317_59; // @[Mux.scala 46:19:@12659.4]
  assign _T_17025 = _T_17024 ? _T_10366_20 : _T_17023; // @[Mux.scala 46:16:@12660.4]
  assign _T_17026 = 6'h14 == _T_11317_59; // @[Mux.scala 46:19:@12661.4]
  assign _T_17027 = _T_17026 ? _T_10366_19 : _T_17025; // @[Mux.scala 46:16:@12662.4]
  assign _T_17028 = 6'h13 == _T_11317_59; // @[Mux.scala 46:19:@12663.4]
  assign _T_17029 = _T_17028 ? _T_10366_18 : _T_17027; // @[Mux.scala 46:16:@12664.4]
  assign _T_17030 = 6'h12 == _T_11317_59; // @[Mux.scala 46:19:@12665.4]
  assign _T_17031 = _T_17030 ? _T_10366_17 : _T_17029; // @[Mux.scala 46:16:@12666.4]
  assign _T_17032 = 6'h11 == _T_11317_59; // @[Mux.scala 46:19:@12667.4]
  assign _T_17033 = _T_17032 ? _T_10366_16 : _T_17031; // @[Mux.scala 46:16:@12668.4]
  assign _T_17034 = 6'h10 == _T_11317_59; // @[Mux.scala 46:19:@12669.4]
  assign _T_17035 = _T_17034 ? _T_10366_15 : _T_17033; // @[Mux.scala 46:16:@12670.4]
  assign _T_17036 = 6'hf == _T_11317_59; // @[Mux.scala 46:19:@12671.4]
  assign _T_17037 = _T_17036 ? _T_10366_14 : _T_17035; // @[Mux.scala 46:16:@12672.4]
  assign _T_17038 = 6'he == _T_11317_59; // @[Mux.scala 46:19:@12673.4]
  assign _T_17039 = _T_17038 ? _T_10366_13 : _T_17037; // @[Mux.scala 46:16:@12674.4]
  assign _T_17040 = 6'hd == _T_11317_59; // @[Mux.scala 46:19:@12675.4]
  assign _T_17041 = _T_17040 ? _T_10366_12 : _T_17039; // @[Mux.scala 46:16:@12676.4]
  assign _T_17042 = 6'hc == _T_11317_59; // @[Mux.scala 46:19:@12677.4]
  assign _T_17043 = _T_17042 ? _T_10366_11 : _T_17041; // @[Mux.scala 46:16:@12678.4]
  assign _T_17044 = 6'hb == _T_11317_59; // @[Mux.scala 46:19:@12679.4]
  assign _T_17045 = _T_17044 ? _T_10366_10 : _T_17043; // @[Mux.scala 46:16:@12680.4]
  assign _T_17046 = 6'ha == _T_11317_59; // @[Mux.scala 46:19:@12681.4]
  assign _T_17047 = _T_17046 ? _T_10366_9 : _T_17045; // @[Mux.scala 46:16:@12682.4]
  assign _T_17048 = 6'h9 == _T_11317_59; // @[Mux.scala 46:19:@12683.4]
  assign _T_17049 = _T_17048 ? _T_10366_8 : _T_17047; // @[Mux.scala 46:16:@12684.4]
  assign _T_17050 = 6'h8 == _T_11317_59; // @[Mux.scala 46:19:@12685.4]
  assign _T_17051 = _T_17050 ? _T_10366_7 : _T_17049; // @[Mux.scala 46:16:@12686.4]
  assign _T_17052 = 6'h7 == _T_11317_59; // @[Mux.scala 46:19:@12687.4]
  assign _T_17053 = _T_17052 ? _T_10366_6 : _T_17051; // @[Mux.scala 46:16:@12688.4]
  assign _T_17054 = 6'h6 == _T_11317_59; // @[Mux.scala 46:19:@12689.4]
  assign _T_17055 = _T_17054 ? _T_10366_5 : _T_17053; // @[Mux.scala 46:16:@12690.4]
  assign _T_17056 = 6'h5 == _T_11317_59; // @[Mux.scala 46:19:@12691.4]
  assign _T_17057 = _T_17056 ? _T_10366_4 : _T_17055; // @[Mux.scala 46:16:@12692.4]
  assign _T_17058 = 6'h4 == _T_11317_59; // @[Mux.scala 46:19:@12693.4]
  assign _T_17059 = _T_17058 ? _T_10366_3 : _T_17057; // @[Mux.scala 46:16:@12694.4]
  assign _T_17060 = 6'h3 == _T_11317_59; // @[Mux.scala 46:19:@12695.4]
  assign _T_17061 = _T_17060 ? _T_10366_2 : _T_17059; // @[Mux.scala 46:16:@12696.4]
  assign _T_17062 = 6'h2 == _T_11317_59; // @[Mux.scala 46:19:@12697.4]
  assign _T_17063 = _T_17062 ? _T_10366_1 : _T_17061; // @[Mux.scala 46:16:@12698.4]
  assign _T_17064 = 6'h1 == _T_11317_59; // @[Mux.scala 46:19:@12699.4]
  assign _T_17065 = _T_17064 ? _T_10366_0 : _T_17063; // @[Mux.scala 46:16:@12700.4]
  assign _T_17128 = 6'h3d == _T_11317_60; // @[Mux.scala 46:19:@12702.4]
  assign _T_17129 = _T_17128 ? _T_10366_60 : 8'h0; // @[Mux.scala 46:16:@12703.4]
  assign _T_17130 = 6'h3c == _T_11317_60; // @[Mux.scala 46:19:@12704.4]
  assign _T_17131 = _T_17130 ? _T_10366_59 : _T_17129; // @[Mux.scala 46:16:@12705.4]
  assign _T_17132 = 6'h3b == _T_11317_60; // @[Mux.scala 46:19:@12706.4]
  assign _T_17133 = _T_17132 ? _T_10366_58 : _T_17131; // @[Mux.scala 46:16:@12707.4]
  assign _T_17134 = 6'h3a == _T_11317_60; // @[Mux.scala 46:19:@12708.4]
  assign _T_17135 = _T_17134 ? _T_10366_57 : _T_17133; // @[Mux.scala 46:16:@12709.4]
  assign _T_17136 = 6'h39 == _T_11317_60; // @[Mux.scala 46:19:@12710.4]
  assign _T_17137 = _T_17136 ? _T_10366_56 : _T_17135; // @[Mux.scala 46:16:@12711.4]
  assign _T_17138 = 6'h38 == _T_11317_60; // @[Mux.scala 46:19:@12712.4]
  assign _T_17139 = _T_17138 ? _T_10366_55 : _T_17137; // @[Mux.scala 46:16:@12713.4]
  assign _T_17140 = 6'h37 == _T_11317_60; // @[Mux.scala 46:19:@12714.4]
  assign _T_17141 = _T_17140 ? _T_10366_54 : _T_17139; // @[Mux.scala 46:16:@12715.4]
  assign _T_17142 = 6'h36 == _T_11317_60; // @[Mux.scala 46:19:@12716.4]
  assign _T_17143 = _T_17142 ? _T_10366_53 : _T_17141; // @[Mux.scala 46:16:@12717.4]
  assign _T_17144 = 6'h35 == _T_11317_60; // @[Mux.scala 46:19:@12718.4]
  assign _T_17145 = _T_17144 ? _T_10366_52 : _T_17143; // @[Mux.scala 46:16:@12719.4]
  assign _T_17146 = 6'h34 == _T_11317_60; // @[Mux.scala 46:19:@12720.4]
  assign _T_17147 = _T_17146 ? _T_10366_51 : _T_17145; // @[Mux.scala 46:16:@12721.4]
  assign _T_17148 = 6'h33 == _T_11317_60; // @[Mux.scala 46:19:@12722.4]
  assign _T_17149 = _T_17148 ? _T_10366_50 : _T_17147; // @[Mux.scala 46:16:@12723.4]
  assign _T_17150 = 6'h32 == _T_11317_60; // @[Mux.scala 46:19:@12724.4]
  assign _T_17151 = _T_17150 ? _T_10366_49 : _T_17149; // @[Mux.scala 46:16:@12725.4]
  assign _T_17152 = 6'h31 == _T_11317_60; // @[Mux.scala 46:19:@12726.4]
  assign _T_17153 = _T_17152 ? _T_10366_48 : _T_17151; // @[Mux.scala 46:16:@12727.4]
  assign _T_17154 = 6'h30 == _T_11317_60; // @[Mux.scala 46:19:@12728.4]
  assign _T_17155 = _T_17154 ? _T_10366_47 : _T_17153; // @[Mux.scala 46:16:@12729.4]
  assign _T_17156 = 6'h2f == _T_11317_60; // @[Mux.scala 46:19:@12730.4]
  assign _T_17157 = _T_17156 ? _T_10366_46 : _T_17155; // @[Mux.scala 46:16:@12731.4]
  assign _T_17158 = 6'h2e == _T_11317_60; // @[Mux.scala 46:19:@12732.4]
  assign _T_17159 = _T_17158 ? _T_10366_45 : _T_17157; // @[Mux.scala 46:16:@12733.4]
  assign _T_17160 = 6'h2d == _T_11317_60; // @[Mux.scala 46:19:@12734.4]
  assign _T_17161 = _T_17160 ? _T_10366_44 : _T_17159; // @[Mux.scala 46:16:@12735.4]
  assign _T_17162 = 6'h2c == _T_11317_60; // @[Mux.scala 46:19:@12736.4]
  assign _T_17163 = _T_17162 ? _T_10366_43 : _T_17161; // @[Mux.scala 46:16:@12737.4]
  assign _T_17164 = 6'h2b == _T_11317_60; // @[Mux.scala 46:19:@12738.4]
  assign _T_17165 = _T_17164 ? _T_10366_42 : _T_17163; // @[Mux.scala 46:16:@12739.4]
  assign _T_17166 = 6'h2a == _T_11317_60; // @[Mux.scala 46:19:@12740.4]
  assign _T_17167 = _T_17166 ? _T_10366_41 : _T_17165; // @[Mux.scala 46:16:@12741.4]
  assign _T_17168 = 6'h29 == _T_11317_60; // @[Mux.scala 46:19:@12742.4]
  assign _T_17169 = _T_17168 ? _T_10366_40 : _T_17167; // @[Mux.scala 46:16:@12743.4]
  assign _T_17170 = 6'h28 == _T_11317_60; // @[Mux.scala 46:19:@12744.4]
  assign _T_17171 = _T_17170 ? _T_10366_39 : _T_17169; // @[Mux.scala 46:16:@12745.4]
  assign _T_17172 = 6'h27 == _T_11317_60; // @[Mux.scala 46:19:@12746.4]
  assign _T_17173 = _T_17172 ? _T_10366_38 : _T_17171; // @[Mux.scala 46:16:@12747.4]
  assign _T_17174 = 6'h26 == _T_11317_60; // @[Mux.scala 46:19:@12748.4]
  assign _T_17175 = _T_17174 ? _T_10366_37 : _T_17173; // @[Mux.scala 46:16:@12749.4]
  assign _T_17176 = 6'h25 == _T_11317_60; // @[Mux.scala 46:19:@12750.4]
  assign _T_17177 = _T_17176 ? _T_10366_36 : _T_17175; // @[Mux.scala 46:16:@12751.4]
  assign _T_17178 = 6'h24 == _T_11317_60; // @[Mux.scala 46:19:@12752.4]
  assign _T_17179 = _T_17178 ? _T_10366_35 : _T_17177; // @[Mux.scala 46:16:@12753.4]
  assign _T_17180 = 6'h23 == _T_11317_60; // @[Mux.scala 46:19:@12754.4]
  assign _T_17181 = _T_17180 ? _T_10366_34 : _T_17179; // @[Mux.scala 46:16:@12755.4]
  assign _T_17182 = 6'h22 == _T_11317_60; // @[Mux.scala 46:19:@12756.4]
  assign _T_17183 = _T_17182 ? _T_10366_33 : _T_17181; // @[Mux.scala 46:16:@12757.4]
  assign _T_17184 = 6'h21 == _T_11317_60; // @[Mux.scala 46:19:@12758.4]
  assign _T_17185 = _T_17184 ? _T_10366_32 : _T_17183; // @[Mux.scala 46:16:@12759.4]
  assign _T_17186 = 6'h20 == _T_11317_60; // @[Mux.scala 46:19:@12760.4]
  assign _T_17187 = _T_17186 ? _T_10366_31 : _T_17185; // @[Mux.scala 46:16:@12761.4]
  assign _T_17188 = 6'h1f == _T_11317_60; // @[Mux.scala 46:19:@12762.4]
  assign _T_17189 = _T_17188 ? _T_10366_30 : _T_17187; // @[Mux.scala 46:16:@12763.4]
  assign _T_17190 = 6'h1e == _T_11317_60; // @[Mux.scala 46:19:@12764.4]
  assign _T_17191 = _T_17190 ? _T_10366_29 : _T_17189; // @[Mux.scala 46:16:@12765.4]
  assign _T_17192 = 6'h1d == _T_11317_60; // @[Mux.scala 46:19:@12766.4]
  assign _T_17193 = _T_17192 ? _T_10366_28 : _T_17191; // @[Mux.scala 46:16:@12767.4]
  assign _T_17194 = 6'h1c == _T_11317_60; // @[Mux.scala 46:19:@12768.4]
  assign _T_17195 = _T_17194 ? _T_10366_27 : _T_17193; // @[Mux.scala 46:16:@12769.4]
  assign _T_17196 = 6'h1b == _T_11317_60; // @[Mux.scala 46:19:@12770.4]
  assign _T_17197 = _T_17196 ? _T_10366_26 : _T_17195; // @[Mux.scala 46:16:@12771.4]
  assign _T_17198 = 6'h1a == _T_11317_60; // @[Mux.scala 46:19:@12772.4]
  assign _T_17199 = _T_17198 ? _T_10366_25 : _T_17197; // @[Mux.scala 46:16:@12773.4]
  assign _T_17200 = 6'h19 == _T_11317_60; // @[Mux.scala 46:19:@12774.4]
  assign _T_17201 = _T_17200 ? _T_10366_24 : _T_17199; // @[Mux.scala 46:16:@12775.4]
  assign _T_17202 = 6'h18 == _T_11317_60; // @[Mux.scala 46:19:@12776.4]
  assign _T_17203 = _T_17202 ? _T_10366_23 : _T_17201; // @[Mux.scala 46:16:@12777.4]
  assign _T_17204 = 6'h17 == _T_11317_60; // @[Mux.scala 46:19:@12778.4]
  assign _T_17205 = _T_17204 ? _T_10366_22 : _T_17203; // @[Mux.scala 46:16:@12779.4]
  assign _T_17206 = 6'h16 == _T_11317_60; // @[Mux.scala 46:19:@12780.4]
  assign _T_17207 = _T_17206 ? _T_10366_21 : _T_17205; // @[Mux.scala 46:16:@12781.4]
  assign _T_17208 = 6'h15 == _T_11317_60; // @[Mux.scala 46:19:@12782.4]
  assign _T_17209 = _T_17208 ? _T_10366_20 : _T_17207; // @[Mux.scala 46:16:@12783.4]
  assign _T_17210 = 6'h14 == _T_11317_60; // @[Mux.scala 46:19:@12784.4]
  assign _T_17211 = _T_17210 ? _T_10366_19 : _T_17209; // @[Mux.scala 46:16:@12785.4]
  assign _T_17212 = 6'h13 == _T_11317_60; // @[Mux.scala 46:19:@12786.4]
  assign _T_17213 = _T_17212 ? _T_10366_18 : _T_17211; // @[Mux.scala 46:16:@12787.4]
  assign _T_17214 = 6'h12 == _T_11317_60; // @[Mux.scala 46:19:@12788.4]
  assign _T_17215 = _T_17214 ? _T_10366_17 : _T_17213; // @[Mux.scala 46:16:@12789.4]
  assign _T_17216 = 6'h11 == _T_11317_60; // @[Mux.scala 46:19:@12790.4]
  assign _T_17217 = _T_17216 ? _T_10366_16 : _T_17215; // @[Mux.scala 46:16:@12791.4]
  assign _T_17218 = 6'h10 == _T_11317_60; // @[Mux.scala 46:19:@12792.4]
  assign _T_17219 = _T_17218 ? _T_10366_15 : _T_17217; // @[Mux.scala 46:16:@12793.4]
  assign _T_17220 = 6'hf == _T_11317_60; // @[Mux.scala 46:19:@12794.4]
  assign _T_17221 = _T_17220 ? _T_10366_14 : _T_17219; // @[Mux.scala 46:16:@12795.4]
  assign _T_17222 = 6'he == _T_11317_60; // @[Mux.scala 46:19:@12796.4]
  assign _T_17223 = _T_17222 ? _T_10366_13 : _T_17221; // @[Mux.scala 46:16:@12797.4]
  assign _T_17224 = 6'hd == _T_11317_60; // @[Mux.scala 46:19:@12798.4]
  assign _T_17225 = _T_17224 ? _T_10366_12 : _T_17223; // @[Mux.scala 46:16:@12799.4]
  assign _T_17226 = 6'hc == _T_11317_60; // @[Mux.scala 46:19:@12800.4]
  assign _T_17227 = _T_17226 ? _T_10366_11 : _T_17225; // @[Mux.scala 46:16:@12801.4]
  assign _T_17228 = 6'hb == _T_11317_60; // @[Mux.scala 46:19:@12802.4]
  assign _T_17229 = _T_17228 ? _T_10366_10 : _T_17227; // @[Mux.scala 46:16:@12803.4]
  assign _T_17230 = 6'ha == _T_11317_60; // @[Mux.scala 46:19:@12804.4]
  assign _T_17231 = _T_17230 ? _T_10366_9 : _T_17229; // @[Mux.scala 46:16:@12805.4]
  assign _T_17232 = 6'h9 == _T_11317_60; // @[Mux.scala 46:19:@12806.4]
  assign _T_17233 = _T_17232 ? _T_10366_8 : _T_17231; // @[Mux.scala 46:16:@12807.4]
  assign _T_17234 = 6'h8 == _T_11317_60; // @[Mux.scala 46:19:@12808.4]
  assign _T_17235 = _T_17234 ? _T_10366_7 : _T_17233; // @[Mux.scala 46:16:@12809.4]
  assign _T_17236 = 6'h7 == _T_11317_60; // @[Mux.scala 46:19:@12810.4]
  assign _T_17237 = _T_17236 ? _T_10366_6 : _T_17235; // @[Mux.scala 46:16:@12811.4]
  assign _T_17238 = 6'h6 == _T_11317_60; // @[Mux.scala 46:19:@12812.4]
  assign _T_17239 = _T_17238 ? _T_10366_5 : _T_17237; // @[Mux.scala 46:16:@12813.4]
  assign _T_17240 = 6'h5 == _T_11317_60; // @[Mux.scala 46:19:@12814.4]
  assign _T_17241 = _T_17240 ? _T_10366_4 : _T_17239; // @[Mux.scala 46:16:@12815.4]
  assign _T_17242 = 6'h4 == _T_11317_60; // @[Mux.scala 46:19:@12816.4]
  assign _T_17243 = _T_17242 ? _T_10366_3 : _T_17241; // @[Mux.scala 46:16:@12817.4]
  assign _T_17244 = 6'h3 == _T_11317_60; // @[Mux.scala 46:19:@12818.4]
  assign _T_17245 = _T_17244 ? _T_10366_2 : _T_17243; // @[Mux.scala 46:16:@12819.4]
  assign _T_17246 = 6'h2 == _T_11317_60; // @[Mux.scala 46:19:@12820.4]
  assign _T_17247 = _T_17246 ? _T_10366_1 : _T_17245; // @[Mux.scala 46:16:@12821.4]
  assign _T_17248 = 6'h1 == _T_11317_60; // @[Mux.scala 46:19:@12822.4]
  assign _T_17249 = _T_17248 ? _T_10366_0 : _T_17247; // @[Mux.scala 46:16:@12823.4]
  assign _T_17313 = 6'h3e == _T_11317_61; // @[Mux.scala 46:19:@12825.4]
  assign _T_17314 = _T_17313 ? _T_10366_61 : 8'h0; // @[Mux.scala 46:16:@12826.4]
  assign _T_17315 = 6'h3d == _T_11317_61; // @[Mux.scala 46:19:@12827.4]
  assign _T_17316 = _T_17315 ? _T_10366_60 : _T_17314; // @[Mux.scala 46:16:@12828.4]
  assign _T_17317 = 6'h3c == _T_11317_61; // @[Mux.scala 46:19:@12829.4]
  assign _T_17318 = _T_17317 ? _T_10366_59 : _T_17316; // @[Mux.scala 46:16:@12830.4]
  assign _T_17319 = 6'h3b == _T_11317_61; // @[Mux.scala 46:19:@12831.4]
  assign _T_17320 = _T_17319 ? _T_10366_58 : _T_17318; // @[Mux.scala 46:16:@12832.4]
  assign _T_17321 = 6'h3a == _T_11317_61; // @[Mux.scala 46:19:@12833.4]
  assign _T_17322 = _T_17321 ? _T_10366_57 : _T_17320; // @[Mux.scala 46:16:@12834.4]
  assign _T_17323 = 6'h39 == _T_11317_61; // @[Mux.scala 46:19:@12835.4]
  assign _T_17324 = _T_17323 ? _T_10366_56 : _T_17322; // @[Mux.scala 46:16:@12836.4]
  assign _T_17325 = 6'h38 == _T_11317_61; // @[Mux.scala 46:19:@12837.4]
  assign _T_17326 = _T_17325 ? _T_10366_55 : _T_17324; // @[Mux.scala 46:16:@12838.4]
  assign _T_17327 = 6'h37 == _T_11317_61; // @[Mux.scala 46:19:@12839.4]
  assign _T_17328 = _T_17327 ? _T_10366_54 : _T_17326; // @[Mux.scala 46:16:@12840.4]
  assign _T_17329 = 6'h36 == _T_11317_61; // @[Mux.scala 46:19:@12841.4]
  assign _T_17330 = _T_17329 ? _T_10366_53 : _T_17328; // @[Mux.scala 46:16:@12842.4]
  assign _T_17331 = 6'h35 == _T_11317_61; // @[Mux.scala 46:19:@12843.4]
  assign _T_17332 = _T_17331 ? _T_10366_52 : _T_17330; // @[Mux.scala 46:16:@12844.4]
  assign _T_17333 = 6'h34 == _T_11317_61; // @[Mux.scala 46:19:@12845.4]
  assign _T_17334 = _T_17333 ? _T_10366_51 : _T_17332; // @[Mux.scala 46:16:@12846.4]
  assign _T_17335 = 6'h33 == _T_11317_61; // @[Mux.scala 46:19:@12847.4]
  assign _T_17336 = _T_17335 ? _T_10366_50 : _T_17334; // @[Mux.scala 46:16:@12848.4]
  assign _T_17337 = 6'h32 == _T_11317_61; // @[Mux.scala 46:19:@12849.4]
  assign _T_17338 = _T_17337 ? _T_10366_49 : _T_17336; // @[Mux.scala 46:16:@12850.4]
  assign _T_17339 = 6'h31 == _T_11317_61; // @[Mux.scala 46:19:@12851.4]
  assign _T_17340 = _T_17339 ? _T_10366_48 : _T_17338; // @[Mux.scala 46:16:@12852.4]
  assign _T_17341 = 6'h30 == _T_11317_61; // @[Mux.scala 46:19:@12853.4]
  assign _T_17342 = _T_17341 ? _T_10366_47 : _T_17340; // @[Mux.scala 46:16:@12854.4]
  assign _T_17343 = 6'h2f == _T_11317_61; // @[Mux.scala 46:19:@12855.4]
  assign _T_17344 = _T_17343 ? _T_10366_46 : _T_17342; // @[Mux.scala 46:16:@12856.4]
  assign _T_17345 = 6'h2e == _T_11317_61; // @[Mux.scala 46:19:@12857.4]
  assign _T_17346 = _T_17345 ? _T_10366_45 : _T_17344; // @[Mux.scala 46:16:@12858.4]
  assign _T_17347 = 6'h2d == _T_11317_61; // @[Mux.scala 46:19:@12859.4]
  assign _T_17348 = _T_17347 ? _T_10366_44 : _T_17346; // @[Mux.scala 46:16:@12860.4]
  assign _T_17349 = 6'h2c == _T_11317_61; // @[Mux.scala 46:19:@12861.4]
  assign _T_17350 = _T_17349 ? _T_10366_43 : _T_17348; // @[Mux.scala 46:16:@12862.4]
  assign _T_17351 = 6'h2b == _T_11317_61; // @[Mux.scala 46:19:@12863.4]
  assign _T_17352 = _T_17351 ? _T_10366_42 : _T_17350; // @[Mux.scala 46:16:@12864.4]
  assign _T_17353 = 6'h2a == _T_11317_61; // @[Mux.scala 46:19:@12865.4]
  assign _T_17354 = _T_17353 ? _T_10366_41 : _T_17352; // @[Mux.scala 46:16:@12866.4]
  assign _T_17355 = 6'h29 == _T_11317_61; // @[Mux.scala 46:19:@12867.4]
  assign _T_17356 = _T_17355 ? _T_10366_40 : _T_17354; // @[Mux.scala 46:16:@12868.4]
  assign _T_17357 = 6'h28 == _T_11317_61; // @[Mux.scala 46:19:@12869.4]
  assign _T_17358 = _T_17357 ? _T_10366_39 : _T_17356; // @[Mux.scala 46:16:@12870.4]
  assign _T_17359 = 6'h27 == _T_11317_61; // @[Mux.scala 46:19:@12871.4]
  assign _T_17360 = _T_17359 ? _T_10366_38 : _T_17358; // @[Mux.scala 46:16:@12872.4]
  assign _T_17361 = 6'h26 == _T_11317_61; // @[Mux.scala 46:19:@12873.4]
  assign _T_17362 = _T_17361 ? _T_10366_37 : _T_17360; // @[Mux.scala 46:16:@12874.4]
  assign _T_17363 = 6'h25 == _T_11317_61; // @[Mux.scala 46:19:@12875.4]
  assign _T_17364 = _T_17363 ? _T_10366_36 : _T_17362; // @[Mux.scala 46:16:@12876.4]
  assign _T_17365 = 6'h24 == _T_11317_61; // @[Mux.scala 46:19:@12877.4]
  assign _T_17366 = _T_17365 ? _T_10366_35 : _T_17364; // @[Mux.scala 46:16:@12878.4]
  assign _T_17367 = 6'h23 == _T_11317_61; // @[Mux.scala 46:19:@12879.4]
  assign _T_17368 = _T_17367 ? _T_10366_34 : _T_17366; // @[Mux.scala 46:16:@12880.4]
  assign _T_17369 = 6'h22 == _T_11317_61; // @[Mux.scala 46:19:@12881.4]
  assign _T_17370 = _T_17369 ? _T_10366_33 : _T_17368; // @[Mux.scala 46:16:@12882.4]
  assign _T_17371 = 6'h21 == _T_11317_61; // @[Mux.scala 46:19:@12883.4]
  assign _T_17372 = _T_17371 ? _T_10366_32 : _T_17370; // @[Mux.scala 46:16:@12884.4]
  assign _T_17373 = 6'h20 == _T_11317_61; // @[Mux.scala 46:19:@12885.4]
  assign _T_17374 = _T_17373 ? _T_10366_31 : _T_17372; // @[Mux.scala 46:16:@12886.4]
  assign _T_17375 = 6'h1f == _T_11317_61; // @[Mux.scala 46:19:@12887.4]
  assign _T_17376 = _T_17375 ? _T_10366_30 : _T_17374; // @[Mux.scala 46:16:@12888.4]
  assign _T_17377 = 6'h1e == _T_11317_61; // @[Mux.scala 46:19:@12889.4]
  assign _T_17378 = _T_17377 ? _T_10366_29 : _T_17376; // @[Mux.scala 46:16:@12890.4]
  assign _T_17379 = 6'h1d == _T_11317_61; // @[Mux.scala 46:19:@12891.4]
  assign _T_17380 = _T_17379 ? _T_10366_28 : _T_17378; // @[Mux.scala 46:16:@12892.4]
  assign _T_17381 = 6'h1c == _T_11317_61; // @[Mux.scala 46:19:@12893.4]
  assign _T_17382 = _T_17381 ? _T_10366_27 : _T_17380; // @[Mux.scala 46:16:@12894.4]
  assign _T_17383 = 6'h1b == _T_11317_61; // @[Mux.scala 46:19:@12895.4]
  assign _T_17384 = _T_17383 ? _T_10366_26 : _T_17382; // @[Mux.scala 46:16:@12896.4]
  assign _T_17385 = 6'h1a == _T_11317_61; // @[Mux.scala 46:19:@12897.4]
  assign _T_17386 = _T_17385 ? _T_10366_25 : _T_17384; // @[Mux.scala 46:16:@12898.4]
  assign _T_17387 = 6'h19 == _T_11317_61; // @[Mux.scala 46:19:@12899.4]
  assign _T_17388 = _T_17387 ? _T_10366_24 : _T_17386; // @[Mux.scala 46:16:@12900.4]
  assign _T_17389 = 6'h18 == _T_11317_61; // @[Mux.scala 46:19:@12901.4]
  assign _T_17390 = _T_17389 ? _T_10366_23 : _T_17388; // @[Mux.scala 46:16:@12902.4]
  assign _T_17391 = 6'h17 == _T_11317_61; // @[Mux.scala 46:19:@12903.4]
  assign _T_17392 = _T_17391 ? _T_10366_22 : _T_17390; // @[Mux.scala 46:16:@12904.4]
  assign _T_17393 = 6'h16 == _T_11317_61; // @[Mux.scala 46:19:@12905.4]
  assign _T_17394 = _T_17393 ? _T_10366_21 : _T_17392; // @[Mux.scala 46:16:@12906.4]
  assign _T_17395 = 6'h15 == _T_11317_61; // @[Mux.scala 46:19:@12907.4]
  assign _T_17396 = _T_17395 ? _T_10366_20 : _T_17394; // @[Mux.scala 46:16:@12908.4]
  assign _T_17397 = 6'h14 == _T_11317_61; // @[Mux.scala 46:19:@12909.4]
  assign _T_17398 = _T_17397 ? _T_10366_19 : _T_17396; // @[Mux.scala 46:16:@12910.4]
  assign _T_17399 = 6'h13 == _T_11317_61; // @[Mux.scala 46:19:@12911.4]
  assign _T_17400 = _T_17399 ? _T_10366_18 : _T_17398; // @[Mux.scala 46:16:@12912.4]
  assign _T_17401 = 6'h12 == _T_11317_61; // @[Mux.scala 46:19:@12913.4]
  assign _T_17402 = _T_17401 ? _T_10366_17 : _T_17400; // @[Mux.scala 46:16:@12914.4]
  assign _T_17403 = 6'h11 == _T_11317_61; // @[Mux.scala 46:19:@12915.4]
  assign _T_17404 = _T_17403 ? _T_10366_16 : _T_17402; // @[Mux.scala 46:16:@12916.4]
  assign _T_17405 = 6'h10 == _T_11317_61; // @[Mux.scala 46:19:@12917.4]
  assign _T_17406 = _T_17405 ? _T_10366_15 : _T_17404; // @[Mux.scala 46:16:@12918.4]
  assign _T_17407 = 6'hf == _T_11317_61; // @[Mux.scala 46:19:@12919.4]
  assign _T_17408 = _T_17407 ? _T_10366_14 : _T_17406; // @[Mux.scala 46:16:@12920.4]
  assign _T_17409 = 6'he == _T_11317_61; // @[Mux.scala 46:19:@12921.4]
  assign _T_17410 = _T_17409 ? _T_10366_13 : _T_17408; // @[Mux.scala 46:16:@12922.4]
  assign _T_17411 = 6'hd == _T_11317_61; // @[Mux.scala 46:19:@12923.4]
  assign _T_17412 = _T_17411 ? _T_10366_12 : _T_17410; // @[Mux.scala 46:16:@12924.4]
  assign _T_17413 = 6'hc == _T_11317_61; // @[Mux.scala 46:19:@12925.4]
  assign _T_17414 = _T_17413 ? _T_10366_11 : _T_17412; // @[Mux.scala 46:16:@12926.4]
  assign _T_17415 = 6'hb == _T_11317_61; // @[Mux.scala 46:19:@12927.4]
  assign _T_17416 = _T_17415 ? _T_10366_10 : _T_17414; // @[Mux.scala 46:16:@12928.4]
  assign _T_17417 = 6'ha == _T_11317_61; // @[Mux.scala 46:19:@12929.4]
  assign _T_17418 = _T_17417 ? _T_10366_9 : _T_17416; // @[Mux.scala 46:16:@12930.4]
  assign _T_17419 = 6'h9 == _T_11317_61; // @[Mux.scala 46:19:@12931.4]
  assign _T_17420 = _T_17419 ? _T_10366_8 : _T_17418; // @[Mux.scala 46:16:@12932.4]
  assign _T_17421 = 6'h8 == _T_11317_61; // @[Mux.scala 46:19:@12933.4]
  assign _T_17422 = _T_17421 ? _T_10366_7 : _T_17420; // @[Mux.scala 46:16:@12934.4]
  assign _T_17423 = 6'h7 == _T_11317_61; // @[Mux.scala 46:19:@12935.4]
  assign _T_17424 = _T_17423 ? _T_10366_6 : _T_17422; // @[Mux.scala 46:16:@12936.4]
  assign _T_17425 = 6'h6 == _T_11317_61; // @[Mux.scala 46:19:@12937.4]
  assign _T_17426 = _T_17425 ? _T_10366_5 : _T_17424; // @[Mux.scala 46:16:@12938.4]
  assign _T_17427 = 6'h5 == _T_11317_61; // @[Mux.scala 46:19:@12939.4]
  assign _T_17428 = _T_17427 ? _T_10366_4 : _T_17426; // @[Mux.scala 46:16:@12940.4]
  assign _T_17429 = 6'h4 == _T_11317_61; // @[Mux.scala 46:19:@12941.4]
  assign _T_17430 = _T_17429 ? _T_10366_3 : _T_17428; // @[Mux.scala 46:16:@12942.4]
  assign _T_17431 = 6'h3 == _T_11317_61; // @[Mux.scala 46:19:@12943.4]
  assign _T_17432 = _T_17431 ? _T_10366_2 : _T_17430; // @[Mux.scala 46:16:@12944.4]
  assign _T_17433 = 6'h2 == _T_11317_61; // @[Mux.scala 46:19:@12945.4]
  assign _T_17434 = _T_17433 ? _T_10366_1 : _T_17432; // @[Mux.scala 46:16:@12946.4]
  assign _T_17435 = 6'h1 == _T_11317_61; // @[Mux.scala 46:19:@12947.4]
  assign _T_17436 = _T_17435 ? _T_10366_0 : _T_17434; // @[Mux.scala 46:16:@12948.4]
  assign _T_17501 = 6'h3f == _T_11317_62; // @[Mux.scala 46:19:@12950.4]
  assign _T_17502 = _T_17501 ? _T_10366_62 : 8'h0; // @[Mux.scala 46:16:@12951.4]
  assign _T_17503 = 6'h3e == _T_11317_62; // @[Mux.scala 46:19:@12952.4]
  assign _T_17504 = _T_17503 ? _T_10366_61 : _T_17502; // @[Mux.scala 46:16:@12953.4]
  assign _T_17505 = 6'h3d == _T_11317_62; // @[Mux.scala 46:19:@12954.4]
  assign _T_17506 = _T_17505 ? _T_10366_60 : _T_17504; // @[Mux.scala 46:16:@12955.4]
  assign _T_17507 = 6'h3c == _T_11317_62; // @[Mux.scala 46:19:@12956.4]
  assign _T_17508 = _T_17507 ? _T_10366_59 : _T_17506; // @[Mux.scala 46:16:@12957.4]
  assign _T_17509 = 6'h3b == _T_11317_62; // @[Mux.scala 46:19:@12958.4]
  assign _T_17510 = _T_17509 ? _T_10366_58 : _T_17508; // @[Mux.scala 46:16:@12959.4]
  assign _T_17511 = 6'h3a == _T_11317_62; // @[Mux.scala 46:19:@12960.4]
  assign _T_17512 = _T_17511 ? _T_10366_57 : _T_17510; // @[Mux.scala 46:16:@12961.4]
  assign _T_17513 = 6'h39 == _T_11317_62; // @[Mux.scala 46:19:@12962.4]
  assign _T_17514 = _T_17513 ? _T_10366_56 : _T_17512; // @[Mux.scala 46:16:@12963.4]
  assign _T_17515 = 6'h38 == _T_11317_62; // @[Mux.scala 46:19:@12964.4]
  assign _T_17516 = _T_17515 ? _T_10366_55 : _T_17514; // @[Mux.scala 46:16:@12965.4]
  assign _T_17517 = 6'h37 == _T_11317_62; // @[Mux.scala 46:19:@12966.4]
  assign _T_17518 = _T_17517 ? _T_10366_54 : _T_17516; // @[Mux.scala 46:16:@12967.4]
  assign _T_17519 = 6'h36 == _T_11317_62; // @[Mux.scala 46:19:@12968.4]
  assign _T_17520 = _T_17519 ? _T_10366_53 : _T_17518; // @[Mux.scala 46:16:@12969.4]
  assign _T_17521 = 6'h35 == _T_11317_62; // @[Mux.scala 46:19:@12970.4]
  assign _T_17522 = _T_17521 ? _T_10366_52 : _T_17520; // @[Mux.scala 46:16:@12971.4]
  assign _T_17523 = 6'h34 == _T_11317_62; // @[Mux.scala 46:19:@12972.4]
  assign _T_17524 = _T_17523 ? _T_10366_51 : _T_17522; // @[Mux.scala 46:16:@12973.4]
  assign _T_17525 = 6'h33 == _T_11317_62; // @[Mux.scala 46:19:@12974.4]
  assign _T_17526 = _T_17525 ? _T_10366_50 : _T_17524; // @[Mux.scala 46:16:@12975.4]
  assign _T_17527 = 6'h32 == _T_11317_62; // @[Mux.scala 46:19:@12976.4]
  assign _T_17528 = _T_17527 ? _T_10366_49 : _T_17526; // @[Mux.scala 46:16:@12977.4]
  assign _T_17529 = 6'h31 == _T_11317_62; // @[Mux.scala 46:19:@12978.4]
  assign _T_17530 = _T_17529 ? _T_10366_48 : _T_17528; // @[Mux.scala 46:16:@12979.4]
  assign _T_17531 = 6'h30 == _T_11317_62; // @[Mux.scala 46:19:@12980.4]
  assign _T_17532 = _T_17531 ? _T_10366_47 : _T_17530; // @[Mux.scala 46:16:@12981.4]
  assign _T_17533 = 6'h2f == _T_11317_62; // @[Mux.scala 46:19:@12982.4]
  assign _T_17534 = _T_17533 ? _T_10366_46 : _T_17532; // @[Mux.scala 46:16:@12983.4]
  assign _T_17535 = 6'h2e == _T_11317_62; // @[Mux.scala 46:19:@12984.4]
  assign _T_17536 = _T_17535 ? _T_10366_45 : _T_17534; // @[Mux.scala 46:16:@12985.4]
  assign _T_17537 = 6'h2d == _T_11317_62; // @[Mux.scala 46:19:@12986.4]
  assign _T_17538 = _T_17537 ? _T_10366_44 : _T_17536; // @[Mux.scala 46:16:@12987.4]
  assign _T_17539 = 6'h2c == _T_11317_62; // @[Mux.scala 46:19:@12988.4]
  assign _T_17540 = _T_17539 ? _T_10366_43 : _T_17538; // @[Mux.scala 46:16:@12989.4]
  assign _T_17541 = 6'h2b == _T_11317_62; // @[Mux.scala 46:19:@12990.4]
  assign _T_17542 = _T_17541 ? _T_10366_42 : _T_17540; // @[Mux.scala 46:16:@12991.4]
  assign _T_17543 = 6'h2a == _T_11317_62; // @[Mux.scala 46:19:@12992.4]
  assign _T_17544 = _T_17543 ? _T_10366_41 : _T_17542; // @[Mux.scala 46:16:@12993.4]
  assign _T_17545 = 6'h29 == _T_11317_62; // @[Mux.scala 46:19:@12994.4]
  assign _T_17546 = _T_17545 ? _T_10366_40 : _T_17544; // @[Mux.scala 46:16:@12995.4]
  assign _T_17547 = 6'h28 == _T_11317_62; // @[Mux.scala 46:19:@12996.4]
  assign _T_17548 = _T_17547 ? _T_10366_39 : _T_17546; // @[Mux.scala 46:16:@12997.4]
  assign _T_17549 = 6'h27 == _T_11317_62; // @[Mux.scala 46:19:@12998.4]
  assign _T_17550 = _T_17549 ? _T_10366_38 : _T_17548; // @[Mux.scala 46:16:@12999.4]
  assign _T_17551 = 6'h26 == _T_11317_62; // @[Mux.scala 46:19:@13000.4]
  assign _T_17552 = _T_17551 ? _T_10366_37 : _T_17550; // @[Mux.scala 46:16:@13001.4]
  assign _T_17553 = 6'h25 == _T_11317_62; // @[Mux.scala 46:19:@13002.4]
  assign _T_17554 = _T_17553 ? _T_10366_36 : _T_17552; // @[Mux.scala 46:16:@13003.4]
  assign _T_17555 = 6'h24 == _T_11317_62; // @[Mux.scala 46:19:@13004.4]
  assign _T_17556 = _T_17555 ? _T_10366_35 : _T_17554; // @[Mux.scala 46:16:@13005.4]
  assign _T_17557 = 6'h23 == _T_11317_62; // @[Mux.scala 46:19:@13006.4]
  assign _T_17558 = _T_17557 ? _T_10366_34 : _T_17556; // @[Mux.scala 46:16:@13007.4]
  assign _T_17559 = 6'h22 == _T_11317_62; // @[Mux.scala 46:19:@13008.4]
  assign _T_17560 = _T_17559 ? _T_10366_33 : _T_17558; // @[Mux.scala 46:16:@13009.4]
  assign _T_17561 = 6'h21 == _T_11317_62; // @[Mux.scala 46:19:@13010.4]
  assign _T_17562 = _T_17561 ? _T_10366_32 : _T_17560; // @[Mux.scala 46:16:@13011.4]
  assign _T_17563 = 6'h20 == _T_11317_62; // @[Mux.scala 46:19:@13012.4]
  assign _T_17564 = _T_17563 ? _T_10366_31 : _T_17562; // @[Mux.scala 46:16:@13013.4]
  assign _T_17565 = 6'h1f == _T_11317_62; // @[Mux.scala 46:19:@13014.4]
  assign _T_17566 = _T_17565 ? _T_10366_30 : _T_17564; // @[Mux.scala 46:16:@13015.4]
  assign _T_17567 = 6'h1e == _T_11317_62; // @[Mux.scala 46:19:@13016.4]
  assign _T_17568 = _T_17567 ? _T_10366_29 : _T_17566; // @[Mux.scala 46:16:@13017.4]
  assign _T_17569 = 6'h1d == _T_11317_62; // @[Mux.scala 46:19:@13018.4]
  assign _T_17570 = _T_17569 ? _T_10366_28 : _T_17568; // @[Mux.scala 46:16:@13019.4]
  assign _T_17571 = 6'h1c == _T_11317_62; // @[Mux.scala 46:19:@13020.4]
  assign _T_17572 = _T_17571 ? _T_10366_27 : _T_17570; // @[Mux.scala 46:16:@13021.4]
  assign _T_17573 = 6'h1b == _T_11317_62; // @[Mux.scala 46:19:@13022.4]
  assign _T_17574 = _T_17573 ? _T_10366_26 : _T_17572; // @[Mux.scala 46:16:@13023.4]
  assign _T_17575 = 6'h1a == _T_11317_62; // @[Mux.scala 46:19:@13024.4]
  assign _T_17576 = _T_17575 ? _T_10366_25 : _T_17574; // @[Mux.scala 46:16:@13025.4]
  assign _T_17577 = 6'h19 == _T_11317_62; // @[Mux.scala 46:19:@13026.4]
  assign _T_17578 = _T_17577 ? _T_10366_24 : _T_17576; // @[Mux.scala 46:16:@13027.4]
  assign _T_17579 = 6'h18 == _T_11317_62; // @[Mux.scala 46:19:@13028.4]
  assign _T_17580 = _T_17579 ? _T_10366_23 : _T_17578; // @[Mux.scala 46:16:@13029.4]
  assign _T_17581 = 6'h17 == _T_11317_62; // @[Mux.scala 46:19:@13030.4]
  assign _T_17582 = _T_17581 ? _T_10366_22 : _T_17580; // @[Mux.scala 46:16:@13031.4]
  assign _T_17583 = 6'h16 == _T_11317_62; // @[Mux.scala 46:19:@13032.4]
  assign _T_17584 = _T_17583 ? _T_10366_21 : _T_17582; // @[Mux.scala 46:16:@13033.4]
  assign _T_17585 = 6'h15 == _T_11317_62; // @[Mux.scala 46:19:@13034.4]
  assign _T_17586 = _T_17585 ? _T_10366_20 : _T_17584; // @[Mux.scala 46:16:@13035.4]
  assign _T_17587 = 6'h14 == _T_11317_62; // @[Mux.scala 46:19:@13036.4]
  assign _T_17588 = _T_17587 ? _T_10366_19 : _T_17586; // @[Mux.scala 46:16:@13037.4]
  assign _T_17589 = 6'h13 == _T_11317_62; // @[Mux.scala 46:19:@13038.4]
  assign _T_17590 = _T_17589 ? _T_10366_18 : _T_17588; // @[Mux.scala 46:16:@13039.4]
  assign _T_17591 = 6'h12 == _T_11317_62; // @[Mux.scala 46:19:@13040.4]
  assign _T_17592 = _T_17591 ? _T_10366_17 : _T_17590; // @[Mux.scala 46:16:@13041.4]
  assign _T_17593 = 6'h11 == _T_11317_62; // @[Mux.scala 46:19:@13042.4]
  assign _T_17594 = _T_17593 ? _T_10366_16 : _T_17592; // @[Mux.scala 46:16:@13043.4]
  assign _T_17595 = 6'h10 == _T_11317_62; // @[Mux.scala 46:19:@13044.4]
  assign _T_17596 = _T_17595 ? _T_10366_15 : _T_17594; // @[Mux.scala 46:16:@13045.4]
  assign _T_17597 = 6'hf == _T_11317_62; // @[Mux.scala 46:19:@13046.4]
  assign _T_17598 = _T_17597 ? _T_10366_14 : _T_17596; // @[Mux.scala 46:16:@13047.4]
  assign _T_17599 = 6'he == _T_11317_62; // @[Mux.scala 46:19:@13048.4]
  assign _T_17600 = _T_17599 ? _T_10366_13 : _T_17598; // @[Mux.scala 46:16:@13049.4]
  assign _T_17601 = 6'hd == _T_11317_62; // @[Mux.scala 46:19:@13050.4]
  assign _T_17602 = _T_17601 ? _T_10366_12 : _T_17600; // @[Mux.scala 46:16:@13051.4]
  assign _T_17603 = 6'hc == _T_11317_62; // @[Mux.scala 46:19:@13052.4]
  assign _T_17604 = _T_17603 ? _T_10366_11 : _T_17602; // @[Mux.scala 46:16:@13053.4]
  assign _T_17605 = 6'hb == _T_11317_62; // @[Mux.scala 46:19:@13054.4]
  assign _T_17606 = _T_17605 ? _T_10366_10 : _T_17604; // @[Mux.scala 46:16:@13055.4]
  assign _T_17607 = 6'ha == _T_11317_62; // @[Mux.scala 46:19:@13056.4]
  assign _T_17608 = _T_17607 ? _T_10366_9 : _T_17606; // @[Mux.scala 46:16:@13057.4]
  assign _T_17609 = 6'h9 == _T_11317_62; // @[Mux.scala 46:19:@13058.4]
  assign _T_17610 = _T_17609 ? _T_10366_8 : _T_17608; // @[Mux.scala 46:16:@13059.4]
  assign _T_17611 = 6'h8 == _T_11317_62; // @[Mux.scala 46:19:@13060.4]
  assign _T_17612 = _T_17611 ? _T_10366_7 : _T_17610; // @[Mux.scala 46:16:@13061.4]
  assign _T_17613 = 6'h7 == _T_11317_62; // @[Mux.scala 46:19:@13062.4]
  assign _T_17614 = _T_17613 ? _T_10366_6 : _T_17612; // @[Mux.scala 46:16:@13063.4]
  assign _T_17615 = 6'h6 == _T_11317_62; // @[Mux.scala 46:19:@13064.4]
  assign _T_17616 = _T_17615 ? _T_10366_5 : _T_17614; // @[Mux.scala 46:16:@13065.4]
  assign _T_17617 = 6'h5 == _T_11317_62; // @[Mux.scala 46:19:@13066.4]
  assign _T_17618 = _T_17617 ? _T_10366_4 : _T_17616; // @[Mux.scala 46:16:@13067.4]
  assign _T_17619 = 6'h4 == _T_11317_62; // @[Mux.scala 46:19:@13068.4]
  assign _T_17620 = _T_17619 ? _T_10366_3 : _T_17618; // @[Mux.scala 46:16:@13069.4]
  assign _T_17621 = 6'h3 == _T_11317_62; // @[Mux.scala 46:19:@13070.4]
  assign _T_17622 = _T_17621 ? _T_10366_2 : _T_17620; // @[Mux.scala 46:16:@13071.4]
  assign _T_17623 = 6'h2 == _T_11317_62; // @[Mux.scala 46:19:@13072.4]
  assign _T_17624 = _T_17623 ? _T_10366_1 : _T_17622; // @[Mux.scala 46:16:@13073.4]
  assign _T_17625 = 6'h1 == _T_11317_62; // @[Mux.scala 46:19:@13074.4]
  assign _T_17626 = _T_17625 ? _T_10366_0 : _T_17624; // @[Mux.scala 46:16:@13075.4]
  assign _T_17692 = 7'h40 == _T_11317_63; // @[Mux.scala 46:19:@13077.4]
  assign _T_17693 = _T_17692 ? _T_10366_63 : 8'h0; // @[Mux.scala 46:16:@13078.4]
  assign _T_17694 = 7'h3f == _T_11317_63; // @[Mux.scala 46:19:@13079.4]
  assign _T_17695 = _T_17694 ? _T_10366_62 : _T_17693; // @[Mux.scala 46:16:@13080.4]
  assign _T_17696 = 7'h3e == _T_11317_63; // @[Mux.scala 46:19:@13081.4]
  assign _T_17697 = _T_17696 ? _T_10366_61 : _T_17695; // @[Mux.scala 46:16:@13082.4]
  assign _T_17698 = 7'h3d == _T_11317_63; // @[Mux.scala 46:19:@13083.4]
  assign _T_17699 = _T_17698 ? _T_10366_60 : _T_17697; // @[Mux.scala 46:16:@13084.4]
  assign _T_17700 = 7'h3c == _T_11317_63; // @[Mux.scala 46:19:@13085.4]
  assign _T_17701 = _T_17700 ? _T_10366_59 : _T_17699; // @[Mux.scala 46:16:@13086.4]
  assign _T_17702 = 7'h3b == _T_11317_63; // @[Mux.scala 46:19:@13087.4]
  assign _T_17703 = _T_17702 ? _T_10366_58 : _T_17701; // @[Mux.scala 46:16:@13088.4]
  assign _T_17704 = 7'h3a == _T_11317_63; // @[Mux.scala 46:19:@13089.4]
  assign _T_17705 = _T_17704 ? _T_10366_57 : _T_17703; // @[Mux.scala 46:16:@13090.4]
  assign _T_17706 = 7'h39 == _T_11317_63; // @[Mux.scala 46:19:@13091.4]
  assign _T_17707 = _T_17706 ? _T_10366_56 : _T_17705; // @[Mux.scala 46:16:@13092.4]
  assign _T_17708 = 7'h38 == _T_11317_63; // @[Mux.scala 46:19:@13093.4]
  assign _T_17709 = _T_17708 ? _T_10366_55 : _T_17707; // @[Mux.scala 46:16:@13094.4]
  assign _T_17710 = 7'h37 == _T_11317_63; // @[Mux.scala 46:19:@13095.4]
  assign _T_17711 = _T_17710 ? _T_10366_54 : _T_17709; // @[Mux.scala 46:16:@13096.4]
  assign _T_17712 = 7'h36 == _T_11317_63; // @[Mux.scala 46:19:@13097.4]
  assign _T_17713 = _T_17712 ? _T_10366_53 : _T_17711; // @[Mux.scala 46:16:@13098.4]
  assign _T_17714 = 7'h35 == _T_11317_63; // @[Mux.scala 46:19:@13099.4]
  assign _T_17715 = _T_17714 ? _T_10366_52 : _T_17713; // @[Mux.scala 46:16:@13100.4]
  assign _T_17716 = 7'h34 == _T_11317_63; // @[Mux.scala 46:19:@13101.4]
  assign _T_17717 = _T_17716 ? _T_10366_51 : _T_17715; // @[Mux.scala 46:16:@13102.4]
  assign _T_17718 = 7'h33 == _T_11317_63; // @[Mux.scala 46:19:@13103.4]
  assign _T_17719 = _T_17718 ? _T_10366_50 : _T_17717; // @[Mux.scala 46:16:@13104.4]
  assign _T_17720 = 7'h32 == _T_11317_63; // @[Mux.scala 46:19:@13105.4]
  assign _T_17721 = _T_17720 ? _T_10366_49 : _T_17719; // @[Mux.scala 46:16:@13106.4]
  assign _T_17722 = 7'h31 == _T_11317_63; // @[Mux.scala 46:19:@13107.4]
  assign _T_17723 = _T_17722 ? _T_10366_48 : _T_17721; // @[Mux.scala 46:16:@13108.4]
  assign _T_17724 = 7'h30 == _T_11317_63; // @[Mux.scala 46:19:@13109.4]
  assign _T_17725 = _T_17724 ? _T_10366_47 : _T_17723; // @[Mux.scala 46:16:@13110.4]
  assign _T_17726 = 7'h2f == _T_11317_63; // @[Mux.scala 46:19:@13111.4]
  assign _T_17727 = _T_17726 ? _T_10366_46 : _T_17725; // @[Mux.scala 46:16:@13112.4]
  assign _T_17728 = 7'h2e == _T_11317_63; // @[Mux.scala 46:19:@13113.4]
  assign _T_17729 = _T_17728 ? _T_10366_45 : _T_17727; // @[Mux.scala 46:16:@13114.4]
  assign _T_17730 = 7'h2d == _T_11317_63; // @[Mux.scala 46:19:@13115.4]
  assign _T_17731 = _T_17730 ? _T_10366_44 : _T_17729; // @[Mux.scala 46:16:@13116.4]
  assign _T_17732 = 7'h2c == _T_11317_63; // @[Mux.scala 46:19:@13117.4]
  assign _T_17733 = _T_17732 ? _T_10366_43 : _T_17731; // @[Mux.scala 46:16:@13118.4]
  assign _T_17734 = 7'h2b == _T_11317_63; // @[Mux.scala 46:19:@13119.4]
  assign _T_17735 = _T_17734 ? _T_10366_42 : _T_17733; // @[Mux.scala 46:16:@13120.4]
  assign _T_17736 = 7'h2a == _T_11317_63; // @[Mux.scala 46:19:@13121.4]
  assign _T_17737 = _T_17736 ? _T_10366_41 : _T_17735; // @[Mux.scala 46:16:@13122.4]
  assign _T_17738 = 7'h29 == _T_11317_63; // @[Mux.scala 46:19:@13123.4]
  assign _T_17739 = _T_17738 ? _T_10366_40 : _T_17737; // @[Mux.scala 46:16:@13124.4]
  assign _T_17740 = 7'h28 == _T_11317_63; // @[Mux.scala 46:19:@13125.4]
  assign _T_17741 = _T_17740 ? _T_10366_39 : _T_17739; // @[Mux.scala 46:16:@13126.4]
  assign _T_17742 = 7'h27 == _T_11317_63; // @[Mux.scala 46:19:@13127.4]
  assign _T_17743 = _T_17742 ? _T_10366_38 : _T_17741; // @[Mux.scala 46:16:@13128.4]
  assign _T_17744 = 7'h26 == _T_11317_63; // @[Mux.scala 46:19:@13129.4]
  assign _T_17745 = _T_17744 ? _T_10366_37 : _T_17743; // @[Mux.scala 46:16:@13130.4]
  assign _T_17746 = 7'h25 == _T_11317_63; // @[Mux.scala 46:19:@13131.4]
  assign _T_17747 = _T_17746 ? _T_10366_36 : _T_17745; // @[Mux.scala 46:16:@13132.4]
  assign _T_17748 = 7'h24 == _T_11317_63; // @[Mux.scala 46:19:@13133.4]
  assign _T_17749 = _T_17748 ? _T_10366_35 : _T_17747; // @[Mux.scala 46:16:@13134.4]
  assign _T_17750 = 7'h23 == _T_11317_63; // @[Mux.scala 46:19:@13135.4]
  assign _T_17751 = _T_17750 ? _T_10366_34 : _T_17749; // @[Mux.scala 46:16:@13136.4]
  assign _T_17752 = 7'h22 == _T_11317_63; // @[Mux.scala 46:19:@13137.4]
  assign _T_17753 = _T_17752 ? _T_10366_33 : _T_17751; // @[Mux.scala 46:16:@13138.4]
  assign _T_17754 = 7'h21 == _T_11317_63; // @[Mux.scala 46:19:@13139.4]
  assign _T_17755 = _T_17754 ? _T_10366_32 : _T_17753; // @[Mux.scala 46:16:@13140.4]
  assign _T_17756 = 7'h20 == _T_11317_63; // @[Mux.scala 46:19:@13141.4]
  assign _T_17757 = _T_17756 ? _T_10366_31 : _T_17755; // @[Mux.scala 46:16:@13142.4]
  assign _T_17758 = 7'h1f == _T_11317_63; // @[Mux.scala 46:19:@13143.4]
  assign _T_17759 = _T_17758 ? _T_10366_30 : _T_17757; // @[Mux.scala 46:16:@13144.4]
  assign _T_17760 = 7'h1e == _T_11317_63; // @[Mux.scala 46:19:@13145.4]
  assign _T_17761 = _T_17760 ? _T_10366_29 : _T_17759; // @[Mux.scala 46:16:@13146.4]
  assign _T_17762 = 7'h1d == _T_11317_63; // @[Mux.scala 46:19:@13147.4]
  assign _T_17763 = _T_17762 ? _T_10366_28 : _T_17761; // @[Mux.scala 46:16:@13148.4]
  assign _T_17764 = 7'h1c == _T_11317_63; // @[Mux.scala 46:19:@13149.4]
  assign _T_17765 = _T_17764 ? _T_10366_27 : _T_17763; // @[Mux.scala 46:16:@13150.4]
  assign _T_17766 = 7'h1b == _T_11317_63; // @[Mux.scala 46:19:@13151.4]
  assign _T_17767 = _T_17766 ? _T_10366_26 : _T_17765; // @[Mux.scala 46:16:@13152.4]
  assign _T_17768 = 7'h1a == _T_11317_63; // @[Mux.scala 46:19:@13153.4]
  assign _T_17769 = _T_17768 ? _T_10366_25 : _T_17767; // @[Mux.scala 46:16:@13154.4]
  assign _T_17770 = 7'h19 == _T_11317_63; // @[Mux.scala 46:19:@13155.4]
  assign _T_17771 = _T_17770 ? _T_10366_24 : _T_17769; // @[Mux.scala 46:16:@13156.4]
  assign _T_17772 = 7'h18 == _T_11317_63; // @[Mux.scala 46:19:@13157.4]
  assign _T_17773 = _T_17772 ? _T_10366_23 : _T_17771; // @[Mux.scala 46:16:@13158.4]
  assign _T_17774 = 7'h17 == _T_11317_63; // @[Mux.scala 46:19:@13159.4]
  assign _T_17775 = _T_17774 ? _T_10366_22 : _T_17773; // @[Mux.scala 46:16:@13160.4]
  assign _T_17776 = 7'h16 == _T_11317_63; // @[Mux.scala 46:19:@13161.4]
  assign _T_17777 = _T_17776 ? _T_10366_21 : _T_17775; // @[Mux.scala 46:16:@13162.4]
  assign _T_17778 = 7'h15 == _T_11317_63; // @[Mux.scala 46:19:@13163.4]
  assign _T_17779 = _T_17778 ? _T_10366_20 : _T_17777; // @[Mux.scala 46:16:@13164.4]
  assign _T_17780 = 7'h14 == _T_11317_63; // @[Mux.scala 46:19:@13165.4]
  assign _T_17781 = _T_17780 ? _T_10366_19 : _T_17779; // @[Mux.scala 46:16:@13166.4]
  assign _T_17782 = 7'h13 == _T_11317_63; // @[Mux.scala 46:19:@13167.4]
  assign _T_17783 = _T_17782 ? _T_10366_18 : _T_17781; // @[Mux.scala 46:16:@13168.4]
  assign _T_17784 = 7'h12 == _T_11317_63; // @[Mux.scala 46:19:@13169.4]
  assign _T_17785 = _T_17784 ? _T_10366_17 : _T_17783; // @[Mux.scala 46:16:@13170.4]
  assign _T_17786 = 7'h11 == _T_11317_63; // @[Mux.scala 46:19:@13171.4]
  assign _T_17787 = _T_17786 ? _T_10366_16 : _T_17785; // @[Mux.scala 46:16:@13172.4]
  assign _T_17788 = 7'h10 == _T_11317_63; // @[Mux.scala 46:19:@13173.4]
  assign _T_17789 = _T_17788 ? _T_10366_15 : _T_17787; // @[Mux.scala 46:16:@13174.4]
  assign _T_17790 = 7'hf == _T_11317_63; // @[Mux.scala 46:19:@13175.4]
  assign _T_17791 = _T_17790 ? _T_10366_14 : _T_17789; // @[Mux.scala 46:16:@13176.4]
  assign _T_17792 = 7'he == _T_11317_63; // @[Mux.scala 46:19:@13177.4]
  assign _T_17793 = _T_17792 ? _T_10366_13 : _T_17791; // @[Mux.scala 46:16:@13178.4]
  assign _T_17794 = 7'hd == _T_11317_63; // @[Mux.scala 46:19:@13179.4]
  assign _T_17795 = _T_17794 ? _T_10366_12 : _T_17793; // @[Mux.scala 46:16:@13180.4]
  assign _T_17796 = 7'hc == _T_11317_63; // @[Mux.scala 46:19:@13181.4]
  assign _T_17797 = _T_17796 ? _T_10366_11 : _T_17795; // @[Mux.scala 46:16:@13182.4]
  assign _T_17798 = 7'hb == _T_11317_63; // @[Mux.scala 46:19:@13183.4]
  assign _T_17799 = _T_17798 ? _T_10366_10 : _T_17797; // @[Mux.scala 46:16:@13184.4]
  assign _T_17800 = 7'ha == _T_11317_63; // @[Mux.scala 46:19:@13185.4]
  assign _T_17801 = _T_17800 ? _T_10366_9 : _T_17799; // @[Mux.scala 46:16:@13186.4]
  assign _T_17802 = 7'h9 == _T_11317_63; // @[Mux.scala 46:19:@13187.4]
  assign _T_17803 = _T_17802 ? _T_10366_8 : _T_17801; // @[Mux.scala 46:16:@13188.4]
  assign _T_17804 = 7'h8 == _T_11317_63; // @[Mux.scala 46:19:@13189.4]
  assign _T_17805 = _T_17804 ? _T_10366_7 : _T_17803; // @[Mux.scala 46:16:@13190.4]
  assign _T_17806 = 7'h7 == _T_11317_63; // @[Mux.scala 46:19:@13191.4]
  assign _T_17807 = _T_17806 ? _T_10366_6 : _T_17805; // @[Mux.scala 46:16:@13192.4]
  assign _T_17808 = 7'h6 == _T_11317_63; // @[Mux.scala 46:19:@13193.4]
  assign _T_17809 = _T_17808 ? _T_10366_5 : _T_17807; // @[Mux.scala 46:16:@13194.4]
  assign _T_17810 = 7'h5 == _T_11317_63; // @[Mux.scala 46:19:@13195.4]
  assign _T_17811 = _T_17810 ? _T_10366_4 : _T_17809; // @[Mux.scala 46:16:@13196.4]
  assign _T_17812 = 7'h4 == _T_11317_63; // @[Mux.scala 46:19:@13197.4]
  assign _T_17813 = _T_17812 ? _T_10366_3 : _T_17811; // @[Mux.scala 46:16:@13198.4]
  assign _T_17814 = 7'h3 == _T_11317_63; // @[Mux.scala 46:19:@13199.4]
  assign _T_17815 = _T_17814 ? _T_10366_2 : _T_17813; // @[Mux.scala 46:16:@13200.4]
  assign _T_17816 = 7'h2 == _T_11317_63; // @[Mux.scala 46:19:@13201.4]
  assign _T_17817 = _T_17816 ? _T_10366_1 : _T_17815; // @[Mux.scala 46:16:@13202.4]
  assign _T_17818 = 7'h1 == _T_11317_63; // @[Mux.scala 46:19:@13203.4]
  assign _T_17819 = _T_17818 ? _T_10366_0 : _T_17817; // @[Mux.scala 46:16:@13204.4]
  assign _GEN_224 = _T_10362 ? _T_10641_0 : _T_17961_0; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_225 = _T_10362 ? _T_10641_1 : _T_17961_1; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_226 = _T_10362 ? _T_10641_2 : _T_17961_2; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_227 = _T_10362 ? _T_10641_3 : _T_17961_3; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_228 = _T_10362 ? _T_10641_4 : _T_17961_4; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_229 = _T_10362 ? _T_10641_5 : _T_17961_5; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_230 = _T_10362 ? _T_10641_6 : _T_17961_6; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_231 = _T_10362 ? _T_10641_7 : _T_17961_7; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_232 = _T_10362 ? _T_10641_8 : _T_17961_8; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_233 = _T_10362 ? _T_10641_9 : _T_17961_9; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_234 = _T_10362 ? _T_10641_10 : _T_17961_10; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_235 = _T_10362 ? _T_10641_11 : _T_17961_11; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_236 = _T_10362 ? _T_10641_12 : _T_17961_12; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_237 = _T_10362 ? _T_10641_13 : _T_17961_13; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_238 = _T_10362 ? _T_10641_14 : _T_17961_14; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_239 = _T_10362 ? _T_10641_15 : _T_17961_15; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_240 = _T_10362 ? _T_10641_16 : _T_17961_16; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_241 = _T_10362 ? _T_10641_17 : _T_17961_17; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_242 = _T_10362 ? _T_10641_18 : _T_17961_18; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_243 = _T_10362 ? _T_10641_19 : _T_17961_19; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_244 = _T_10362 ? _T_10641_20 : _T_17961_20; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_245 = _T_10362 ? _T_10641_21 : _T_17961_21; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_246 = _T_10362 ? _T_10641_22 : _T_17961_22; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_247 = _T_10362 ? _T_10641_23 : _T_17961_23; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_248 = _T_10362 ? _T_10641_24 : _T_17961_24; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_249 = _T_10362 ? _T_10641_25 : _T_17961_25; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_250 = _T_10362 ? _T_10641_26 : _T_17961_26; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_251 = _T_10362 ? _T_10641_27 : _T_17961_27; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_252 = _T_10362 ? _T_10641_28 : _T_17961_28; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_253 = _T_10362 ? _T_10641_29 : _T_17961_29; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_254 = _T_10362 ? _T_10641_30 : _T_17961_30; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_255 = _T_10362 ? _T_10641_31 : _T_17961_31; // @[NV_NVDLA_CSC_WL_dec.scala 99:19:@13243.4]
  assign _GEN_256 = _T_10436_0 ? _T_11519 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13278.6]
  assign _GEN_258 = _T_10436_1 ? _T_11526 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13286.6]
  assign _GEN_260 = _T_10436_2 ? _T_11536 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13294.6]
  assign _GEN_262 = _T_10436_3 ? _T_11549 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13302.6]
  assign _GEN_264 = _T_10436_4 ? _T_11565 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13310.6]
  assign _GEN_266 = _T_10436_5 ? _T_11584 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13318.6]
  assign _GEN_268 = _T_10436_6 ? _T_11606 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13326.6]
  assign _GEN_270 = _T_10436_7 ? _T_11631 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13334.6]
  assign _GEN_272 = _T_10436_8 ? _T_11659 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13342.6]
  assign _GEN_274 = _T_10436_9 ? _T_11690 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13350.6]
  assign _GEN_276 = _T_10436_10 ? _T_11724 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13358.6]
  assign _GEN_278 = _T_10436_11 ? _T_11761 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13366.6]
  assign _GEN_280 = _T_10436_12 ? _T_11801 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13374.6]
  assign _GEN_282 = _T_10436_13 ? _T_11844 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13382.6]
  assign _GEN_284 = _T_10436_14 ? _T_11890 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13390.6]
  assign _GEN_286 = _T_10436_15 ? _T_11939 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13398.6]
  assign _GEN_288 = _T_10436_16 ? _T_11991 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13406.6]
  assign _GEN_290 = _T_10436_17 ? _T_12046 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13414.6]
  assign _GEN_292 = _T_10436_18 ? _T_12104 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13422.6]
  assign _GEN_294 = _T_10436_19 ? _T_12165 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13430.6]
  assign _GEN_296 = _T_10436_20 ? _T_12229 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13438.6]
  assign _GEN_298 = _T_10436_21 ? _T_12296 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13446.6]
  assign _GEN_300 = _T_10436_22 ? _T_12366 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13454.6]
  assign _GEN_302 = _T_10436_23 ? _T_12439 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13462.6]
  assign _GEN_304 = _T_10436_24 ? _T_12515 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13470.6]
  assign _GEN_306 = _T_10436_25 ? _T_12594 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13478.6]
  assign _GEN_308 = _T_10436_26 ? _T_12676 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13486.6]
  assign _GEN_310 = _T_10436_27 ? _T_12761 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13494.6]
  assign _GEN_312 = _T_10436_28 ? _T_12849 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13502.6]
  assign _GEN_314 = _T_10436_29 ? _T_12940 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13510.6]
  assign _GEN_316 = _T_10436_30 ? _T_13034 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13518.6]
  assign _GEN_318 = _T_10436_31 ? _T_13131 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13526.6]
  assign _GEN_320 = _T_10436_32 ? _T_13231 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13534.6]
  assign _GEN_322 = _T_10436_33 ? _T_13334 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13542.6]
  assign _GEN_324 = _T_10436_34 ? _T_13440 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13550.6]
  assign _GEN_326 = _T_10436_35 ? _T_13549 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13558.6]
  assign _GEN_328 = _T_10436_36 ? _T_13661 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13566.6]
  assign _GEN_330 = _T_10436_37 ? _T_13776 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13574.6]
  assign _GEN_332 = _T_10436_38 ? _T_13894 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13582.6]
  assign _GEN_334 = _T_10436_39 ? _T_14015 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13590.6]
  assign _GEN_336 = _T_10436_40 ? _T_14139 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13598.6]
  assign _GEN_338 = _T_10436_41 ? _T_14266 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13606.6]
  assign _GEN_340 = _T_10436_42 ? _T_14396 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13614.6]
  assign _GEN_342 = _T_10436_43 ? _T_14529 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13622.6]
  assign _GEN_344 = _T_10436_44 ? _T_14665 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13630.6]
  assign _GEN_346 = _T_10436_45 ? _T_14804 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13638.6]
  assign _GEN_348 = _T_10436_46 ? _T_14946 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13646.6]
  assign _GEN_350 = _T_10436_47 ? _T_15091 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13654.6]
  assign _GEN_352 = _T_10436_48 ? _T_15239 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13662.6]
  assign _GEN_354 = _T_10436_49 ? _T_15390 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13670.6]
  assign _GEN_356 = _T_10436_50 ? _T_15544 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13678.6]
  assign _GEN_358 = _T_10436_51 ? _T_15701 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13686.6]
  assign _GEN_360 = _T_10436_52 ? _T_15861 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13694.6]
  assign _GEN_362 = _T_10436_53 ? _T_16024 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13702.6]
  assign _GEN_364 = _T_10436_54 ? _T_16190 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13710.6]
  assign _GEN_366 = _T_10436_55 ? _T_16359 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13718.6]
  assign _GEN_368 = _T_10436_56 ? _T_16531 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13726.6]
  assign _GEN_370 = _T_10436_57 ? _T_16706 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13734.6]
  assign _GEN_372 = _T_10436_58 ? _T_16884 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13742.6]
  assign _GEN_374 = _T_10436_59 ? _T_17065 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13750.6]
  assign _GEN_376 = _T_10436_60 ? _T_17249 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13758.6]
  assign _GEN_378 = _T_10436_61 ? _T_17436 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13766.6]
  assign _GEN_380 = _T_10436_62 ? _T_17626 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13774.6]
  assign _GEN_382 = _T_10436_63 ? _T_17819 : 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 104:29:@13782.6]
  assign _T_18267 = _T_11519 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13790.4]
  assign _T_18269 = _T_11526 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13792.4]
  assign _T_18271 = _T_11536 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13794.4]
  assign _T_18273 = _T_11549 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13796.4]
  assign _T_18275 = _T_11565 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13798.4]
  assign _T_18277 = _T_11584 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13800.4]
  assign _T_18279 = _T_11606 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13802.4]
  assign _T_18281 = _T_11631 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13804.4]
  assign _T_18283 = _T_11659 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13806.4]
  assign _T_18285 = _T_11690 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13808.4]
  assign _T_18287 = _T_11724 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13810.4]
  assign _T_18289 = _T_11761 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13812.4]
  assign _T_18291 = _T_11801 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13814.4]
  assign _T_18293 = _T_11844 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13816.4]
  assign _T_18295 = _T_11890 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13818.4]
  assign _T_18297 = _T_11939 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13820.4]
  assign _T_18299 = _T_11991 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13822.4]
  assign _T_18301 = _T_12046 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13824.4]
  assign _T_18303 = _T_12104 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13826.4]
  assign _T_18305 = _T_12165 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13828.4]
  assign _T_18307 = _T_12229 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13830.4]
  assign _T_18309 = _T_12296 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13832.4]
  assign _T_18311 = _T_12366 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13834.4]
  assign _T_18313 = _T_12439 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13836.4]
  assign _T_18315 = _T_12515 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13838.4]
  assign _T_18317 = _T_12594 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13840.4]
  assign _T_18319 = _T_12676 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13842.4]
  assign _T_18321 = _T_12761 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13844.4]
  assign _T_18323 = _T_12849 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13846.4]
  assign _T_18325 = _T_12940 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13848.4]
  assign _T_18327 = _T_13034 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13850.4]
  assign _T_18329 = _T_13131 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13852.4]
  assign _T_18331 = _T_13231 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13854.4]
  assign _T_18333 = _T_13334 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13856.4]
  assign _T_18335 = _T_13440 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13858.4]
  assign _T_18337 = _T_13549 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13860.4]
  assign _T_18339 = _T_13661 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13862.4]
  assign _T_18341 = _T_13776 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13864.4]
  assign _T_18343 = _T_13894 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13866.4]
  assign _T_18345 = _T_14015 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13868.4]
  assign _T_18347 = _T_14139 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13870.4]
  assign _T_18349 = _T_14266 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13872.4]
  assign _T_18351 = _T_14396 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13874.4]
  assign _T_18353 = _T_14529 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13876.4]
  assign _T_18355 = _T_14665 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13878.4]
  assign _T_18357 = _T_14804 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13880.4]
  assign _T_18359 = _T_14946 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13882.4]
  assign _T_18361 = _T_15091 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13884.4]
  assign _T_18363 = _T_15239 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13886.4]
  assign _T_18365 = _T_15390 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13888.4]
  assign _T_18367 = _T_15544 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13890.4]
  assign _T_18369 = _T_15701 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13892.4]
  assign _T_18371 = _T_15861 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13894.4]
  assign _T_18373 = _T_16024 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13896.4]
  assign _T_18375 = _T_16190 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13898.4]
  assign _T_18377 = _T_16359 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13900.4]
  assign _T_18379 = _T_16531 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13902.4]
  assign _T_18381 = _T_16706 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13904.4]
  assign _T_18383 = _T_16884 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13906.4]
  assign _T_18385 = _T_17065 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13908.4]
  assign _T_18387 = _T_17249 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13910.4]
  assign _T_18389 = _T_17436 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13912.4]
  assign _T_18391 = _T_17626 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13914.4]
  assign _T_18393 = _T_17819 != 8'h0; // @[NV_NVDLA_CSC_WL_dec.scala 117:49:@13916.4]
  assign _GEN_448 = _T_17822 ? _T_17961_0 : _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_449 = _T_17822 ? _T_17961_1 : _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_450 = _T_17822 ? _T_17961_2 : _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_451 = _T_17822 ? _T_17961_3 : _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_452 = _T_17822 ? _T_17961_4 : _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_453 = _T_17822 ? _T_17961_5 : _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_454 = _T_17822 ? _T_17961_6 : _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_455 = _T_17822 ? _T_17961_7 : _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_456 = _T_17822 ? _T_17961_8 : _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_457 = _T_17822 ? _T_17961_9 : _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_458 = _T_17822 ? _T_17961_10 : _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_459 = _T_17822 ? _T_17961_11 : _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_460 = _T_17822 ? _T_17961_12 : _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_461 = _T_17822 ? _T_17961_13 : _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_462 = _T_17822 ? _T_17961_14 : _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_463 = _T_17822 ? _T_17961_15 : _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_464 = _T_17822 ? _T_17961_16 : _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_465 = _T_17822 ? _T_17961_17 : _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_466 = _T_17822 ? _T_17961_18 : _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_467 = _T_17822 ? _T_17961_19 : _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_468 = _T_17822 ? _T_17961_20 : _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_469 = _T_17822 ? _T_17961_21 : _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_470 = _T_17822 ? _T_17961_22 : _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_471 = _T_17822 ? _T_17961_23 : _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_472 = _T_17822 ? _T_17961_24 : _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_473 = _T_17822 ? _T_17961_25 : _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_474 = _T_17822 ? _T_17961_26 : _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_475 = _T_17822 ? _T_17961_27 : _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_476 = _T_17822 ? _T_17961_28 : _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_477 = _T_17822 ? _T_17961_29 : _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_478 = _T_17822 ? _T_17961_30 : _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign _GEN_479 = _T_17822 ? _T_17961_31 : _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 128:19:@13956.4]
  assign io_output_valid = _T_18396; // @[NV_NVDLA_CSC_WL_dec.scala 135:21:@14118.4]
  assign io_output_bits_mask_0 = _T_18400_0; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14119.4]
  assign io_output_bits_mask_1 = _T_18400_1; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14120.4]
  assign io_output_bits_mask_2 = _T_18400_2; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14121.4]
  assign io_output_bits_mask_3 = _T_18400_3; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14122.4]
  assign io_output_bits_mask_4 = _T_18400_4; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14123.4]
  assign io_output_bits_mask_5 = _T_18400_5; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14124.4]
  assign io_output_bits_mask_6 = _T_18400_6; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14125.4]
  assign io_output_bits_mask_7 = _T_18400_7; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14126.4]
  assign io_output_bits_mask_8 = _T_18400_8; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14127.4]
  assign io_output_bits_mask_9 = _T_18400_9; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14128.4]
  assign io_output_bits_mask_10 = _T_18400_10; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14129.4]
  assign io_output_bits_mask_11 = _T_18400_11; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14130.4]
  assign io_output_bits_mask_12 = _T_18400_12; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14131.4]
  assign io_output_bits_mask_13 = _T_18400_13; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14132.4]
  assign io_output_bits_mask_14 = _T_18400_14; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14133.4]
  assign io_output_bits_mask_15 = _T_18400_15; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14134.4]
  assign io_output_bits_mask_16 = _T_18400_16; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14135.4]
  assign io_output_bits_mask_17 = _T_18400_17; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14136.4]
  assign io_output_bits_mask_18 = _T_18400_18; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14137.4]
  assign io_output_bits_mask_19 = _T_18400_19; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14138.4]
  assign io_output_bits_mask_20 = _T_18400_20; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14139.4]
  assign io_output_bits_mask_21 = _T_18400_21; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14140.4]
  assign io_output_bits_mask_22 = _T_18400_22; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14141.4]
  assign io_output_bits_mask_23 = _T_18400_23; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14142.4]
  assign io_output_bits_mask_24 = _T_18400_24; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14143.4]
  assign io_output_bits_mask_25 = _T_18400_25; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14144.4]
  assign io_output_bits_mask_26 = _T_18400_26; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14145.4]
  assign io_output_bits_mask_27 = _T_18400_27; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14146.4]
  assign io_output_bits_mask_28 = _T_18400_28; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14147.4]
  assign io_output_bits_mask_29 = _T_18400_29; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14148.4]
  assign io_output_bits_mask_30 = _T_18400_30; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14149.4]
  assign io_output_bits_mask_31 = _T_18400_31; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14150.4]
  assign io_output_bits_mask_32 = _T_18400_32; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14151.4]
  assign io_output_bits_mask_33 = _T_18400_33; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14152.4]
  assign io_output_bits_mask_34 = _T_18400_34; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14153.4]
  assign io_output_bits_mask_35 = _T_18400_35; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14154.4]
  assign io_output_bits_mask_36 = _T_18400_36; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14155.4]
  assign io_output_bits_mask_37 = _T_18400_37; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14156.4]
  assign io_output_bits_mask_38 = _T_18400_38; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14157.4]
  assign io_output_bits_mask_39 = _T_18400_39; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14158.4]
  assign io_output_bits_mask_40 = _T_18400_40; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14159.4]
  assign io_output_bits_mask_41 = _T_18400_41; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14160.4]
  assign io_output_bits_mask_42 = _T_18400_42; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14161.4]
  assign io_output_bits_mask_43 = _T_18400_43; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14162.4]
  assign io_output_bits_mask_44 = _T_18400_44; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14163.4]
  assign io_output_bits_mask_45 = _T_18400_45; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14164.4]
  assign io_output_bits_mask_46 = _T_18400_46; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14165.4]
  assign io_output_bits_mask_47 = _T_18400_47; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14166.4]
  assign io_output_bits_mask_48 = _T_18400_48; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14167.4]
  assign io_output_bits_mask_49 = _T_18400_49; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14168.4]
  assign io_output_bits_mask_50 = _T_18400_50; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14169.4]
  assign io_output_bits_mask_51 = _T_18400_51; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14170.4]
  assign io_output_bits_mask_52 = _T_18400_52; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14171.4]
  assign io_output_bits_mask_53 = _T_18400_53; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14172.4]
  assign io_output_bits_mask_54 = _T_18400_54; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14173.4]
  assign io_output_bits_mask_55 = _T_18400_55; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14174.4]
  assign io_output_bits_mask_56 = _T_18400_56; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14175.4]
  assign io_output_bits_mask_57 = _T_18400_57; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14176.4]
  assign io_output_bits_mask_58 = _T_18400_58; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14177.4]
  assign io_output_bits_mask_59 = _T_18400_59; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14178.4]
  assign io_output_bits_mask_60 = _T_18400_60; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14179.4]
  assign io_output_bits_mask_61 = _T_18400_61; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14180.4]
  assign io_output_bits_mask_62 = _T_18400_62; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14181.4]
  assign io_output_bits_mask_63 = _T_18400_63; // @[NV_NVDLA_CSC_WL_dec.scala 136:25:@14182.4]
  assign io_output_bits_data_0 = _T_18709_0; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14215.4]
  assign io_output_bits_data_1 = _T_18709_1; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14216.4]
  assign io_output_bits_data_2 = _T_18709_2; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14217.4]
  assign io_output_bits_data_3 = _T_18709_3; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14218.4]
  assign io_output_bits_data_4 = _T_18709_4; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14219.4]
  assign io_output_bits_data_5 = _T_18709_5; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14220.4]
  assign io_output_bits_data_6 = _T_18709_6; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14221.4]
  assign io_output_bits_data_7 = _T_18709_7; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14222.4]
  assign io_output_bits_data_8 = _T_18709_8; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14223.4]
  assign io_output_bits_data_9 = _T_18709_9; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14224.4]
  assign io_output_bits_data_10 = _T_18709_10; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14225.4]
  assign io_output_bits_data_11 = _T_18709_11; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14226.4]
  assign io_output_bits_data_12 = _T_18709_12; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14227.4]
  assign io_output_bits_data_13 = _T_18709_13; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14228.4]
  assign io_output_bits_data_14 = _T_18709_14; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14229.4]
  assign io_output_bits_data_15 = _T_18709_15; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14230.4]
  assign io_output_bits_data_16 = _T_18709_16; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14231.4]
  assign io_output_bits_data_17 = _T_18709_17; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14232.4]
  assign io_output_bits_data_18 = _T_18709_18; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14233.4]
  assign io_output_bits_data_19 = _T_18709_19; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14234.4]
  assign io_output_bits_data_20 = _T_18709_20; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14235.4]
  assign io_output_bits_data_21 = _T_18709_21; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14236.4]
  assign io_output_bits_data_22 = _T_18709_22; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14237.4]
  assign io_output_bits_data_23 = _T_18709_23; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14238.4]
  assign io_output_bits_data_24 = _T_18709_24; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14239.4]
  assign io_output_bits_data_25 = _T_18709_25; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14240.4]
  assign io_output_bits_data_26 = _T_18709_26; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14241.4]
  assign io_output_bits_data_27 = _T_18709_27; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14242.4]
  assign io_output_bits_data_28 = _T_18709_28; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14243.4]
  assign io_output_bits_data_29 = _T_18709_29; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14244.4]
  assign io_output_bits_data_30 = _T_18709_30; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14245.4]
  assign io_output_bits_data_31 = _T_18709_31; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14246.4]
  assign io_output_bits_data_32 = _T_18709_32; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14247.4]
  assign io_output_bits_data_33 = _T_18709_33; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14248.4]
  assign io_output_bits_data_34 = _T_18709_34; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14249.4]
  assign io_output_bits_data_35 = _T_18709_35; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14250.4]
  assign io_output_bits_data_36 = _T_18709_36; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14251.4]
  assign io_output_bits_data_37 = _T_18709_37; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14252.4]
  assign io_output_bits_data_38 = _T_18709_38; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14253.4]
  assign io_output_bits_data_39 = _T_18709_39; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14254.4]
  assign io_output_bits_data_40 = _T_18709_40; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14255.4]
  assign io_output_bits_data_41 = _T_18709_41; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14256.4]
  assign io_output_bits_data_42 = _T_18709_42; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14257.4]
  assign io_output_bits_data_43 = _T_18709_43; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14258.4]
  assign io_output_bits_data_44 = _T_18709_44; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14259.4]
  assign io_output_bits_data_45 = _T_18709_45; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14260.4]
  assign io_output_bits_data_46 = _T_18709_46; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14261.4]
  assign io_output_bits_data_47 = _T_18709_47; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14262.4]
  assign io_output_bits_data_48 = _T_18709_48; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14263.4]
  assign io_output_bits_data_49 = _T_18709_49; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14264.4]
  assign io_output_bits_data_50 = _T_18709_50; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14265.4]
  assign io_output_bits_data_51 = _T_18709_51; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14266.4]
  assign io_output_bits_data_52 = _T_18709_52; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14267.4]
  assign io_output_bits_data_53 = _T_18709_53; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14268.4]
  assign io_output_bits_data_54 = _T_18709_54; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14269.4]
  assign io_output_bits_data_55 = _T_18709_55; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14270.4]
  assign io_output_bits_data_56 = _T_18709_56; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14271.4]
  assign io_output_bits_data_57 = _T_18709_57; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14272.4]
  assign io_output_bits_data_58 = _T_18709_58; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14273.4]
  assign io_output_bits_data_59 = _T_18709_59; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14274.4]
  assign io_output_bits_data_60 = _T_18709_60; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14275.4]
  assign io_output_bits_data_61 = _T_18709_61; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14276.4]
  assign io_output_bits_data_62 = _T_18709_62; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14277.4]
  assign io_output_bits_data_63 = _T_18709_63; // @[NV_NVDLA_CSC_WL_dec.scala 138:25:@14278.4]
  assign io_output_bits_sel_0 = _T_18605_0; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14183.4]
  assign io_output_bits_sel_1 = _T_18605_1; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14184.4]
  assign io_output_bits_sel_2 = _T_18605_2; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14185.4]
  assign io_output_bits_sel_3 = _T_18605_3; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14186.4]
  assign io_output_bits_sel_4 = _T_18605_4; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14187.4]
  assign io_output_bits_sel_5 = _T_18605_5; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14188.4]
  assign io_output_bits_sel_6 = _T_18605_6; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14189.4]
  assign io_output_bits_sel_7 = _T_18605_7; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14190.4]
  assign io_output_bits_sel_8 = _T_18605_8; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14191.4]
  assign io_output_bits_sel_9 = _T_18605_9; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14192.4]
  assign io_output_bits_sel_10 = _T_18605_10; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14193.4]
  assign io_output_bits_sel_11 = _T_18605_11; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14194.4]
  assign io_output_bits_sel_12 = _T_18605_12; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14195.4]
  assign io_output_bits_sel_13 = _T_18605_13; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14196.4]
  assign io_output_bits_sel_14 = _T_18605_14; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14197.4]
  assign io_output_bits_sel_15 = _T_18605_15; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14198.4]
  assign io_output_bits_sel_16 = _T_18605_16; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14199.4]
  assign io_output_bits_sel_17 = _T_18605_17; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14200.4]
  assign io_output_bits_sel_18 = _T_18605_18; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14201.4]
  assign io_output_bits_sel_19 = _T_18605_19; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14202.4]
  assign io_output_bits_sel_20 = _T_18605_20; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14203.4]
  assign io_output_bits_sel_21 = _T_18605_21; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14204.4]
  assign io_output_bits_sel_22 = _T_18605_22; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14205.4]
  assign io_output_bits_sel_23 = _T_18605_23; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14206.4]
  assign io_output_bits_sel_24 = _T_18605_24; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14207.4]
  assign io_output_bits_sel_25 = _T_18605_25; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14208.4]
  assign io_output_bits_sel_26 = _T_18605_26; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14209.4]
  assign io_output_bits_sel_27 = _T_18605_27; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14210.4]
  assign io_output_bits_sel_28 = _T_18605_28; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14211.4]
  assign io_output_bits_sel_29 = _T_18605_29; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14212.4]
  assign io_output_bits_sel_30 = _T_18605_30; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14213.4]
  assign io_output_bits_sel_31 = _T_18605_31; // @[NV_NVDLA_CSC_WL_dec.scala 137:24:@14214.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_10362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_10366_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_10366_1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_10366_2 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_10366_3 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_10366_4 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_10366_5 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_10366_6 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_10366_7 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_10366_8 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10366_9 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_10366_10 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_10366_11 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_10366_12 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_10366_13 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_10366_14 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_10366_15 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_10366_16 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_10366_17 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_10366_18 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_10366_19 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_10366_20 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_10366_21 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_10366_22 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_10366_23 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_10366_24 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_10366_25 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_10366_26 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_10366_27 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_10366_28 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_10366_29 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_10366_30 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_10366_31 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_10366_32 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_10366_33 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_10366_34 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_10366_35 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_10366_36 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_10366_37 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_10366_38 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_10366_39 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_10366_40 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_10366_41 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_10366_42 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_10366_43 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_10366_44 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_10366_45 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_10366_46 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_10366_47 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_10366_48 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_10366_49 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_10366_50 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_10366_51 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_10366_52 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_10366_53 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_10366_54 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_10366_55 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_10366_56 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_10366_57 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_10366_58 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_10366_59 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_10366_60 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_10366_61 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_10366_62 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_10366_63 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_10436_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_10436_1 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_10436_2 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_10436_3 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_10436_4 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_10436_5 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_10436_6 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_10436_7 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_10436_8 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_10436_9 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_10436_10 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_10436_11 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_10436_12 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_10436_13 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_10436_14 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_10436_15 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_10436_16 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_10436_17 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_10436_18 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_10436_19 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_10436_20 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_10436_21 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_10436_22 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_10436_23 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_10436_24 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_10436_25 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_10436_26 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_10436_27 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_10436_28 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_10436_29 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_10436_30 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_10436_31 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_10436_32 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_10436_33 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_10436_34 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_10436_35 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_10436_36 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_10436_37 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_10436_38 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_10436_39 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_10436_40 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_10436_41 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_10436_42 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_10436_43 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_10436_44 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_10436_45 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_10436_46 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_10436_47 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_10436_48 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_10436_49 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_10436_50 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_10436_51 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_10436_52 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_10436_53 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_10436_54 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_10436_55 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_10436_56 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_10436_57 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_10436_58 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_10436_59 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_10436_60 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_10436_61 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_10436_62 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_10436_63 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_10641_0 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_10641_1 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_10641_2 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_10641_3 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_10641_4 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_10641_5 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_10641_6 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_10641_7 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_10641_8 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_10641_9 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_10641_10 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_10641_11 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_10641_12 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_10641_13 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_10641_14 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_10641_15 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_10641_16 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_10641_17 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_10641_18 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_10641_19 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_10641_20 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_10641_21 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_10641_22 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_10641_23 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_10641_24 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_10641_25 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_10641_26 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_10641_27 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_10641_28 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_10641_29 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_10641_30 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_10641_31 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_11317_63 = _RAND_161[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_11317_62 = _RAND_162[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_11317_61 = _RAND_163[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_11317_60 = _RAND_164[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_11317_59 = _RAND_165[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_11317_58 = _RAND_166[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_11317_57 = _RAND_167[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_11317_56 = _RAND_168[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_11317_55 = _RAND_169[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_11317_54 = _RAND_170[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_11317_53 = _RAND_171[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_11317_52 = _RAND_172[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_11317_51 = _RAND_173[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_11317_50 = _RAND_174[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_11317_49 = _RAND_175[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_11317_48 = _RAND_176[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_11317_47 = _RAND_177[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_11317_46 = _RAND_178[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_11317_45 = _RAND_179[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_11317_44 = _RAND_180[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_11317_43 = _RAND_181[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_11317_42 = _RAND_182[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_11317_41 = _RAND_183[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_11317_40 = _RAND_184[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_11317_39 = _RAND_185[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_11317_38 = _RAND_186[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_11317_37 = _RAND_187[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_11317_36 = _RAND_188[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_11317_35 = _RAND_189[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_11317_34 = _RAND_190[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_11317_33 = _RAND_191[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_11317_32 = _RAND_192[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_11317_31 = _RAND_193[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_11317_30 = _RAND_194[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_11317_29 = _RAND_195[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_11317_28 = _RAND_196[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_11317_27 = _RAND_197[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_11317_26 = _RAND_198[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_11317_25 = _RAND_199[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_11317_24 = _RAND_200[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_11317_23 = _RAND_201[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_11317_22 = _RAND_202[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_11317_21 = _RAND_203[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_11317_20 = _RAND_204[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_11317_19 = _RAND_205[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_11317_18 = _RAND_206[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_11317_17 = _RAND_207[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_11317_16 = _RAND_208[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_11317_15 = _RAND_209[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_11317_14 = _RAND_210[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_11317_13 = _RAND_211[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_11317_12 = _RAND_212[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_11317_11 = _RAND_213[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_11317_10 = _RAND_214[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_11317_9 = _RAND_215[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_11317_8 = _RAND_216[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_11317_7 = _RAND_217[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_11317_6 = _RAND_218[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_11317_5 = _RAND_219[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_11317_4 = _RAND_220[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_11317_3 = _RAND_221[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_11317_2 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_11317_1 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_11317_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_17822 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_17961_0 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_17961_1 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_17961_2 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_17961_3 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_17961_4 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_17961_5 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_17961_6 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_17961_7 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_17961_8 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_17961_9 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_17961_10 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_17961_11 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_17961_12 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_17961_13 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_17961_14 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_17961_15 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_17961_16 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_17961_17 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_17961_18 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_17961_19 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_17961_20 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_17961_21 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_17961_22 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_17961_23 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_17961_24 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_17961_25 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_17961_26 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_17961_27 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_17961_28 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_17961_29 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_17961_30 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_17961_31 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_18065_0 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_18065_1 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_18065_2 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_18065_3 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_18065_4 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_18065_5 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_18065_6 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_18065_7 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_18065_8 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_18065_9 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_18065_10 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_18065_11 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_18065_12 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_18065_13 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_18065_14 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_18065_15 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_18065_16 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_18065_17 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_18065_18 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_18065_19 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_18065_20 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_18065_21 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_18065_22 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_18065_23 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_18065_24 = _RAND_282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_18065_25 = _RAND_283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_18065_26 = _RAND_284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_18065_27 = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_18065_28 = _RAND_286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_18065_29 = _RAND_287[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_18065_30 = _RAND_288[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_18065_31 = _RAND_289[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_18065_32 = _RAND_290[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_18065_33 = _RAND_291[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_18065_34 = _RAND_292[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_18065_35 = _RAND_293[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_18065_36 = _RAND_294[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_18065_37 = _RAND_295[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_18065_38 = _RAND_296[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_18065_39 = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_18065_40 = _RAND_298[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_18065_41 = _RAND_299[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_18065_42 = _RAND_300[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_18065_43 = _RAND_301[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_18065_44 = _RAND_302[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_18065_45 = _RAND_303[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_18065_46 = _RAND_304[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_18065_47 = _RAND_305[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_18065_48 = _RAND_306[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_18065_49 = _RAND_307[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_18065_50 = _RAND_308[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_18065_51 = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_18065_52 = _RAND_310[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_18065_53 = _RAND_311[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_18065_54 = _RAND_312[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_18065_55 = _RAND_313[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_18065_56 = _RAND_314[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_18065_57 = _RAND_315[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_18065_58 = _RAND_316[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_18065_59 = _RAND_317[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_18065_60 = _RAND_318[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_18065_61 = _RAND_319[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_18065_62 = _RAND_320[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_18065_63 = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_18396 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_18400_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_18400_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_18400_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_18400_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_18400_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_18400_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_18400_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_18400_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_18400_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_18400_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_18400_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_18400_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_18400_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_18400_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_18400_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_18400_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_18400_16 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_18400_17 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_18400_18 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_18400_19 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_18400_20 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_18400_21 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_18400_22 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_18400_23 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_18400_24 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_18400_25 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_18400_26 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_18400_27 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_18400_28 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_18400_29 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_18400_30 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_18400_31 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_18400_32 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_18400_33 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_18400_34 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_18400_35 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_18400_36 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_18400_37 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_18400_38 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_18400_39 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_18400_40 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_18400_41 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_18400_42 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_18400_43 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_18400_44 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_18400_45 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_18400_46 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_18400_47 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_18400_48 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_18400_49 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_18400_50 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_18400_51 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_18400_52 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_18400_53 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_18400_54 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_18400_55 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_18400_56 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_18400_57 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_18400_58 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_18400_59 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_18400_60 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_18400_61 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_18400_62 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_18400_63 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_18605_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_18605_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_18605_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_18605_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_18605_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_18605_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_18605_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_18605_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_18605_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_18605_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_18605_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_18605_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_18605_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_18605_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_18605_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_18605_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_18605_16 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_18605_17 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_18605_18 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_18605_19 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_18605_20 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_18605_21 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_18605_22 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_18605_23 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_18605_24 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_18605_25 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_18605_26 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_18605_27 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_18605_28 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_18605_29 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_18605_30 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_18605_31 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_18709_0 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_18709_1 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_18709_2 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_18709_3 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_18709_4 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_18709_5 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_18709_6 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_18709_7 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_18709_8 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_18709_9 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_18709_10 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_18709_11 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_18709_12 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_18709_13 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_18709_14 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_18709_15 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_18709_16 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_18709_17 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_18709_18 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_18709_19 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_18709_20 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_18709_21 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_18709_22 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_18709_23 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_18709_24 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_18709_25 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_18709_26 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_18709_27 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_18709_28 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_18709_29 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_18709_30 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_18709_31 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_18709_32 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_18709_33 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_18709_34 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_18709_35 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_18709_36 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_18709_37 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_18709_38 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_18709_39 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_18709_40 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_18709_41 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_18709_42 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_18709_43 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_18709_44 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_18709_45 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_18709_46 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_18709_47 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_18709_48 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_18709_49 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_18709_50 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_18709_51 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_18709_52 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_18709_53 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_18709_54 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_18709_55 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_18709_56 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_18709_57 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_18709_58 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_18709_59 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_18709_60 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_18709_61 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_18709_62 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_18709_63 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_10362 <= 1'h0;
    end else begin
      _T_10362 <= io_input_valid;
    end
    if (io_input_valid) begin
      _T_10366_0 <= io_input_bits_data_0;
    end
    if (io_input_valid) begin
      _T_10366_1 <= io_input_bits_data_1;
    end
    if (io_input_valid) begin
      _T_10366_2 <= io_input_bits_data_2;
    end
    if (io_input_valid) begin
      _T_10366_3 <= io_input_bits_data_3;
    end
    if (io_input_valid) begin
      _T_10366_4 <= io_input_bits_data_4;
    end
    if (io_input_valid) begin
      _T_10366_5 <= io_input_bits_data_5;
    end
    if (io_input_valid) begin
      _T_10366_6 <= io_input_bits_data_6;
    end
    if (io_input_valid) begin
      _T_10366_7 <= io_input_bits_data_7;
    end
    if (io_input_valid) begin
      _T_10366_8 <= io_input_bits_data_8;
    end
    if (io_input_valid) begin
      _T_10366_9 <= io_input_bits_data_9;
    end
    if (io_input_valid) begin
      _T_10366_10 <= io_input_bits_data_10;
    end
    if (io_input_valid) begin
      _T_10366_11 <= io_input_bits_data_11;
    end
    if (io_input_valid) begin
      _T_10366_12 <= io_input_bits_data_12;
    end
    if (io_input_valid) begin
      _T_10366_13 <= io_input_bits_data_13;
    end
    if (io_input_valid) begin
      _T_10366_14 <= io_input_bits_data_14;
    end
    if (io_input_valid) begin
      _T_10366_15 <= io_input_bits_data_15;
    end
    if (io_input_valid) begin
      _T_10366_16 <= io_input_bits_data_16;
    end
    if (io_input_valid) begin
      _T_10366_17 <= io_input_bits_data_17;
    end
    if (io_input_valid) begin
      _T_10366_18 <= io_input_bits_data_18;
    end
    if (io_input_valid) begin
      _T_10366_19 <= io_input_bits_data_19;
    end
    if (io_input_valid) begin
      _T_10366_20 <= io_input_bits_data_20;
    end
    if (io_input_valid) begin
      _T_10366_21 <= io_input_bits_data_21;
    end
    if (io_input_valid) begin
      _T_10366_22 <= io_input_bits_data_22;
    end
    if (io_input_valid) begin
      _T_10366_23 <= io_input_bits_data_23;
    end
    if (io_input_valid) begin
      _T_10366_24 <= io_input_bits_data_24;
    end
    if (io_input_valid) begin
      _T_10366_25 <= io_input_bits_data_25;
    end
    if (io_input_valid) begin
      _T_10366_26 <= io_input_bits_data_26;
    end
    if (io_input_valid) begin
      _T_10366_27 <= io_input_bits_data_27;
    end
    if (io_input_valid) begin
      _T_10366_28 <= io_input_bits_data_28;
    end
    if (io_input_valid) begin
      _T_10366_29 <= io_input_bits_data_29;
    end
    if (io_input_valid) begin
      _T_10366_30 <= io_input_bits_data_30;
    end
    if (io_input_valid) begin
      _T_10366_31 <= io_input_bits_data_31;
    end
    if (io_input_valid) begin
      _T_10366_32 <= io_input_bits_data_32;
    end
    if (io_input_valid) begin
      _T_10366_33 <= io_input_bits_data_33;
    end
    if (io_input_valid) begin
      _T_10366_34 <= io_input_bits_data_34;
    end
    if (io_input_valid) begin
      _T_10366_35 <= io_input_bits_data_35;
    end
    if (io_input_valid) begin
      _T_10366_36 <= io_input_bits_data_36;
    end
    if (io_input_valid) begin
      _T_10366_37 <= io_input_bits_data_37;
    end
    if (io_input_valid) begin
      _T_10366_38 <= io_input_bits_data_38;
    end
    if (io_input_valid) begin
      _T_10366_39 <= io_input_bits_data_39;
    end
    if (io_input_valid) begin
      _T_10366_40 <= io_input_bits_data_40;
    end
    if (io_input_valid) begin
      _T_10366_41 <= io_input_bits_data_41;
    end
    if (io_input_valid) begin
      _T_10366_42 <= io_input_bits_data_42;
    end
    if (io_input_valid) begin
      _T_10366_43 <= io_input_bits_data_43;
    end
    if (io_input_valid) begin
      _T_10366_44 <= io_input_bits_data_44;
    end
    if (io_input_valid) begin
      _T_10366_45 <= io_input_bits_data_45;
    end
    if (io_input_valid) begin
      _T_10366_46 <= io_input_bits_data_46;
    end
    if (io_input_valid) begin
      _T_10366_47 <= io_input_bits_data_47;
    end
    if (io_input_valid) begin
      _T_10366_48 <= io_input_bits_data_48;
    end
    if (io_input_valid) begin
      _T_10366_49 <= io_input_bits_data_49;
    end
    if (io_input_valid) begin
      _T_10366_50 <= io_input_bits_data_50;
    end
    if (io_input_valid) begin
      _T_10366_51 <= io_input_bits_data_51;
    end
    if (io_input_valid) begin
      _T_10366_52 <= io_input_bits_data_52;
    end
    if (io_input_valid) begin
      _T_10366_53 <= io_input_bits_data_53;
    end
    if (io_input_valid) begin
      _T_10366_54 <= io_input_bits_data_54;
    end
    if (io_input_valid) begin
      _T_10366_55 <= io_input_bits_data_55;
    end
    if (io_input_valid) begin
      _T_10366_56 <= io_input_bits_data_56;
    end
    if (io_input_valid) begin
      _T_10366_57 <= io_input_bits_data_57;
    end
    if (io_input_valid) begin
      _T_10366_58 <= io_input_bits_data_58;
    end
    if (io_input_valid) begin
      _T_10366_59 <= io_input_bits_data_59;
    end
    if (io_input_valid) begin
      _T_10366_60 <= io_input_bits_data_60;
    end
    if (io_input_valid) begin
      _T_10366_61 <= io_input_bits_data_61;
    end
    if (io_input_valid) begin
      _T_10366_62 <= io_input_bits_data_62;
    end
    if (io_input_valid) begin
      _T_10366_63 <= io_input_bits_data_63;
    end
    if (io_input_valid) begin
      _T_10436_0 <= io_input_bits_mask_0;
    end
    if (io_input_valid) begin
      _T_10436_1 <= io_input_bits_mask_1;
    end
    if (io_input_valid) begin
      _T_10436_2 <= io_input_bits_mask_2;
    end
    if (io_input_valid) begin
      _T_10436_3 <= io_input_bits_mask_3;
    end
    if (io_input_valid) begin
      _T_10436_4 <= io_input_bits_mask_4;
    end
    if (io_input_valid) begin
      _T_10436_5 <= io_input_bits_mask_5;
    end
    if (io_input_valid) begin
      _T_10436_6 <= io_input_bits_mask_6;
    end
    if (io_input_valid) begin
      _T_10436_7 <= io_input_bits_mask_7;
    end
    if (io_input_valid) begin
      _T_10436_8 <= io_input_bits_mask_8;
    end
    if (io_input_valid) begin
      _T_10436_9 <= io_input_bits_mask_9;
    end
    if (io_input_valid) begin
      _T_10436_10 <= io_input_bits_mask_10;
    end
    if (io_input_valid) begin
      _T_10436_11 <= io_input_bits_mask_11;
    end
    if (io_input_valid) begin
      _T_10436_12 <= io_input_bits_mask_12;
    end
    if (io_input_valid) begin
      _T_10436_13 <= io_input_bits_mask_13;
    end
    if (io_input_valid) begin
      _T_10436_14 <= io_input_bits_mask_14;
    end
    if (io_input_valid) begin
      _T_10436_15 <= io_input_bits_mask_15;
    end
    if (io_input_valid) begin
      _T_10436_16 <= io_input_bits_mask_16;
    end
    if (io_input_valid) begin
      _T_10436_17 <= io_input_bits_mask_17;
    end
    if (io_input_valid) begin
      _T_10436_18 <= io_input_bits_mask_18;
    end
    if (io_input_valid) begin
      _T_10436_19 <= io_input_bits_mask_19;
    end
    if (io_input_valid) begin
      _T_10436_20 <= io_input_bits_mask_20;
    end
    if (io_input_valid) begin
      _T_10436_21 <= io_input_bits_mask_21;
    end
    if (io_input_valid) begin
      _T_10436_22 <= io_input_bits_mask_22;
    end
    if (io_input_valid) begin
      _T_10436_23 <= io_input_bits_mask_23;
    end
    if (io_input_valid) begin
      _T_10436_24 <= io_input_bits_mask_24;
    end
    if (io_input_valid) begin
      _T_10436_25 <= io_input_bits_mask_25;
    end
    if (io_input_valid) begin
      _T_10436_26 <= io_input_bits_mask_26;
    end
    if (io_input_valid) begin
      _T_10436_27 <= io_input_bits_mask_27;
    end
    if (io_input_valid) begin
      _T_10436_28 <= io_input_bits_mask_28;
    end
    if (io_input_valid) begin
      _T_10436_29 <= io_input_bits_mask_29;
    end
    if (io_input_valid) begin
      _T_10436_30 <= io_input_bits_mask_30;
    end
    if (io_input_valid) begin
      _T_10436_31 <= io_input_bits_mask_31;
    end
    if (io_input_valid) begin
      _T_10436_32 <= io_input_bits_mask_32;
    end
    if (io_input_valid) begin
      _T_10436_33 <= io_input_bits_mask_33;
    end
    if (io_input_valid) begin
      _T_10436_34 <= io_input_bits_mask_34;
    end
    if (io_input_valid) begin
      _T_10436_35 <= io_input_bits_mask_35;
    end
    if (io_input_valid) begin
      _T_10436_36 <= io_input_bits_mask_36;
    end
    if (io_input_valid) begin
      _T_10436_37 <= io_input_bits_mask_37;
    end
    if (io_input_valid) begin
      _T_10436_38 <= io_input_bits_mask_38;
    end
    if (io_input_valid) begin
      _T_10436_39 <= io_input_bits_mask_39;
    end
    if (io_input_valid) begin
      _T_10436_40 <= io_input_bits_mask_40;
    end
    if (io_input_valid) begin
      _T_10436_41 <= io_input_bits_mask_41;
    end
    if (io_input_valid) begin
      _T_10436_42 <= io_input_bits_mask_42;
    end
    if (io_input_valid) begin
      _T_10436_43 <= io_input_bits_mask_43;
    end
    if (io_input_valid) begin
      _T_10436_44 <= io_input_bits_mask_44;
    end
    if (io_input_valid) begin
      _T_10436_45 <= io_input_bits_mask_45;
    end
    if (io_input_valid) begin
      _T_10436_46 <= io_input_bits_mask_46;
    end
    if (io_input_valid) begin
      _T_10436_47 <= io_input_bits_mask_47;
    end
    if (io_input_valid) begin
      _T_10436_48 <= io_input_bits_mask_48;
    end
    if (io_input_valid) begin
      _T_10436_49 <= io_input_bits_mask_49;
    end
    if (io_input_valid) begin
      _T_10436_50 <= io_input_bits_mask_50;
    end
    if (io_input_valid) begin
      _T_10436_51 <= io_input_bits_mask_51;
    end
    if (io_input_valid) begin
      _T_10436_52 <= io_input_bits_mask_52;
    end
    if (io_input_valid) begin
      _T_10436_53 <= io_input_bits_mask_53;
    end
    if (io_input_valid) begin
      _T_10436_54 <= io_input_bits_mask_54;
    end
    if (io_input_valid) begin
      _T_10436_55 <= io_input_bits_mask_55;
    end
    if (io_input_valid) begin
      _T_10436_56 <= io_input_bits_mask_56;
    end
    if (io_input_valid) begin
      _T_10436_57 <= io_input_bits_mask_57;
    end
    if (io_input_valid) begin
      _T_10436_58 <= io_input_bits_mask_58;
    end
    if (io_input_valid) begin
      _T_10436_59 <= io_input_bits_mask_59;
    end
    if (io_input_valid) begin
      _T_10436_60 <= io_input_bits_mask_60;
    end
    if (io_input_valid) begin
      _T_10436_61 <= io_input_bits_mask_61;
    end
    if (io_input_valid) begin
      _T_10436_62 <= io_input_bits_mask_62;
    end
    if (io_input_valid) begin
      _T_10436_63 <= io_input_bits_mask_63;
    end
    if (reset) begin
      _T_10641_0 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_0 <= io_input_bits_sel_0;
      end
    end
    if (reset) begin
      _T_10641_1 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_1 <= io_input_bits_sel_1;
      end
    end
    if (reset) begin
      _T_10641_2 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_2 <= io_input_bits_sel_2;
      end
    end
    if (reset) begin
      _T_10641_3 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_3 <= io_input_bits_sel_3;
      end
    end
    if (reset) begin
      _T_10641_4 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_4 <= io_input_bits_sel_4;
      end
    end
    if (reset) begin
      _T_10641_5 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_5 <= io_input_bits_sel_5;
      end
    end
    if (reset) begin
      _T_10641_6 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_6 <= io_input_bits_sel_6;
      end
    end
    if (reset) begin
      _T_10641_7 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_7 <= io_input_bits_sel_7;
      end
    end
    if (reset) begin
      _T_10641_8 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_8 <= io_input_bits_sel_8;
      end
    end
    if (reset) begin
      _T_10641_9 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_9 <= io_input_bits_sel_9;
      end
    end
    if (reset) begin
      _T_10641_10 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_10 <= io_input_bits_sel_10;
      end
    end
    if (reset) begin
      _T_10641_11 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_11 <= io_input_bits_sel_11;
      end
    end
    if (reset) begin
      _T_10641_12 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_12 <= io_input_bits_sel_12;
      end
    end
    if (reset) begin
      _T_10641_13 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_13 <= io_input_bits_sel_13;
      end
    end
    if (reset) begin
      _T_10641_14 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_14 <= io_input_bits_sel_14;
      end
    end
    if (reset) begin
      _T_10641_15 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_15 <= io_input_bits_sel_15;
      end
    end
    if (reset) begin
      _T_10641_16 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_16 <= io_input_bits_sel_16;
      end
    end
    if (reset) begin
      _T_10641_17 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_17 <= io_input_bits_sel_17;
      end
    end
    if (reset) begin
      _T_10641_18 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_18 <= io_input_bits_sel_18;
      end
    end
    if (reset) begin
      _T_10641_19 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_19 <= io_input_bits_sel_19;
      end
    end
    if (reset) begin
      _T_10641_20 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_20 <= io_input_bits_sel_20;
      end
    end
    if (reset) begin
      _T_10641_21 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_21 <= io_input_bits_sel_21;
      end
    end
    if (reset) begin
      _T_10641_22 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_22 <= io_input_bits_sel_22;
      end
    end
    if (reset) begin
      _T_10641_23 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_23 <= io_input_bits_sel_23;
      end
    end
    if (reset) begin
      _T_10641_24 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_24 <= io_input_bits_sel_24;
      end
    end
    if (reset) begin
      _T_10641_25 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_25 <= io_input_bits_sel_25;
      end
    end
    if (reset) begin
      _T_10641_26 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_26 <= io_input_bits_sel_26;
      end
    end
    if (reset) begin
      _T_10641_27 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_27 <= io_input_bits_sel_27;
      end
    end
    if (reset) begin
      _T_10641_28 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_28 <= io_input_bits_sel_28;
      end
    end
    if (reset) begin
      _T_10641_29 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_29 <= io_input_bits_sel_29;
      end
    end
    if (reset) begin
      _T_10641_30 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_30 <= io_input_bits_sel_30;
      end
    end
    if (reset) begin
      _T_10641_31 <= 1'h0;
    end else begin
      if (io_input_valid) begin
        _T_10641_31 <= io_input_bits_sel_31;
      end
    end
    if (reset) begin
      _T_11317_63 <= 7'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_63 <= _T_10359;
      end
    end
    if (reset) begin
      _T_11317_62 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_62 <= _T_2167_62;
      end
    end
    if (reset) begin
      _T_11317_61 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_61 <= _T_2167_61;
      end
    end
    if (reset) begin
      _T_11317_60 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_60 <= _T_2167_60;
      end
    end
    if (reset) begin
      _T_11317_59 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_59 <= _T_2167_59;
      end
    end
    if (reset) begin
      _T_11317_58 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_58 <= _T_2167_58;
      end
    end
    if (reset) begin
      _T_11317_57 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_57 <= _T_2167_57;
      end
    end
    if (reset) begin
      _T_11317_56 <= 6'h0;
    end else begin
      if (_T_11431) begin
        _T_11317_56 <= _T_2167_56;
      end
    end
    if (reset) begin
      _T_11317_55 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_55 <= _T_2167_55;
      end
    end
    if (reset) begin
      _T_11317_54 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_54 <= _T_2167_54;
      end
    end
    if (reset) begin
      _T_11317_53 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_53 <= _T_2167_53;
      end
    end
    if (reset) begin
      _T_11317_52 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_52 <= _T_2167_52;
      end
    end
    if (reset) begin
      _T_11317_51 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_51 <= _T_2167_51;
      end
    end
    if (reset) begin
      _T_11317_50 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_50 <= _T_2167_50;
      end
    end
    if (reset) begin
      _T_11317_49 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_49 <= _T_2167_49;
      end
    end
    if (reset) begin
      _T_11317_48 <= 6'h0;
    end else begin
      if (_T_11415) begin
        _T_11317_48 <= _T_2167_48;
      end
    end
    if (reset) begin
      _T_11317_47 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_47 <= _T_2167_47;
      end
    end
    if (reset) begin
      _T_11317_46 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_46 <= _T_2167_46;
      end
    end
    if (reset) begin
      _T_11317_45 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_45 <= _T_2167_45;
      end
    end
    if (reset) begin
      _T_11317_44 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_44 <= _T_2167_44;
      end
    end
    if (reset) begin
      _T_11317_43 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_43 <= _T_2167_43;
      end
    end
    if (reset) begin
      _T_11317_42 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_42 <= _T_2167_42;
      end
    end
    if (reset) begin
      _T_11317_41 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_41 <= _T_2167_41;
      end
    end
    if (reset) begin
      _T_11317_40 <= 6'h0;
    end else begin
      if (_T_11399) begin
        _T_11317_40 <= _T_2167_40;
      end
    end
    if (reset) begin
      _T_11317_39 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_39 <= _T_2167_39;
      end
    end
    if (reset) begin
      _T_11317_38 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_38 <= _T_2167_38;
      end
    end
    if (reset) begin
      _T_11317_37 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_37 <= _T_2167_37;
      end
    end
    if (reset) begin
      _T_11317_36 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_36 <= _T_2167_36;
      end
    end
    if (reset) begin
      _T_11317_35 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_35 <= _T_2167_35;
      end
    end
    if (reset) begin
      _T_11317_34 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_34 <= _T_2167_34;
      end
    end
    if (reset) begin
      _T_11317_33 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_33 <= _T_2167_33;
      end
    end
    if (reset) begin
      _T_11317_32 <= 6'h0;
    end else begin
      if (_T_11383) begin
        _T_11317_32 <= _T_2167_32;
      end
    end
    if (reset) begin
      _T_11317_31 <= 6'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_31 <= _T_5239;
      end
    end
    if (reset) begin
      _T_11317_30 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_30 <= _T_2167_30;
      end
    end
    if (reset) begin
      _T_11317_29 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_29 <= _T_2167_29;
      end
    end
    if (reset) begin
      _T_11317_28 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_28 <= _T_2167_28;
      end
    end
    if (reset) begin
      _T_11317_27 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_27 <= _T_2167_27;
      end
    end
    if (reset) begin
      _T_11317_26 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_26 <= _T_2167_26;
      end
    end
    if (reset) begin
      _T_11317_25 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_25 <= _T_2167_25;
      end
    end
    if (reset) begin
      _T_11317_24 <= 5'h0;
    end else begin
      if (_T_11367) begin
        _T_11317_24 <= _T_2167_24;
      end
    end
    if (reset) begin
      _T_11317_23 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_23 <= _T_2167_23;
      end
    end
    if (reset) begin
      _T_11317_22 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_22 <= _T_2167_22;
      end
    end
    if (reset) begin
      _T_11317_21 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_21 <= _T_2167_21;
      end
    end
    if (reset) begin
      _T_11317_20 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_20 <= _T_2167_20;
      end
    end
    if (reset) begin
      _T_11317_19 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_19 <= _T_2167_19;
      end
    end
    if (reset) begin
      _T_11317_18 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_18 <= _T_2167_18;
      end
    end
    if (reset) begin
      _T_11317_17 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_17 <= _T_2167_17;
      end
    end
    if (reset) begin
      _T_11317_16 <= 5'h0;
    end else begin
      if (_T_11351) begin
        _T_11317_16 <= _T_2167_16;
      end
    end
    if (reset) begin
      _T_11317_15 <= 5'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_15 <= _T_3447;
      end
    end
    if (reset) begin
      _T_11317_14 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_14 <= _T_2167_14;
      end
    end
    if (reset) begin
      _T_11317_13 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_13 <= _T_2167_13;
      end
    end
    if (reset) begin
      _T_11317_12 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_12 <= _T_2167_12;
      end
    end
    if (reset) begin
      _T_11317_11 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_11 <= _T_2167_11;
      end
    end
    if (reset) begin
      _T_11317_10 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_10 <= _T_2167_10;
      end
    end
    if (reset) begin
      _T_11317_9 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_9 <= _T_2167_9;
      end
    end
    if (reset) begin
      _T_11317_8 <= 4'h0;
    end else begin
      if (_T_11335) begin
        _T_11317_8 <= _T_2167_8;
      end
    end
    if (reset) begin
      _T_11317_7 <= 4'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_7 <= _T_2743;
      end
    end
    if (reset) begin
      _T_11317_6 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_6 <= _T_2167_6;
      end
    end
    if (reset) begin
      _T_11317_5 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_5 <= _T_2167_5;
      end
    end
    if (reset) begin
      _T_11317_4 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_4 <= _T_2167_4;
      end
    end
    if (reset) begin
      _T_11317_3 <= 3'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_3 <= _T_2439;
      end
    end
    if (reset) begin
      _T_11317_2 <= 2'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_2 <= _T_2167_2;
      end
    end
    if (reset) begin
      _T_11317_1 <= 2'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_1 <= _T_2299;
      end
    end
    if (reset) begin
      _T_11317_0 <= 1'h0;
    end else begin
      if (_T_11319) begin
        _T_11317_0 <= _T_2231;
      end
    end
    if (reset) begin
      _T_17822 <= 1'h0;
    end else begin
      _T_17822 <= _T_10362;
    end
    if (reset) begin
      _T_17961_0 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_0 <= _T_10641_0;
      end
    end
    if (reset) begin
      _T_17961_1 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_1 <= _T_10641_1;
      end
    end
    if (reset) begin
      _T_17961_2 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_2 <= _T_10641_2;
      end
    end
    if (reset) begin
      _T_17961_3 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_3 <= _T_10641_3;
      end
    end
    if (reset) begin
      _T_17961_4 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_4 <= _T_10641_4;
      end
    end
    if (reset) begin
      _T_17961_5 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_5 <= _T_10641_5;
      end
    end
    if (reset) begin
      _T_17961_6 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_6 <= _T_10641_6;
      end
    end
    if (reset) begin
      _T_17961_7 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_7 <= _T_10641_7;
      end
    end
    if (reset) begin
      _T_17961_8 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_8 <= _T_10641_8;
      end
    end
    if (reset) begin
      _T_17961_9 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_9 <= _T_10641_9;
      end
    end
    if (reset) begin
      _T_17961_10 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_10 <= _T_10641_10;
      end
    end
    if (reset) begin
      _T_17961_11 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_11 <= _T_10641_11;
      end
    end
    if (reset) begin
      _T_17961_12 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_12 <= _T_10641_12;
      end
    end
    if (reset) begin
      _T_17961_13 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_13 <= _T_10641_13;
      end
    end
    if (reset) begin
      _T_17961_14 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_14 <= _T_10641_14;
      end
    end
    if (reset) begin
      _T_17961_15 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_15 <= _T_10641_15;
      end
    end
    if (reset) begin
      _T_17961_16 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_16 <= _T_10641_16;
      end
    end
    if (reset) begin
      _T_17961_17 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_17 <= _T_10641_17;
      end
    end
    if (reset) begin
      _T_17961_18 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_18 <= _T_10641_18;
      end
    end
    if (reset) begin
      _T_17961_19 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_19 <= _T_10641_19;
      end
    end
    if (reset) begin
      _T_17961_20 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_20 <= _T_10641_20;
      end
    end
    if (reset) begin
      _T_17961_21 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_21 <= _T_10641_21;
      end
    end
    if (reset) begin
      _T_17961_22 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_22 <= _T_10641_22;
      end
    end
    if (reset) begin
      _T_17961_23 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_23 <= _T_10641_23;
      end
    end
    if (reset) begin
      _T_17961_24 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_24 <= _T_10641_24;
      end
    end
    if (reset) begin
      _T_17961_25 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_25 <= _T_10641_25;
      end
    end
    if (reset) begin
      _T_17961_26 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_26 <= _T_10641_26;
      end
    end
    if (reset) begin
      _T_17961_27 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_27 <= _T_10641_27;
      end
    end
    if (reset) begin
      _T_17961_28 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_28 <= _T_10641_28;
      end
    end
    if (reset) begin
      _T_17961_29 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_29 <= _T_10641_29;
      end
    end
    if (reset) begin
      _T_17961_30 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_30 <= _T_10641_30;
      end
    end
    if (reset) begin
      _T_17961_31 <= 1'h0;
    end else begin
      if (_T_10362) begin
        _T_17961_31 <= _T_10641_31;
      end
    end
    if (_T_10362) begin
      if (_T_10436_0) begin
        if (_T_11317_0) begin
          _T_18065_0 <= _T_10366_0;
        end else begin
          _T_18065_0 <= 8'h0;
        end
      end else begin
        _T_18065_0 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_1) begin
        if (_T_11525) begin
          _T_18065_1 <= _T_10366_0;
        end else begin
          if (_T_11523) begin
            _T_18065_1 <= _T_10366_1;
          end else begin
            _T_18065_1 <= 8'h0;
          end
        end
      end else begin
        _T_18065_1 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_2) begin
        if (_T_11535) begin
          _T_18065_2 <= _T_10366_0;
        end else begin
          if (_T_11533) begin
            _T_18065_2 <= _T_10366_1;
          end else begin
            if (_T_11531) begin
              _T_18065_2 <= _T_10366_2;
            end else begin
              _T_18065_2 <= 8'h0;
            end
          end
        end
      end else begin
        _T_18065_2 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_3) begin
        if (_T_11548) begin
          _T_18065_3 <= _T_10366_0;
        end else begin
          if (_T_11546) begin
            _T_18065_3 <= _T_10366_1;
          end else begin
            if (_T_11544) begin
              _T_18065_3 <= _T_10366_2;
            end else begin
              if (_T_11542) begin
                _T_18065_3 <= _T_10366_3;
              end else begin
                _T_18065_3 <= 8'h0;
              end
            end
          end
        end
      end else begin
        _T_18065_3 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_4) begin
        if (_T_11564) begin
          _T_18065_4 <= _T_10366_0;
        end else begin
          if (_T_11562) begin
            _T_18065_4 <= _T_10366_1;
          end else begin
            if (_T_11560) begin
              _T_18065_4 <= _T_10366_2;
            end else begin
              if (_T_11558) begin
                _T_18065_4 <= _T_10366_3;
              end else begin
                if (_T_11556) begin
                  _T_18065_4 <= _T_10366_4;
                end else begin
                  _T_18065_4 <= 8'h0;
                end
              end
            end
          end
        end
      end else begin
        _T_18065_4 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_5) begin
        if (_T_11583) begin
          _T_18065_5 <= _T_10366_0;
        end else begin
          if (_T_11581) begin
            _T_18065_5 <= _T_10366_1;
          end else begin
            if (_T_11579) begin
              _T_18065_5 <= _T_10366_2;
            end else begin
              if (_T_11577) begin
                _T_18065_5 <= _T_10366_3;
              end else begin
                if (_T_11575) begin
                  _T_18065_5 <= _T_10366_4;
                end else begin
                  if (_T_11573) begin
                    _T_18065_5 <= _T_10366_5;
                  end else begin
                    _T_18065_5 <= 8'h0;
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_5 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_6) begin
        if (_T_11605) begin
          _T_18065_6 <= _T_10366_0;
        end else begin
          if (_T_11603) begin
            _T_18065_6 <= _T_10366_1;
          end else begin
            if (_T_11601) begin
              _T_18065_6 <= _T_10366_2;
            end else begin
              if (_T_11599) begin
                _T_18065_6 <= _T_10366_3;
              end else begin
                if (_T_11597) begin
                  _T_18065_6 <= _T_10366_4;
                end else begin
                  if (_T_11595) begin
                    _T_18065_6 <= _T_10366_5;
                  end else begin
                    if (_T_11593) begin
                      _T_18065_6 <= _T_10366_6;
                    end else begin
                      _T_18065_6 <= 8'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_6 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_7) begin
        if (_T_11630) begin
          _T_18065_7 <= _T_10366_0;
        end else begin
          if (_T_11628) begin
            _T_18065_7 <= _T_10366_1;
          end else begin
            if (_T_11626) begin
              _T_18065_7 <= _T_10366_2;
            end else begin
              if (_T_11624) begin
                _T_18065_7 <= _T_10366_3;
              end else begin
                if (_T_11622) begin
                  _T_18065_7 <= _T_10366_4;
                end else begin
                  if (_T_11620) begin
                    _T_18065_7 <= _T_10366_5;
                  end else begin
                    if (_T_11618) begin
                      _T_18065_7 <= _T_10366_6;
                    end else begin
                      if (_T_11616) begin
                        _T_18065_7 <= _T_10366_7;
                      end else begin
                        _T_18065_7 <= 8'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_7 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_8) begin
        if (_T_11658) begin
          _T_18065_8 <= _T_10366_0;
        end else begin
          if (_T_11656) begin
            _T_18065_8 <= _T_10366_1;
          end else begin
            if (_T_11654) begin
              _T_18065_8 <= _T_10366_2;
            end else begin
              if (_T_11652) begin
                _T_18065_8 <= _T_10366_3;
              end else begin
                if (_T_11650) begin
                  _T_18065_8 <= _T_10366_4;
                end else begin
                  if (_T_11648) begin
                    _T_18065_8 <= _T_10366_5;
                  end else begin
                    if (_T_11646) begin
                      _T_18065_8 <= _T_10366_6;
                    end else begin
                      if (_T_11644) begin
                        _T_18065_8 <= _T_10366_7;
                      end else begin
                        if (_T_11642) begin
                          _T_18065_8 <= _T_10366_8;
                        end else begin
                          _T_18065_8 <= 8'h0;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_8 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_9) begin
        if (_T_11689) begin
          _T_18065_9 <= _T_10366_0;
        end else begin
          if (_T_11687) begin
            _T_18065_9 <= _T_10366_1;
          end else begin
            if (_T_11685) begin
              _T_18065_9 <= _T_10366_2;
            end else begin
              if (_T_11683) begin
                _T_18065_9 <= _T_10366_3;
              end else begin
                if (_T_11681) begin
                  _T_18065_9 <= _T_10366_4;
                end else begin
                  if (_T_11679) begin
                    _T_18065_9 <= _T_10366_5;
                  end else begin
                    if (_T_11677) begin
                      _T_18065_9 <= _T_10366_6;
                    end else begin
                      if (_T_11675) begin
                        _T_18065_9 <= _T_10366_7;
                      end else begin
                        if (_T_11673) begin
                          _T_18065_9 <= _T_10366_8;
                        end else begin
                          if (_T_11671) begin
                            _T_18065_9 <= _T_10366_9;
                          end else begin
                            _T_18065_9 <= 8'h0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_9 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_10) begin
        if (_T_11723) begin
          _T_18065_10 <= _T_10366_0;
        end else begin
          if (_T_11721) begin
            _T_18065_10 <= _T_10366_1;
          end else begin
            if (_T_11719) begin
              _T_18065_10 <= _T_10366_2;
            end else begin
              if (_T_11717) begin
                _T_18065_10 <= _T_10366_3;
              end else begin
                if (_T_11715) begin
                  _T_18065_10 <= _T_10366_4;
                end else begin
                  if (_T_11713) begin
                    _T_18065_10 <= _T_10366_5;
                  end else begin
                    if (_T_11711) begin
                      _T_18065_10 <= _T_10366_6;
                    end else begin
                      if (_T_11709) begin
                        _T_18065_10 <= _T_10366_7;
                      end else begin
                        if (_T_11707) begin
                          _T_18065_10 <= _T_10366_8;
                        end else begin
                          if (_T_11705) begin
                            _T_18065_10 <= _T_10366_9;
                          end else begin
                            if (_T_11703) begin
                              _T_18065_10 <= _T_10366_10;
                            end else begin
                              _T_18065_10 <= 8'h0;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_10 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_11) begin
        if (_T_11760) begin
          _T_18065_11 <= _T_10366_0;
        end else begin
          if (_T_11758) begin
            _T_18065_11 <= _T_10366_1;
          end else begin
            if (_T_11756) begin
              _T_18065_11 <= _T_10366_2;
            end else begin
              if (_T_11754) begin
                _T_18065_11 <= _T_10366_3;
              end else begin
                if (_T_11752) begin
                  _T_18065_11 <= _T_10366_4;
                end else begin
                  if (_T_11750) begin
                    _T_18065_11 <= _T_10366_5;
                  end else begin
                    if (_T_11748) begin
                      _T_18065_11 <= _T_10366_6;
                    end else begin
                      if (_T_11746) begin
                        _T_18065_11 <= _T_10366_7;
                      end else begin
                        if (_T_11744) begin
                          _T_18065_11 <= _T_10366_8;
                        end else begin
                          if (_T_11742) begin
                            _T_18065_11 <= _T_10366_9;
                          end else begin
                            if (_T_11740) begin
                              _T_18065_11 <= _T_10366_10;
                            end else begin
                              if (_T_11738) begin
                                _T_18065_11 <= _T_10366_11;
                              end else begin
                                _T_18065_11 <= 8'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_11 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_12) begin
        if (_T_11800) begin
          _T_18065_12 <= _T_10366_0;
        end else begin
          if (_T_11798) begin
            _T_18065_12 <= _T_10366_1;
          end else begin
            if (_T_11796) begin
              _T_18065_12 <= _T_10366_2;
            end else begin
              if (_T_11794) begin
                _T_18065_12 <= _T_10366_3;
              end else begin
                if (_T_11792) begin
                  _T_18065_12 <= _T_10366_4;
                end else begin
                  if (_T_11790) begin
                    _T_18065_12 <= _T_10366_5;
                  end else begin
                    if (_T_11788) begin
                      _T_18065_12 <= _T_10366_6;
                    end else begin
                      if (_T_11786) begin
                        _T_18065_12 <= _T_10366_7;
                      end else begin
                        if (_T_11784) begin
                          _T_18065_12 <= _T_10366_8;
                        end else begin
                          if (_T_11782) begin
                            _T_18065_12 <= _T_10366_9;
                          end else begin
                            if (_T_11780) begin
                              _T_18065_12 <= _T_10366_10;
                            end else begin
                              if (_T_11778) begin
                                _T_18065_12 <= _T_10366_11;
                              end else begin
                                if (_T_11776) begin
                                  _T_18065_12 <= _T_10366_12;
                                end else begin
                                  _T_18065_12 <= 8'h0;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_12 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_13) begin
        if (_T_11843) begin
          _T_18065_13 <= _T_10366_0;
        end else begin
          if (_T_11841) begin
            _T_18065_13 <= _T_10366_1;
          end else begin
            if (_T_11839) begin
              _T_18065_13 <= _T_10366_2;
            end else begin
              if (_T_11837) begin
                _T_18065_13 <= _T_10366_3;
              end else begin
                if (_T_11835) begin
                  _T_18065_13 <= _T_10366_4;
                end else begin
                  if (_T_11833) begin
                    _T_18065_13 <= _T_10366_5;
                  end else begin
                    if (_T_11831) begin
                      _T_18065_13 <= _T_10366_6;
                    end else begin
                      if (_T_11829) begin
                        _T_18065_13 <= _T_10366_7;
                      end else begin
                        if (_T_11827) begin
                          _T_18065_13 <= _T_10366_8;
                        end else begin
                          if (_T_11825) begin
                            _T_18065_13 <= _T_10366_9;
                          end else begin
                            if (_T_11823) begin
                              _T_18065_13 <= _T_10366_10;
                            end else begin
                              if (_T_11821) begin
                                _T_18065_13 <= _T_10366_11;
                              end else begin
                                if (_T_11819) begin
                                  _T_18065_13 <= _T_10366_12;
                                end else begin
                                  if (_T_11817) begin
                                    _T_18065_13 <= _T_10366_13;
                                  end else begin
                                    _T_18065_13 <= 8'h0;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_13 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_14) begin
        if (_T_11889) begin
          _T_18065_14 <= _T_10366_0;
        end else begin
          if (_T_11887) begin
            _T_18065_14 <= _T_10366_1;
          end else begin
            if (_T_11885) begin
              _T_18065_14 <= _T_10366_2;
            end else begin
              if (_T_11883) begin
                _T_18065_14 <= _T_10366_3;
              end else begin
                if (_T_11881) begin
                  _T_18065_14 <= _T_10366_4;
                end else begin
                  if (_T_11879) begin
                    _T_18065_14 <= _T_10366_5;
                  end else begin
                    if (_T_11877) begin
                      _T_18065_14 <= _T_10366_6;
                    end else begin
                      if (_T_11875) begin
                        _T_18065_14 <= _T_10366_7;
                      end else begin
                        if (_T_11873) begin
                          _T_18065_14 <= _T_10366_8;
                        end else begin
                          if (_T_11871) begin
                            _T_18065_14 <= _T_10366_9;
                          end else begin
                            if (_T_11869) begin
                              _T_18065_14 <= _T_10366_10;
                            end else begin
                              if (_T_11867) begin
                                _T_18065_14 <= _T_10366_11;
                              end else begin
                                if (_T_11865) begin
                                  _T_18065_14 <= _T_10366_12;
                                end else begin
                                  if (_T_11863) begin
                                    _T_18065_14 <= _T_10366_13;
                                  end else begin
                                    if (_T_11861) begin
                                      _T_18065_14 <= _T_10366_14;
                                    end else begin
                                      _T_18065_14 <= 8'h0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_14 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_15) begin
        if (_T_11938) begin
          _T_18065_15 <= _T_10366_0;
        end else begin
          if (_T_11936) begin
            _T_18065_15 <= _T_10366_1;
          end else begin
            if (_T_11934) begin
              _T_18065_15 <= _T_10366_2;
            end else begin
              if (_T_11932) begin
                _T_18065_15 <= _T_10366_3;
              end else begin
                if (_T_11930) begin
                  _T_18065_15 <= _T_10366_4;
                end else begin
                  if (_T_11928) begin
                    _T_18065_15 <= _T_10366_5;
                  end else begin
                    if (_T_11926) begin
                      _T_18065_15 <= _T_10366_6;
                    end else begin
                      if (_T_11924) begin
                        _T_18065_15 <= _T_10366_7;
                      end else begin
                        if (_T_11922) begin
                          _T_18065_15 <= _T_10366_8;
                        end else begin
                          if (_T_11920) begin
                            _T_18065_15 <= _T_10366_9;
                          end else begin
                            if (_T_11918) begin
                              _T_18065_15 <= _T_10366_10;
                            end else begin
                              if (_T_11916) begin
                                _T_18065_15 <= _T_10366_11;
                              end else begin
                                if (_T_11914) begin
                                  _T_18065_15 <= _T_10366_12;
                                end else begin
                                  if (_T_11912) begin
                                    _T_18065_15 <= _T_10366_13;
                                  end else begin
                                    if (_T_11910) begin
                                      _T_18065_15 <= _T_10366_14;
                                    end else begin
                                      if (_T_11908) begin
                                        _T_18065_15 <= _T_10366_15;
                                      end else begin
                                        _T_18065_15 <= 8'h0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_15 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_16) begin
        if (_T_11990) begin
          _T_18065_16 <= _T_10366_0;
        end else begin
          if (_T_11988) begin
            _T_18065_16 <= _T_10366_1;
          end else begin
            if (_T_11986) begin
              _T_18065_16 <= _T_10366_2;
            end else begin
              if (_T_11984) begin
                _T_18065_16 <= _T_10366_3;
              end else begin
                if (_T_11982) begin
                  _T_18065_16 <= _T_10366_4;
                end else begin
                  if (_T_11980) begin
                    _T_18065_16 <= _T_10366_5;
                  end else begin
                    if (_T_11978) begin
                      _T_18065_16 <= _T_10366_6;
                    end else begin
                      if (_T_11976) begin
                        _T_18065_16 <= _T_10366_7;
                      end else begin
                        if (_T_11974) begin
                          _T_18065_16 <= _T_10366_8;
                        end else begin
                          if (_T_11972) begin
                            _T_18065_16 <= _T_10366_9;
                          end else begin
                            if (_T_11970) begin
                              _T_18065_16 <= _T_10366_10;
                            end else begin
                              if (_T_11968) begin
                                _T_18065_16 <= _T_10366_11;
                              end else begin
                                if (_T_11966) begin
                                  _T_18065_16 <= _T_10366_12;
                                end else begin
                                  if (_T_11964) begin
                                    _T_18065_16 <= _T_10366_13;
                                  end else begin
                                    if (_T_11962) begin
                                      _T_18065_16 <= _T_10366_14;
                                    end else begin
                                      if (_T_11960) begin
                                        _T_18065_16 <= _T_10366_15;
                                      end else begin
                                        if (_T_11958) begin
                                          _T_18065_16 <= _T_10366_16;
                                        end else begin
                                          _T_18065_16 <= 8'h0;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_16 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_17) begin
        if (_T_12045) begin
          _T_18065_17 <= _T_10366_0;
        end else begin
          if (_T_12043) begin
            _T_18065_17 <= _T_10366_1;
          end else begin
            if (_T_12041) begin
              _T_18065_17 <= _T_10366_2;
            end else begin
              if (_T_12039) begin
                _T_18065_17 <= _T_10366_3;
              end else begin
                if (_T_12037) begin
                  _T_18065_17 <= _T_10366_4;
                end else begin
                  if (_T_12035) begin
                    _T_18065_17 <= _T_10366_5;
                  end else begin
                    if (_T_12033) begin
                      _T_18065_17 <= _T_10366_6;
                    end else begin
                      if (_T_12031) begin
                        _T_18065_17 <= _T_10366_7;
                      end else begin
                        if (_T_12029) begin
                          _T_18065_17 <= _T_10366_8;
                        end else begin
                          if (_T_12027) begin
                            _T_18065_17 <= _T_10366_9;
                          end else begin
                            if (_T_12025) begin
                              _T_18065_17 <= _T_10366_10;
                            end else begin
                              if (_T_12023) begin
                                _T_18065_17 <= _T_10366_11;
                              end else begin
                                if (_T_12021) begin
                                  _T_18065_17 <= _T_10366_12;
                                end else begin
                                  if (_T_12019) begin
                                    _T_18065_17 <= _T_10366_13;
                                  end else begin
                                    if (_T_12017) begin
                                      _T_18065_17 <= _T_10366_14;
                                    end else begin
                                      if (_T_12015) begin
                                        _T_18065_17 <= _T_10366_15;
                                      end else begin
                                        if (_T_12013) begin
                                          _T_18065_17 <= _T_10366_16;
                                        end else begin
                                          if (_T_12011) begin
                                            _T_18065_17 <= _T_10366_17;
                                          end else begin
                                            _T_18065_17 <= 8'h0;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_17 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_18) begin
        if (_T_12103) begin
          _T_18065_18 <= _T_10366_0;
        end else begin
          if (_T_12101) begin
            _T_18065_18 <= _T_10366_1;
          end else begin
            if (_T_12099) begin
              _T_18065_18 <= _T_10366_2;
            end else begin
              if (_T_12097) begin
                _T_18065_18 <= _T_10366_3;
              end else begin
                if (_T_12095) begin
                  _T_18065_18 <= _T_10366_4;
                end else begin
                  if (_T_12093) begin
                    _T_18065_18 <= _T_10366_5;
                  end else begin
                    if (_T_12091) begin
                      _T_18065_18 <= _T_10366_6;
                    end else begin
                      if (_T_12089) begin
                        _T_18065_18 <= _T_10366_7;
                      end else begin
                        if (_T_12087) begin
                          _T_18065_18 <= _T_10366_8;
                        end else begin
                          if (_T_12085) begin
                            _T_18065_18 <= _T_10366_9;
                          end else begin
                            if (_T_12083) begin
                              _T_18065_18 <= _T_10366_10;
                            end else begin
                              if (_T_12081) begin
                                _T_18065_18 <= _T_10366_11;
                              end else begin
                                if (_T_12079) begin
                                  _T_18065_18 <= _T_10366_12;
                                end else begin
                                  if (_T_12077) begin
                                    _T_18065_18 <= _T_10366_13;
                                  end else begin
                                    if (_T_12075) begin
                                      _T_18065_18 <= _T_10366_14;
                                    end else begin
                                      if (_T_12073) begin
                                        _T_18065_18 <= _T_10366_15;
                                      end else begin
                                        if (_T_12071) begin
                                          _T_18065_18 <= _T_10366_16;
                                        end else begin
                                          if (_T_12069) begin
                                            _T_18065_18 <= _T_10366_17;
                                          end else begin
                                            if (_T_12067) begin
                                              _T_18065_18 <= _T_10366_18;
                                            end else begin
                                              _T_18065_18 <= 8'h0;
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_18 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_19) begin
        if (_T_12164) begin
          _T_18065_19 <= _T_10366_0;
        end else begin
          if (_T_12162) begin
            _T_18065_19 <= _T_10366_1;
          end else begin
            if (_T_12160) begin
              _T_18065_19 <= _T_10366_2;
            end else begin
              if (_T_12158) begin
                _T_18065_19 <= _T_10366_3;
              end else begin
                if (_T_12156) begin
                  _T_18065_19 <= _T_10366_4;
                end else begin
                  if (_T_12154) begin
                    _T_18065_19 <= _T_10366_5;
                  end else begin
                    if (_T_12152) begin
                      _T_18065_19 <= _T_10366_6;
                    end else begin
                      if (_T_12150) begin
                        _T_18065_19 <= _T_10366_7;
                      end else begin
                        if (_T_12148) begin
                          _T_18065_19 <= _T_10366_8;
                        end else begin
                          if (_T_12146) begin
                            _T_18065_19 <= _T_10366_9;
                          end else begin
                            if (_T_12144) begin
                              _T_18065_19 <= _T_10366_10;
                            end else begin
                              if (_T_12142) begin
                                _T_18065_19 <= _T_10366_11;
                              end else begin
                                if (_T_12140) begin
                                  _T_18065_19 <= _T_10366_12;
                                end else begin
                                  if (_T_12138) begin
                                    _T_18065_19 <= _T_10366_13;
                                  end else begin
                                    if (_T_12136) begin
                                      _T_18065_19 <= _T_10366_14;
                                    end else begin
                                      if (_T_12134) begin
                                        _T_18065_19 <= _T_10366_15;
                                      end else begin
                                        if (_T_12132) begin
                                          _T_18065_19 <= _T_10366_16;
                                        end else begin
                                          if (_T_12130) begin
                                            _T_18065_19 <= _T_10366_17;
                                          end else begin
                                            if (_T_12128) begin
                                              _T_18065_19 <= _T_10366_18;
                                            end else begin
                                              if (_T_12126) begin
                                                _T_18065_19 <= _T_10366_19;
                                              end else begin
                                                _T_18065_19 <= 8'h0;
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_19 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_20) begin
        if (_T_12228) begin
          _T_18065_20 <= _T_10366_0;
        end else begin
          if (_T_12226) begin
            _T_18065_20 <= _T_10366_1;
          end else begin
            if (_T_12224) begin
              _T_18065_20 <= _T_10366_2;
            end else begin
              if (_T_12222) begin
                _T_18065_20 <= _T_10366_3;
              end else begin
                if (_T_12220) begin
                  _T_18065_20 <= _T_10366_4;
                end else begin
                  if (_T_12218) begin
                    _T_18065_20 <= _T_10366_5;
                  end else begin
                    if (_T_12216) begin
                      _T_18065_20 <= _T_10366_6;
                    end else begin
                      if (_T_12214) begin
                        _T_18065_20 <= _T_10366_7;
                      end else begin
                        if (_T_12212) begin
                          _T_18065_20 <= _T_10366_8;
                        end else begin
                          if (_T_12210) begin
                            _T_18065_20 <= _T_10366_9;
                          end else begin
                            if (_T_12208) begin
                              _T_18065_20 <= _T_10366_10;
                            end else begin
                              if (_T_12206) begin
                                _T_18065_20 <= _T_10366_11;
                              end else begin
                                if (_T_12204) begin
                                  _T_18065_20 <= _T_10366_12;
                                end else begin
                                  if (_T_12202) begin
                                    _T_18065_20 <= _T_10366_13;
                                  end else begin
                                    if (_T_12200) begin
                                      _T_18065_20 <= _T_10366_14;
                                    end else begin
                                      if (_T_12198) begin
                                        _T_18065_20 <= _T_10366_15;
                                      end else begin
                                        if (_T_12196) begin
                                          _T_18065_20 <= _T_10366_16;
                                        end else begin
                                          if (_T_12194) begin
                                            _T_18065_20 <= _T_10366_17;
                                          end else begin
                                            if (_T_12192) begin
                                              _T_18065_20 <= _T_10366_18;
                                            end else begin
                                              if (_T_12190) begin
                                                _T_18065_20 <= _T_10366_19;
                                              end else begin
                                                if (_T_12188) begin
                                                  _T_18065_20 <= _T_10366_20;
                                                end else begin
                                                  _T_18065_20 <= 8'h0;
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_20 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_21) begin
        if (_T_12295) begin
          _T_18065_21 <= _T_10366_0;
        end else begin
          if (_T_12293) begin
            _T_18065_21 <= _T_10366_1;
          end else begin
            if (_T_12291) begin
              _T_18065_21 <= _T_10366_2;
            end else begin
              if (_T_12289) begin
                _T_18065_21 <= _T_10366_3;
              end else begin
                if (_T_12287) begin
                  _T_18065_21 <= _T_10366_4;
                end else begin
                  if (_T_12285) begin
                    _T_18065_21 <= _T_10366_5;
                  end else begin
                    if (_T_12283) begin
                      _T_18065_21 <= _T_10366_6;
                    end else begin
                      if (_T_12281) begin
                        _T_18065_21 <= _T_10366_7;
                      end else begin
                        if (_T_12279) begin
                          _T_18065_21 <= _T_10366_8;
                        end else begin
                          if (_T_12277) begin
                            _T_18065_21 <= _T_10366_9;
                          end else begin
                            if (_T_12275) begin
                              _T_18065_21 <= _T_10366_10;
                            end else begin
                              if (_T_12273) begin
                                _T_18065_21 <= _T_10366_11;
                              end else begin
                                if (_T_12271) begin
                                  _T_18065_21 <= _T_10366_12;
                                end else begin
                                  if (_T_12269) begin
                                    _T_18065_21 <= _T_10366_13;
                                  end else begin
                                    if (_T_12267) begin
                                      _T_18065_21 <= _T_10366_14;
                                    end else begin
                                      if (_T_12265) begin
                                        _T_18065_21 <= _T_10366_15;
                                      end else begin
                                        if (_T_12263) begin
                                          _T_18065_21 <= _T_10366_16;
                                        end else begin
                                          if (_T_12261) begin
                                            _T_18065_21 <= _T_10366_17;
                                          end else begin
                                            if (_T_12259) begin
                                              _T_18065_21 <= _T_10366_18;
                                            end else begin
                                              if (_T_12257) begin
                                                _T_18065_21 <= _T_10366_19;
                                              end else begin
                                                if (_T_12255) begin
                                                  _T_18065_21 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12253) begin
                                                    _T_18065_21 <= _T_10366_21;
                                                  end else begin
                                                    _T_18065_21 <= 8'h0;
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_21 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_22) begin
        if (_T_12365) begin
          _T_18065_22 <= _T_10366_0;
        end else begin
          if (_T_12363) begin
            _T_18065_22 <= _T_10366_1;
          end else begin
            if (_T_12361) begin
              _T_18065_22 <= _T_10366_2;
            end else begin
              if (_T_12359) begin
                _T_18065_22 <= _T_10366_3;
              end else begin
                if (_T_12357) begin
                  _T_18065_22 <= _T_10366_4;
                end else begin
                  if (_T_12355) begin
                    _T_18065_22 <= _T_10366_5;
                  end else begin
                    if (_T_12353) begin
                      _T_18065_22 <= _T_10366_6;
                    end else begin
                      if (_T_12351) begin
                        _T_18065_22 <= _T_10366_7;
                      end else begin
                        if (_T_12349) begin
                          _T_18065_22 <= _T_10366_8;
                        end else begin
                          if (_T_12347) begin
                            _T_18065_22 <= _T_10366_9;
                          end else begin
                            if (_T_12345) begin
                              _T_18065_22 <= _T_10366_10;
                            end else begin
                              if (_T_12343) begin
                                _T_18065_22 <= _T_10366_11;
                              end else begin
                                if (_T_12341) begin
                                  _T_18065_22 <= _T_10366_12;
                                end else begin
                                  if (_T_12339) begin
                                    _T_18065_22 <= _T_10366_13;
                                  end else begin
                                    if (_T_12337) begin
                                      _T_18065_22 <= _T_10366_14;
                                    end else begin
                                      if (_T_12335) begin
                                        _T_18065_22 <= _T_10366_15;
                                      end else begin
                                        if (_T_12333) begin
                                          _T_18065_22 <= _T_10366_16;
                                        end else begin
                                          if (_T_12331) begin
                                            _T_18065_22 <= _T_10366_17;
                                          end else begin
                                            if (_T_12329) begin
                                              _T_18065_22 <= _T_10366_18;
                                            end else begin
                                              if (_T_12327) begin
                                                _T_18065_22 <= _T_10366_19;
                                              end else begin
                                                if (_T_12325) begin
                                                  _T_18065_22 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12323) begin
                                                    _T_18065_22 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12321) begin
                                                      _T_18065_22 <= _T_10366_22;
                                                    end else begin
                                                      _T_18065_22 <= 8'h0;
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_22 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_23) begin
        if (_T_12438) begin
          _T_18065_23 <= _T_10366_0;
        end else begin
          if (_T_12436) begin
            _T_18065_23 <= _T_10366_1;
          end else begin
            if (_T_12434) begin
              _T_18065_23 <= _T_10366_2;
            end else begin
              if (_T_12432) begin
                _T_18065_23 <= _T_10366_3;
              end else begin
                if (_T_12430) begin
                  _T_18065_23 <= _T_10366_4;
                end else begin
                  if (_T_12428) begin
                    _T_18065_23 <= _T_10366_5;
                  end else begin
                    if (_T_12426) begin
                      _T_18065_23 <= _T_10366_6;
                    end else begin
                      if (_T_12424) begin
                        _T_18065_23 <= _T_10366_7;
                      end else begin
                        if (_T_12422) begin
                          _T_18065_23 <= _T_10366_8;
                        end else begin
                          if (_T_12420) begin
                            _T_18065_23 <= _T_10366_9;
                          end else begin
                            if (_T_12418) begin
                              _T_18065_23 <= _T_10366_10;
                            end else begin
                              if (_T_12416) begin
                                _T_18065_23 <= _T_10366_11;
                              end else begin
                                if (_T_12414) begin
                                  _T_18065_23 <= _T_10366_12;
                                end else begin
                                  if (_T_12412) begin
                                    _T_18065_23 <= _T_10366_13;
                                  end else begin
                                    if (_T_12410) begin
                                      _T_18065_23 <= _T_10366_14;
                                    end else begin
                                      if (_T_12408) begin
                                        _T_18065_23 <= _T_10366_15;
                                      end else begin
                                        if (_T_12406) begin
                                          _T_18065_23 <= _T_10366_16;
                                        end else begin
                                          if (_T_12404) begin
                                            _T_18065_23 <= _T_10366_17;
                                          end else begin
                                            if (_T_12402) begin
                                              _T_18065_23 <= _T_10366_18;
                                            end else begin
                                              if (_T_12400) begin
                                                _T_18065_23 <= _T_10366_19;
                                              end else begin
                                                if (_T_12398) begin
                                                  _T_18065_23 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12396) begin
                                                    _T_18065_23 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12394) begin
                                                      _T_18065_23 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12392) begin
                                                        _T_18065_23 <= _T_10366_23;
                                                      end else begin
                                                        _T_18065_23 <= 8'h0;
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_23 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_24) begin
        if (_T_12514) begin
          _T_18065_24 <= _T_10366_0;
        end else begin
          if (_T_12512) begin
            _T_18065_24 <= _T_10366_1;
          end else begin
            if (_T_12510) begin
              _T_18065_24 <= _T_10366_2;
            end else begin
              if (_T_12508) begin
                _T_18065_24 <= _T_10366_3;
              end else begin
                if (_T_12506) begin
                  _T_18065_24 <= _T_10366_4;
                end else begin
                  if (_T_12504) begin
                    _T_18065_24 <= _T_10366_5;
                  end else begin
                    if (_T_12502) begin
                      _T_18065_24 <= _T_10366_6;
                    end else begin
                      if (_T_12500) begin
                        _T_18065_24 <= _T_10366_7;
                      end else begin
                        if (_T_12498) begin
                          _T_18065_24 <= _T_10366_8;
                        end else begin
                          if (_T_12496) begin
                            _T_18065_24 <= _T_10366_9;
                          end else begin
                            if (_T_12494) begin
                              _T_18065_24 <= _T_10366_10;
                            end else begin
                              if (_T_12492) begin
                                _T_18065_24 <= _T_10366_11;
                              end else begin
                                if (_T_12490) begin
                                  _T_18065_24 <= _T_10366_12;
                                end else begin
                                  if (_T_12488) begin
                                    _T_18065_24 <= _T_10366_13;
                                  end else begin
                                    if (_T_12486) begin
                                      _T_18065_24 <= _T_10366_14;
                                    end else begin
                                      if (_T_12484) begin
                                        _T_18065_24 <= _T_10366_15;
                                      end else begin
                                        if (_T_12482) begin
                                          _T_18065_24 <= _T_10366_16;
                                        end else begin
                                          if (_T_12480) begin
                                            _T_18065_24 <= _T_10366_17;
                                          end else begin
                                            if (_T_12478) begin
                                              _T_18065_24 <= _T_10366_18;
                                            end else begin
                                              if (_T_12476) begin
                                                _T_18065_24 <= _T_10366_19;
                                              end else begin
                                                if (_T_12474) begin
                                                  _T_18065_24 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12472) begin
                                                    _T_18065_24 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12470) begin
                                                      _T_18065_24 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12468) begin
                                                        _T_18065_24 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12466) begin
                                                          _T_18065_24 <= _T_10366_24;
                                                        end else begin
                                                          _T_18065_24 <= 8'h0;
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_24 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_25) begin
        if (_T_12593) begin
          _T_18065_25 <= _T_10366_0;
        end else begin
          if (_T_12591) begin
            _T_18065_25 <= _T_10366_1;
          end else begin
            if (_T_12589) begin
              _T_18065_25 <= _T_10366_2;
            end else begin
              if (_T_12587) begin
                _T_18065_25 <= _T_10366_3;
              end else begin
                if (_T_12585) begin
                  _T_18065_25 <= _T_10366_4;
                end else begin
                  if (_T_12583) begin
                    _T_18065_25 <= _T_10366_5;
                  end else begin
                    if (_T_12581) begin
                      _T_18065_25 <= _T_10366_6;
                    end else begin
                      if (_T_12579) begin
                        _T_18065_25 <= _T_10366_7;
                      end else begin
                        if (_T_12577) begin
                          _T_18065_25 <= _T_10366_8;
                        end else begin
                          if (_T_12575) begin
                            _T_18065_25 <= _T_10366_9;
                          end else begin
                            if (_T_12573) begin
                              _T_18065_25 <= _T_10366_10;
                            end else begin
                              if (_T_12571) begin
                                _T_18065_25 <= _T_10366_11;
                              end else begin
                                if (_T_12569) begin
                                  _T_18065_25 <= _T_10366_12;
                                end else begin
                                  if (_T_12567) begin
                                    _T_18065_25 <= _T_10366_13;
                                  end else begin
                                    if (_T_12565) begin
                                      _T_18065_25 <= _T_10366_14;
                                    end else begin
                                      if (_T_12563) begin
                                        _T_18065_25 <= _T_10366_15;
                                      end else begin
                                        if (_T_12561) begin
                                          _T_18065_25 <= _T_10366_16;
                                        end else begin
                                          if (_T_12559) begin
                                            _T_18065_25 <= _T_10366_17;
                                          end else begin
                                            if (_T_12557) begin
                                              _T_18065_25 <= _T_10366_18;
                                            end else begin
                                              if (_T_12555) begin
                                                _T_18065_25 <= _T_10366_19;
                                              end else begin
                                                if (_T_12553) begin
                                                  _T_18065_25 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12551) begin
                                                    _T_18065_25 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12549) begin
                                                      _T_18065_25 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12547) begin
                                                        _T_18065_25 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12545) begin
                                                          _T_18065_25 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12543) begin
                                                            _T_18065_25 <= _T_10366_25;
                                                          end else begin
                                                            _T_18065_25 <= 8'h0;
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_25 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_26) begin
        if (_T_12675) begin
          _T_18065_26 <= _T_10366_0;
        end else begin
          if (_T_12673) begin
            _T_18065_26 <= _T_10366_1;
          end else begin
            if (_T_12671) begin
              _T_18065_26 <= _T_10366_2;
            end else begin
              if (_T_12669) begin
                _T_18065_26 <= _T_10366_3;
              end else begin
                if (_T_12667) begin
                  _T_18065_26 <= _T_10366_4;
                end else begin
                  if (_T_12665) begin
                    _T_18065_26 <= _T_10366_5;
                  end else begin
                    if (_T_12663) begin
                      _T_18065_26 <= _T_10366_6;
                    end else begin
                      if (_T_12661) begin
                        _T_18065_26 <= _T_10366_7;
                      end else begin
                        if (_T_12659) begin
                          _T_18065_26 <= _T_10366_8;
                        end else begin
                          if (_T_12657) begin
                            _T_18065_26 <= _T_10366_9;
                          end else begin
                            if (_T_12655) begin
                              _T_18065_26 <= _T_10366_10;
                            end else begin
                              if (_T_12653) begin
                                _T_18065_26 <= _T_10366_11;
                              end else begin
                                if (_T_12651) begin
                                  _T_18065_26 <= _T_10366_12;
                                end else begin
                                  if (_T_12649) begin
                                    _T_18065_26 <= _T_10366_13;
                                  end else begin
                                    if (_T_12647) begin
                                      _T_18065_26 <= _T_10366_14;
                                    end else begin
                                      if (_T_12645) begin
                                        _T_18065_26 <= _T_10366_15;
                                      end else begin
                                        if (_T_12643) begin
                                          _T_18065_26 <= _T_10366_16;
                                        end else begin
                                          if (_T_12641) begin
                                            _T_18065_26 <= _T_10366_17;
                                          end else begin
                                            if (_T_12639) begin
                                              _T_18065_26 <= _T_10366_18;
                                            end else begin
                                              if (_T_12637) begin
                                                _T_18065_26 <= _T_10366_19;
                                              end else begin
                                                if (_T_12635) begin
                                                  _T_18065_26 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12633) begin
                                                    _T_18065_26 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12631) begin
                                                      _T_18065_26 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12629) begin
                                                        _T_18065_26 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12627) begin
                                                          _T_18065_26 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12625) begin
                                                            _T_18065_26 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12623) begin
                                                              _T_18065_26 <= _T_10366_26;
                                                            end else begin
                                                              _T_18065_26 <= 8'h0;
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_26 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_27) begin
        if (_T_12760) begin
          _T_18065_27 <= _T_10366_0;
        end else begin
          if (_T_12758) begin
            _T_18065_27 <= _T_10366_1;
          end else begin
            if (_T_12756) begin
              _T_18065_27 <= _T_10366_2;
            end else begin
              if (_T_12754) begin
                _T_18065_27 <= _T_10366_3;
              end else begin
                if (_T_12752) begin
                  _T_18065_27 <= _T_10366_4;
                end else begin
                  if (_T_12750) begin
                    _T_18065_27 <= _T_10366_5;
                  end else begin
                    if (_T_12748) begin
                      _T_18065_27 <= _T_10366_6;
                    end else begin
                      if (_T_12746) begin
                        _T_18065_27 <= _T_10366_7;
                      end else begin
                        if (_T_12744) begin
                          _T_18065_27 <= _T_10366_8;
                        end else begin
                          if (_T_12742) begin
                            _T_18065_27 <= _T_10366_9;
                          end else begin
                            if (_T_12740) begin
                              _T_18065_27 <= _T_10366_10;
                            end else begin
                              if (_T_12738) begin
                                _T_18065_27 <= _T_10366_11;
                              end else begin
                                if (_T_12736) begin
                                  _T_18065_27 <= _T_10366_12;
                                end else begin
                                  if (_T_12734) begin
                                    _T_18065_27 <= _T_10366_13;
                                  end else begin
                                    if (_T_12732) begin
                                      _T_18065_27 <= _T_10366_14;
                                    end else begin
                                      if (_T_12730) begin
                                        _T_18065_27 <= _T_10366_15;
                                      end else begin
                                        if (_T_12728) begin
                                          _T_18065_27 <= _T_10366_16;
                                        end else begin
                                          if (_T_12726) begin
                                            _T_18065_27 <= _T_10366_17;
                                          end else begin
                                            if (_T_12724) begin
                                              _T_18065_27 <= _T_10366_18;
                                            end else begin
                                              if (_T_12722) begin
                                                _T_18065_27 <= _T_10366_19;
                                              end else begin
                                                if (_T_12720) begin
                                                  _T_18065_27 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12718) begin
                                                    _T_18065_27 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12716) begin
                                                      _T_18065_27 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12714) begin
                                                        _T_18065_27 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12712) begin
                                                          _T_18065_27 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12710) begin
                                                            _T_18065_27 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12708) begin
                                                              _T_18065_27 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12706) begin
                                                                _T_18065_27 <= _T_10366_27;
                                                              end else begin
                                                                _T_18065_27 <= 8'h0;
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_27 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_28) begin
        if (_T_12848) begin
          _T_18065_28 <= _T_10366_0;
        end else begin
          if (_T_12846) begin
            _T_18065_28 <= _T_10366_1;
          end else begin
            if (_T_12844) begin
              _T_18065_28 <= _T_10366_2;
            end else begin
              if (_T_12842) begin
                _T_18065_28 <= _T_10366_3;
              end else begin
                if (_T_12840) begin
                  _T_18065_28 <= _T_10366_4;
                end else begin
                  if (_T_12838) begin
                    _T_18065_28 <= _T_10366_5;
                  end else begin
                    if (_T_12836) begin
                      _T_18065_28 <= _T_10366_6;
                    end else begin
                      if (_T_12834) begin
                        _T_18065_28 <= _T_10366_7;
                      end else begin
                        if (_T_12832) begin
                          _T_18065_28 <= _T_10366_8;
                        end else begin
                          if (_T_12830) begin
                            _T_18065_28 <= _T_10366_9;
                          end else begin
                            if (_T_12828) begin
                              _T_18065_28 <= _T_10366_10;
                            end else begin
                              if (_T_12826) begin
                                _T_18065_28 <= _T_10366_11;
                              end else begin
                                if (_T_12824) begin
                                  _T_18065_28 <= _T_10366_12;
                                end else begin
                                  if (_T_12822) begin
                                    _T_18065_28 <= _T_10366_13;
                                  end else begin
                                    if (_T_12820) begin
                                      _T_18065_28 <= _T_10366_14;
                                    end else begin
                                      if (_T_12818) begin
                                        _T_18065_28 <= _T_10366_15;
                                      end else begin
                                        if (_T_12816) begin
                                          _T_18065_28 <= _T_10366_16;
                                        end else begin
                                          if (_T_12814) begin
                                            _T_18065_28 <= _T_10366_17;
                                          end else begin
                                            if (_T_12812) begin
                                              _T_18065_28 <= _T_10366_18;
                                            end else begin
                                              if (_T_12810) begin
                                                _T_18065_28 <= _T_10366_19;
                                              end else begin
                                                if (_T_12808) begin
                                                  _T_18065_28 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12806) begin
                                                    _T_18065_28 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12804) begin
                                                      _T_18065_28 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12802) begin
                                                        _T_18065_28 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12800) begin
                                                          _T_18065_28 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12798) begin
                                                            _T_18065_28 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12796) begin
                                                              _T_18065_28 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12794) begin
                                                                _T_18065_28 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12792) begin
                                                                  _T_18065_28 <= _T_10366_28;
                                                                end else begin
                                                                  _T_18065_28 <= 8'h0;
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_28 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_29) begin
        if (_T_12939) begin
          _T_18065_29 <= _T_10366_0;
        end else begin
          if (_T_12937) begin
            _T_18065_29 <= _T_10366_1;
          end else begin
            if (_T_12935) begin
              _T_18065_29 <= _T_10366_2;
            end else begin
              if (_T_12933) begin
                _T_18065_29 <= _T_10366_3;
              end else begin
                if (_T_12931) begin
                  _T_18065_29 <= _T_10366_4;
                end else begin
                  if (_T_12929) begin
                    _T_18065_29 <= _T_10366_5;
                  end else begin
                    if (_T_12927) begin
                      _T_18065_29 <= _T_10366_6;
                    end else begin
                      if (_T_12925) begin
                        _T_18065_29 <= _T_10366_7;
                      end else begin
                        if (_T_12923) begin
                          _T_18065_29 <= _T_10366_8;
                        end else begin
                          if (_T_12921) begin
                            _T_18065_29 <= _T_10366_9;
                          end else begin
                            if (_T_12919) begin
                              _T_18065_29 <= _T_10366_10;
                            end else begin
                              if (_T_12917) begin
                                _T_18065_29 <= _T_10366_11;
                              end else begin
                                if (_T_12915) begin
                                  _T_18065_29 <= _T_10366_12;
                                end else begin
                                  if (_T_12913) begin
                                    _T_18065_29 <= _T_10366_13;
                                  end else begin
                                    if (_T_12911) begin
                                      _T_18065_29 <= _T_10366_14;
                                    end else begin
                                      if (_T_12909) begin
                                        _T_18065_29 <= _T_10366_15;
                                      end else begin
                                        if (_T_12907) begin
                                          _T_18065_29 <= _T_10366_16;
                                        end else begin
                                          if (_T_12905) begin
                                            _T_18065_29 <= _T_10366_17;
                                          end else begin
                                            if (_T_12903) begin
                                              _T_18065_29 <= _T_10366_18;
                                            end else begin
                                              if (_T_12901) begin
                                                _T_18065_29 <= _T_10366_19;
                                              end else begin
                                                if (_T_12899) begin
                                                  _T_18065_29 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12897) begin
                                                    _T_18065_29 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12895) begin
                                                      _T_18065_29 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12893) begin
                                                        _T_18065_29 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12891) begin
                                                          _T_18065_29 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12889) begin
                                                            _T_18065_29 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12887) begin
                                                              _T_18065_29 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12885) begin
                                                                _T_18065_29 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12883) begin
                                                                  _T_18065_29 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_12881) begin
                                                                    _T_18065_29 <= _T_10366_29;
                                                                  end else begin
                                                                    _T_18065_29 <= 8'h0;
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_29 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_30) begin
        if (_T_13033) begin
          _T_18065_30 <= _T_10366_0;
        end else begin
          if (_T_13031) begin
            _T_18065_30 <= _T_10366_1;
          end else begin
            if (_T_13029) begin
              _T_18065_30 <= _T_10366_2;
            end else begin
              if (_T_13027) begin
                _T_18065_30 <= _T_10366_3;
              end else begin
                if (_T_13025) begin
                  _T_18065_30 <= _T_10366_4;
                end else begin
                  if (_T_13023) begin
                    _T_18065_30 <= _T_10366_5;
                  end else begin
                    if (_T_13021) begin
                      _T_18065_30 <= _T_10366_6;
                    end else begin
                      if (_T_13019) begin
                        _T_18065_30 <= _T_10366_7;
                      end else begin
                        if (_T_13017) begin
                          _T_18065_30 <= _T_10366_8;
                        end else begin
                          if (_T_13015) begin
                            _T_18065_30 <= _T_10366_9;
                          end else begin
                            if (_T_13013) begin
                              _T_18065_30 <= _T_10366_10;
                            end else begin
                              if (_T_13011) begin
                                _T_18065_30 <= _T_10366_11;
                              end else begin
                                if (_T_13009) begin
                                  _T_18065_30 <= _T_10366_12;
                                end else begin
                                  if (_T_13007) begin
                                    _T_18065_30 <= _T_10366_13;
                                  end else begin
                                    if (_T_13005) begin
                                      _T_18065_30 <= _T_10366_14;
                                    end else begin
                                      if (_T_13003) begin
                                        _T_18065_30 <= _T_10366_15;
                                      end else begin
                                        if (_T_13001) begin
                                          _T_18065_30 <= _T_10366_16;
                                        end else begin
                                          if (_T_12999) begin
                                            _T_18065_30 <= _T_10366_17;
                                          end else begin
                                            if (_T_12997) begin
                                              _T_18065_30 <= _T_10366_18;
                                            end else begin
                                              if (_T_12995) begin
                                                _T_18065_30 <= _T_10366_19;
                                              end else begin
                                                if (_T_12993) begin
                                                  _T_18065_30 <= _T_10366_20;
                                                end else begin
                                                  if (_T_12991) begin
                                                    _T_18065_30 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_12989) begin
                                                      _T_18065_30 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_12987) begin
                                                        _T_18065_30 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_12985) begin
                                                          _T_18065_30 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_12983) begin
                                                            _T_18065_30 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_12981) begin
                                                              _T_18065_30 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_12979) begin
                                                                _T_18065_30 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_12977) begin
                                                                  _T_18065_30 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_12975) begin
                                                                    _T_18065_30 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_12973) begin
                                                                      _T_18065_30 <= _T_10366_30;
                                                                    end else begin
                                                                      _T_18065_30 <= 8'h0;
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_30 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_31) begin
        if (_T_13130) begin
          _T_18065_31 <= _T_10366_0;
        end else begin
          if (_T_13128) begin
            _T_18065_31 <= _T_10366_1;
          end else begin
            if (_T_13126) begin
              _T_18065_31 <= _T_10366_2;
            end else begin
              if (_T_13124) begin
                _T_18065_31 <= _T_10366_3;
              end else begin
                if (_T_13122) begin
                  _T_18065_31 <= _T_10366_4;
                end else begin
                  if (_T_13120) begin
                    _T_18065_31 <= _T_10366_5;
                  end else begin
                    if (_T_13118) begin
                      _T_18065_31 <= _T_10366_6;
                    end else begin
                      if (_T_13116) begin
                        _T_18065_31 <= _T_10366_7;
                      end else begin
                        if (_T_13114) begin
                          _T_18065_31 <= _T_10366_8;
                        end else begin
                          if (_T_13112) begin
                            _T_18065_31 <= _T_10366_9;
                          end else begin
                            if (_T_13110) begin
                              _T_18065_31 <= _T_10366_10;
                            end else begin
                              if (_T_13108) begin
                                _T_18065_31 <= _T_10366_11;
                              end else begin
                                if (_T_13106) begin
                                  _T_18065_31 <= _T_10366_12;
                                end else begin
                                  if (_T_13104) begin
                                    _T_18065_31 <= _T_10366_13;
                                  end else begin
                                    if (_T_13102) begin
                                      _T_18065_31 <= _T_10366_14;
                                    end else begin
                                      if (_T_13100) begin
                                        _T_18065_31 <= _T_10366_15;
                                      end else begin
                                        if (_T_13098) begin
                                          _T_18065_31 <= _T_10366_16;
                                        end else begin
                                          if (_T_13096) begin
                                            _T_18065_31 <= _T_10366_17;
                                          end else begin
                                            if (_T_13094) begin
                                              _T_18065_31 <= _T_10366_18;
                                            end else begin
                                              if (_T_13092) begin
                                                _T_18065_31 <= _T_10366_19;
                                              end else begin
                                                if (_T_13090) begin
                                                  _T_18065_31 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13088) begin
                                                    _T_18065_31 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13086) begin
                                                      _T_18065_31 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13084) begin
                                                        _T_18065_31 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13082) begin
                                                          _T_18065_31 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13080) begin
                                                            _T_18065_31 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13078) begin
                                                              _T_18065_31 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13076) begin
                                                                _T_18065_31 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13074) begin
                                                                  _T_18065_31 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13072) begin
                                                                    _T_18065_31 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13070) begin
                                                                      _T_18065_31 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13068) begin
                                                                        _T_18065_31 <= _T_10366_31;
                                                                      end else begin
                                                                        _T_18065_31 <= 8'h0;
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_31 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_32) begin
        if (_T_13230) begin
          _T_18065_32 <= _T_10366_0;
        end else begin
          if (_T_13228) begin
            _T_18065_32 <= _T_10366_1;
          end else begin
            if (_T_13226) begin
              _T_18065_32 <= _T_10366_2;
            end else begin
              if (_T_13224) begin
                _T_18065_32 <= _T_10366_3;
              end else begin
                if (_T_13222) begin
                  _T_18065_32 <= _T_10366_4;
                end else begin
                  if (_T_13220) begin
                    _T_18065_32 <= _T_10366_5;
                  end else begin
                    if (_T_13218) begin
                      _T_18065_32 <= _T_10366_6;
                    end else begin
                      if (_T_13216) begin
                        _T_18065_32 <= _T_10366_7;
                      end else begin
                        if (_T_13214) begin
                          _T_18065_32 <= _T_10366_8;
                        end else begin
                          if (_T_13212) begin
                            _T_18065_32 <= _T_10366_9;
                          end else begin
                            if (_T_13210) begin
                              _T_18065_32 <= _T_10366_10;
                            end else begin
                              if (_T_13208) begin
                                _T_18065_32 <= _T_10366_11;
                              end else begin
                                if (_T_13206) begin
                                  _T_18065_32 <= _T_10366_12;
                                end else begin
                                  if (_T_13204) begin
                                    _T_18065_32 <= _T_10366_13;
                                  end else begin
                                    if (_T_13202) begin
                                      _T_18065_32 <= _T_10366_14;
                                    end else begin
                                      if (_T_13200) begin
                                        _T_18065_32 <= _T_10366_15;
                                      end else begin
                                        if (_T_13198) begin
                                          _T_18065_32 <= _T_10366_16;
                                        end else begin
                                          if (_T_13196) begin
                                            _T_18065_32 <= _T_10366_17;
                                          end else begin
                                            if (_T_13194) begin
                                              _T_18065_32 <= _T_10366_18;
                                            end else begin
                                              if (_T_13192) begin
                                                _T_18065_32 <= _T_10366_19;
                                              end else begin
                                                if (_T_13190) begin
                                                  _T_18065_32 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13188) begin
                                                    _T_18065_32 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13186) begin
                                                      _T_18065_32 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13184) begin
                                                        _T_18065_32 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13182) begin
                                                          _T_18065_32 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13180) begin
                                                            _T_18065_32 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13178) begin
                                                              _T_18065_32 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13176) begin
                                                                _T_18065_32 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13174) begin
                                                                  _T_18065_32 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13172) begin
                                                                    _T_18065_32 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13170) begin
                                                                      _T_18065_32 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13168) begin
                                                                        _T_18065_32 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13166) begin
                                                                          _T_18065_32 <= _T_10366_32;
                                                                        end else begin
                                                                          _T_18065_32 <= 8'h0;
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_32 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_33) begin
        if (_T_13333) begin
          _T_18065_33 <= _T_10366_0;
        end else begin
          if (_T_13331) begin
            _T_18065_33 <= _T_10366_1;
          end else begin
            if (_T_13329) begin
              _T_18065_33 <= _T_10366_2;
            end else begin
              if (_T_13327) begin
                _T_18065_33 <= _T_10366_3;
              end else begin
                if (_T_13325) begin
                  _T_18065_33 <= _T_10366_4;
                end else begin
                  if (_T_13323) begin
                    _T_18065_33 <= _T_10366_5;
                  end else begin
                    if (_T_13321) begin
                      _T_18065_33 <= _T_10366_6;
                    end else begin
                      if (_T_13319) begin
                        _T_18065_33 <= _T_10366_7;
                      end else begin
                        if (_T_13317) begin
                          _T_18065_33 <= _T_10366_8;
                        end else begin
                          if (_T_13315) begin
                            _T_18065_33 <= _T_10366_9;
                          end else begin
                            if (_T_13313) begin
                              _T_18065_33 <= _T_10366_10;
                            end else begin
                              if (_T_13311) begin
                                _T_18065_33 <= _T_10366_11;
                              end else begin
                                if (_T_13309) begin
                                  _T_18065_33 <= _T_10366_12;
                                end else begin
                                  if (_T_13307) begin
                                    _T_18065_33 <= _T_10366_13;
                                  end else begin
                                    if (_T_13305) begin
                                      _T_18065_33 <= _T_10366_14;
                                    end else begin
                                      if (_T_13303) begin
                                        _T_18065_33 <= _T_10366_15;
                                      end else begin
                                        if (_T_13301) begin
                                          _T_18065_33 <= _T_10366_16;
                                        end else begin
                                          if (_T_13299) begin
                                            _T_18065_33 <= _T_10366_17;
                                          end else begin
                                            if (_T_13297) begin
                                              _T_18065_33 <= _T_10366_18;
                                            end else begin
                                              if (_T_13295) begin
                                                _T_18065_33 <= _T_10366_19;
                                              end else begin
                                                if (_T_13293) begin
                                                  _T_18065_33 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13291) begin
                                                    _T_18065_33 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13289) begin
                                                      _T_18065_33 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13287) begin
                                                        _T_18065_33 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13285) begin
                                                          _T_18065_33 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13283) begin
                                                            _T_18065_33 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13281) begin
                                                              _T_18065_33 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13279) begin
                                                                _T_18065_33 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13277) begin
                                                                  _T_18065_33 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13275) begin
                                                                    _T_18065_33 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13273) begin
                                                                      _T_18065_33 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13271) begin
                                                                        _T_18065_33 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13269) begin
                                                                          _T_18065_33 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13267) begin
                                                                            _T_18065_33 <= _T_10366_33;
                                                                          end else begin
                                                                            _T_18065_33 <= 8'h0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_33 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_34) begin
        if (_T_13439) begin
          _T_18065_34 <= _T_10366_0;
        end else begin
          if (_T_13437) begin
            _T_18065_34 <= _T_10366_1;
          end else begin
            if (_T_13435) begin
              _T_18065_34 <= _T_10366_2;
            end else begin
              if (_T_13433) begin
                _T_18065_34 <= _T_10366_3;
              end else begin
                if (_T_13431) begin
                  _T_18065_34 <= _T_10366_4;
                end else begin
                  if (_T_13429) begin
                    _T_18065_34 <= _T_10366_5;
                  end else begin
                    if (_T_13427) begin
                      _T_18065_34 <= _T_10366_6;
                    end else begin
                      if (_T_13425) begin
                        _T_18065_34 <= _T_10366_7;
                      end else begin
                        if (_T_13423) begin
                          _T_18065_34 <= _T_10366_8;
                        end else begin
                          if (_T_13421) begin
                            _T_18065_34 <= _T_10366_9;
                          end else begin
                            if (_T_13419) begin
                              _T_18065_34 <= _T_10366_10;
                            end else begin
                              if (_T_13417) begin
                                _T_18065_34 <= _T_10366_11;
                              end else begin
                                if (_T_13415) begin
                                  _T_18065_34 <= _T_10366_12;
                                end else begin
                                  if (_T_13413) begin
                                    _T_18065_34 <= _T_10366_13;
                                  end else begin
                                    if (_T_13411) begin
                                      _T_18065_34 <= _T_10366_14;
                                    end else begin
                                      if (_T_13409) begin
                                        _T_18065_34 <= _T_10366_15;
                                      end else begin
                                        if (_T_13407) begin
                                          _T_18065_34 <= _T_10366_16;
                                        end else begin
                                          if (_T_13405) begin
                                            _T_18065_34 <= _T_10366_17;
                                          end else begin
                                            if (_T_13403) begin
                                              _T_18065_34 <= _T_10366_18;
                                            end else begin
                                              if (_T_13401) begin
                                                _T_18065_34 <= _T_10366_19;
                                              end else begin
                                                if (_T_13399) begin
                                                  _T_18065_34 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13397) begin
                                                    _T_18065_34 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13395) begin
                                                      _T_18065_34 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13393) begin
                                                        _T_18065_34 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13391) begin
                                                          _T_18065_34 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13389) begin
                                                            _T_18065_34 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13387) begin
                                                              _T_18065_34 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13385) begin
                                                                _T_18065_34 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13383) begin
                                                                  _T_18065_34 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13381) begin
                                                                    _T_18065_34 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13379) begin
                                                                      _T_18065_34 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13377) begin
                                                                        _T_18065_34 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13375) begin
                                                                          _T_18065_34 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13373) begin
                                                                            _T_18065_34 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13371) begin
                                                                              _T_18065_34 <= _T_10366_34;
                                                                            end else begin
                                                                              _T_18065_34 <= 8'h0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_34 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_35) begin
        if (_T_13548) begin
          _T_18065_35 <= _T_10366_0;
        end else begin
          if (_T_13546) begin
            _T_18065_35 <= _T_10366_1;
          end else begin
            if (_T_13544) begin
              _T_18065_35 <= _T_10366_2;
            end else begin
              if (_T_13542) begin
                _T_18065_35 <= _T_10366_3;
              end else begin
                if (_T_13540) begin
                  _T_18065_35 <= _T_10366_4;
                end else begin
                  if (_T_13538) begin
                    _T_18065_35 <= _T_10366_5;
                  end else begin
                    if (_T_13536) begin
                      _T_18065_35 <= _T_10366_6;
                    end else begin
                      if (_T_13534) begin
                        _T_18065_35 <= _T_10366_7;
                      end else begin
                        if (_T_13532) begin
                          _T_18065_35 <= _T_10366_8;
                        end else begin
                          if (_T_13530) begin
                            _T_18065_35 <= _T_10366_9;
                          end else begin
                            if (_T_13528) begin
                              _T_18065_35 <= _T_10366_10;
                            end else begin
                              if (_T_13526) begin
                                _T_18065_35 <= _T_10366_11;
                              end else begin
                                if (_T_13524) begin
                                  _T_18065_35 <= _T_10366_12;
                                end else begin
                                  if (_T_13522) begin
                                    _T_18065_35 <= _T_10366_13;
                                  end else begin
                                    if (_T_13520) begin
                                      _T_18065_35 <= _T_10366_14;
                                    end else begin
                                      if (_T_13518) begin
                                        _T_18065_35 <= _T_10366_15;
                                      end else begin
                                        if (_T_13516) begin
                                          _T_18065_35 <= _T_10366_16;
                                        end else begin
                                          if (_T_13514) begin
                                            _T_18065_35 <= _T_10366_17;
                                          end else begin
                                            if (_T_13512) begin
                                              _T_18065_35 <= _T_10366_18;
                                            end else begin
                                              if (_T_13510) begin
                                                _T_18065_35 <= _T_10366_19;
                                              end else begin
                                                if (_T_13508) begin
                                                  _T_18065_35 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13506) begin
                                                    _T_18065_35 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13504) begin
                                                      _T_18065_35 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13502) begin
                                                        _T_18065_35 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13500) begin
                                                          _T_18065_35 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13498) begin
                                                            _T_18065_35 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13496) begin
                                                              _T_18065_35 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13494) begin
                                                                _T_18065_35 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13492) begin
                                                                  _T_18065_35 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13490) begin
                                                                    _T_18065_35 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13488) begin
                                                                      _T_18065_35 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13486) begin
                                                                        _T_18065_35 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13484) begin
                                                                          _T_18065_35 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13482) begin
                                                                            _T_18065_35 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13480) begin
                                                                              _T_18065_35 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13478) begin
                                                                                _T_18065_35 <= _T_10366_35;
                                                                              end else begin
                                                                                _T_18065_35 <= 8'h0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_35 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_36) begin
        if (_T_13660) begin
          _T_18065_36 <= _T_10366_0;
        end else begin
          if (_T_13658) begin
            _T_18065_36 <= _T_10366_1;
          end else begin
            if (_T_13656) begin
              _T_18065_36 <= _T_10366_2;
            end else begin
              if (_T_13654) begin
                _T_18065_36 <= _T_10366_3;
              end else begin
                if (_T_13652) begin
                  _T_18065_36 <= _T_10366_4;
                end else begin
                  if (_T_13650) begin
                    _T_18065_36 <= _T_10366_5;
                  end else begin
                    if (_T_13648) begin
                      _T_18065_36 <= _T_10366_6;
                    end else begin
                      if (_T_13646) begin
                        _T_18065_36 <= _T_10366_7;
                      end else begin
                        if (_T_13644) begin
                          _T_18065_36 <= _T_10366_8;
                        end else begin
                          if (_T_13642) begin
                            _T_18065_36 <= _T_10366_9;
                          end else begin
                            if (_T_13640) begin
                              _T_18065_36 <= _T_10366_10;
                            end else begin
                              if (_T_13638) begin
                                _T_18065_36 <= _T_10366_11;
                              end else begin
                                if (_T_13636) begin
                                  _T_18065_36 <= _T_10366_12;
                                end else begin
                                  if (_T_13634) begin
                                    _T_18065_36 <= _T_10366_13;
                                  end else begin
                                    if (_T_13632) begin
                                      _T_18065_36 <= _T_10366_14;
                                    end else begin
                                      if (_T_13630) begin
                                        _T_18065_36 <= _T_10366_15;
                                      end else begin
                                        if (_T_13628) begin
                                          _T_18065_36 <= _T_10366_16;
                                        end else begin
                                          if (_T_13626) begin
                                            _T_18065_36 <= _T_10366_17;
                                          end else begin
                                            if (_T_13624) begin
                                              _T_18065_36 <= _T_10366_18;
                                            end else begin
                                              if (_T_13622) begin
                                                _T_18065_36 <= _T_10366_19;
                                              end else begin
                                                if (_T_13620) begin
                                                  _T_18065_36 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13618) begin
                                                    _T_18065_36 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13616) begin
                                                      _T_18065_36 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13614) begin
                                                        _T_18065_36 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13612) begin
                                                          _T_18065_36 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13610) begin
                                                            _T_18065_36 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13608) begin
                                                              _T_18065_36 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13606) begin
                                                                _T_18065_36 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13604) begin
                                                                  _T_18065_36 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13602) begin
                                                                    _T_18065_36 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13600) begin
                                                                      _T_18065_36 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13598) begin
                                                                        _T_18065_36 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13596) begin
                                                                          _T_18065_36 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13594) begin
                                                                            _T_18065_36 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13592) begin
                                                                              _T_18065_36 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13590) begin
                                                                                _T_18065_36 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13588) begin
                                                                                  _T_18065_36 <= _T_10366_36;
                                                                                end else begin
                                                                                  _T_18065_36 <= 8'h0;
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_36 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_37) begin
        if (_T_13775) begin
          _T_18065_37 <= _T_10366_0;
        end else begin
          if (_T_13773) begin
            _T_18065_37 <= _T_10366_1;
          end else begin
            if (_T_13771) begin
              _T_18065_37 <= _T_10366_2;
            end else begin
              if (_T_13769) begin
                _T_18065_37 <= _T_10366_3;
              end else begin
                if (_T_13767) begin
                  _T_18065_37 <= _T_10366_4;
                end else begin
                  if (_T_13765) begin
                    _T_18065_37 <= _T_10366_5;
                  end else begin
                    if (_T_13763) begin
                      _T_18065_37 <= _T_10366_6;
                    end else begin
                      if (_T_13761) begin
                        _T_18065_37 <= _T_10366_7;
                      end else begin
                        if (_T_13759) begin
                          _T_18065_37 <= _T_10366_8;
                        end else begin
                          if (_T_13757) begin
                            _T_18065_37 <= _T_10366_9;
                          end else begin
                            if (_T_13755) begin
                              _T_18065_37 <= _T_10366_10;
                            end else begin
                              if (_T_13753) begin
                                _T_18065_37 <= _T_10366_11;
                              end else begin
                                if (_T_13751) begin
                                  _T_18065_37 <= _T_10366_12;
                                end else begin
                                  if (_T_13749) begin
                                    _T_18065_37 <= _T_10366_13;
                                  end else begin
                                    if (_T_13747) begin
                                      _T_18065_37 <= _T_10366_14;
                                    end else begin
                                      if (_T_13745) begin
                                        _T_18065_37 <= _T_10366_15;
                                      end else begin
                                        if (_T_13743) begin
                                          _T_18065_37 <= _T_10366_16;
                                        end else begin
                                          if (_T_13741) begin
                                            _T_18065_37 <= _T_10366_17;
                                          end else begin
                                            if (_T_13739) begin
                                              _T_18065_37 <= _T_10366_18;
                                            end else begin
                                              if (_T_13737) begin
                                                _T_18065_37 <= _T_10366_19;
                                              end else begin
                                                if (_T_13735) begin
                                                  _T_18065_37 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13733) begin
                                                    _T_18065_37 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13731) begin
                                                      _T_18065_37 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13729) begin
                                                        _T_18065_37 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13727) begin
                                                          _T_18065_37 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13725) begin
                                                            _T_18065_37 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13723) begin
                                                              _T_18065_37 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13721) begin
                                                                _T_18065_37 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13719) begin
                                                                  _T_18065_37 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13717) begin
                                                                    _T_18065_37 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13715) begin
                                                                      _T_18065_37 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13713) begin
                                                                        _T_18065_37 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13711) begin
                                                                          _T_18065_37 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13709) begin
                                                                            _T_18065_37 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13707) begin
                                                                              _T_18065_37 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13705) begin
                                                                                _T_18065_37 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13703) begin
                                                                                  _T_18065_37 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13701) begin
                                                                                    _T_18065_37 <= _T_10366_37;
                                                                                  end else begin
                                                                                    _T_18065_37 <= 8'h0;
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_37 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_38) begin
        if (_T_13893) begin
          _T_18065_38 <= _T_10366_0;
        end else begin
          if (_T_13891) begin
            _T_18065_38 <= _T_10366_1;
          end else begin
            if (_T_13889) begin
              _T_18065_38 <= _T_10366_2;
            end else begin
              if (_T_13887) begin
                _T_18065_38 <= _T_10366_3;
              end else begin
                if (_T_13885) begin
                  _T_18065_38 <= _T_10366_4;
                end else begin
                  if (_T_13883) begin
                    _T_18065_38 <= _T_10366_5;
                  end else begin
                    if (_T_13881) begin
                      _T_18065_38 <= _T_10366_6;
                    end else begin
                      if (_T_13879) begin
                        _T_18065_38 <= _T_10366_7;
                      end else begin
                        if (_T_13877) begin
                          _T_18065_38 <= _T_10366_8;
                        end else begin
                          if (_T_13875) begin
                            _T_18065_38 <= _T_10366_9;
                          end else begin
                            if (_T_13873) begin
                              _T_18065_38 <= _T_10366_10;
                            end else begin
                              if (_T_13871) begin
                                _T_18065_38 <= _T_10366_11;
                              end else begin
                                if (_T_13869) begin
                                  _T_18065_38 <= _T_10366_12;
                                end else begin
                                  if (_T_13867) begin
                                    _T_18065_38 <= _T_10366_13;
                                  end else begin
                                    if (_T_13865) begin
                                      _T_18065_38 <= _T_10366_14;
                                    end else begin
                                      if (_T_13863) begin
                                        _T_18065_38 <= _T_10366_15;
                                      end else begin
                                        if (_T_13861) begin
                                          _T_18065_38 <= _T_10366_16;
                                        end else begin
                                          if (_T_13859) begin
                                            _T_18065_38 <= _T_10366_17;
                                          end else begin
                                            if (_T_13857) begin
                                              _T_18065_38 <= _T_10366_18;
                                            end else begin
                                              if (_T_13855) begin
                                                _T_18065_38 <= _T_10366_19;
                                              end else begin
                                                if (_T_13853) begin
                                                  _T_18065_38 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13851) begin
                                                    _T_18065_38 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13849) begin
                                                      _T_18065_38 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13847) begin
                                                        _T_18065_38 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13845) begin
                                                          _T_18065_38 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13843) begin
                                                            _T_18065_38 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13841) begin
                                                              _T_18065_38 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13839) begin
                                                                _T_18065_38 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13837) begin
                                                                  _T_18065_38 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13835) begin
                                                                    _T_18065_38 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13833) begin
                                                                      _T_18065_38 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13831) begin
                                                                        _T_18065_38 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13829) begin
                                                                          _T_18065_38 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13827) begin
                                                                            _T_18065_38 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13825) begin
                                                                              _T_18065_38 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13823) begin
                                                                                _T_18065_38 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13821) begin
                                                                                  _T_18065_38 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13819) begin
                                                                                    _T_18065_38 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_13817) begin
                                                                                      _T_18065_38 <= _T_10366_38;
                                                                                    end else begin
                                                                                      _T_18065_38 <= 8'h0;
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_38 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_39) begin
        if (_T_14014) begin
          _T_18065_39 <= _T_10366_0;
        end else begin
          if (_T_14012) begin
            _T_18065_39 <= _T_10366_1;
          end else begin
            if (_T_14010) begin
              _T_18065_39 <= _T_10366_2;
            end else begin
              if (_T_14008) begin
                _T_18065_39 <= _T_10366_3;
              end else begin
                if (_T_14006) begin
                  _T_18065_39 <= _T_10366_4;
                end else begin
                  if (_T_14004) begin
                    _T_18065_39 <= _T_10366_5;
                  end else begin
                    if (_T_14002) begin
                      _T_18065_39 <= _T_10366_6;
                    end else begin
                      if (_T_14000) begin
                        _T_18065_39 <= _T_10366_7;
                      end else begin
                        if (_T_13998) begin
                          _T_18065_39 <= _T_10366_8;
                        end else begin
                          if (_T_13996) begin
                            _T_18065_39 <= _T_10366_9;
                          end else begin
                            if (_T_13994) begin
                              _T_18065_39 <= _T_10366_10;
                            end else begin
                              if (_T_13992) begin
                                _T_18065_39 <= _T_10366_11;
                              end else begin
                                if (_T_13990) begin
                                  _T_18065_39 <= _T_10366_12;
                                end else begin
                                  if (_T_13988) begin
                                    _T_18065_39 <= _T_10366_13;
                                  end else begin
                                    if (_T_13986) begin
                                      _T_18065_39 <= _T_10366_14;
                                    end else begin
                                      if (_T_13984) begin
                                        _T_18065_39 <= _T_10366_15;
                                      end else begin
                                        if (_T_13982) begin
                                          _T_18065_39 <= _T_10366_16;
                                        end else begin
                                          if (_T_13980) begin
                                            _T_18065_39 <= _T_10366_17;
                                          end else begin
                                            if (_T_13978) begin
                                              _T_18065_39 <= _T_10366_18;
                                            end else begin
                                              if (_T_13976) begin
                                                _T_18065_39 <= _T_10366_19;
                                              end else begin
                                                if (_T_13974) begin
                                                  _T_18065_39 <= _T_10366_20;
                                                end else begin
                                                  if (_T_13972) begin
                                                    _T_18065_39 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_13970) begin
                                                      _T_18065_39 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_13968) begin
                                                        _T_18065_39 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_13966) begin
                                                          _T_18065_39 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_13964) begin
                                                            _T_18065_39 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_13962) begin
                                                              _T_18065_39 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_13960) begin
                                                                _T_18065_39 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_13958) begin
                                                                  _T_18065_39 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_13956) begin
                                                                    _T_18065_39 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_13954) begin
                                                                      _T_18065_39 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_13952) begin
                                                                        _T_18065_39 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_13950) begin
                                                                          _T_18065_39 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_13948) begin
                                                                            _T_18065_39 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_13946) begin
                                                                              _T_18065_39 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_13944) begin
                                                                                _T_18065_39 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_13942) begin
                                                                                  _T_18065_39 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_13940) begin
                                                                                    _T_18065_39 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_13938) begin
                                                                                      _T_18065_39 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_13936) begin
                                                                                        _T_18065_39 <= _T_10366_39;
                                                                                      end else begin
                                                                                        _T_18065_39 <= 8'h0;
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_39 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_40) begin
        if (_T_14138) begin
          _T_18065_40 <= _T_10366_0;
        end else begin
          if (_T_14136) begin
            _T_18065_40 <= _T_10366_1;
          end else begin
            if (_T_14134) begin
              _T_18065_40 <= _T_10366_2;
            end else begin
              if (_T_14132) begin
                _T_18065_40 <= _T_10366_3;
              end else begin
                if (_T_14130) begin
                  _T_18065_40 <= _T_10366_4;
                end else begin
                  if (_T_14128) begin
                    _T_18065_40 <= _T_10366_5;
                  end else begin
                    if (_T_14126) begin
                      _T_18065_40 <= _T_10366_6;
                    end else begin
                      if (_T_14124) begin
                        _T_18065_40 <= _T_10366_7;
                      end else begin
                        if (_T_14122) begin
                          _T_18065_40 <= _T_10366_8;
                        end else begin
                          if (_T_14120) begin
                            _T_18065_40 <= _T_10366_9;
                          end else begin
                            if (_T_14118) begin
                              _T_18065_40 <= _T_10366_10;
                            end else begin
                              if (_T_14116) begin
                                _T_18065_40 <= _T_10366_11;
                              end else begin
                                if (_T_14114) begin
                                  _T_18065_40 <= _T_10366_12;
                                end else begin
                                  if (_T_14112) begin
                                    _T_18065_40 <= _T_10366_13;
                                  end else begin
                                    if (_T_14110) begin
                                      _T_18065_40 <= _T_10366_14;
                                    end else begin
                                      if (_T_14108) begin
                                        _T_18065_40 <= _T_10366_15;
                                      end else begin
                                        if (_T_14106) begin
                                          _T_18065_40 <= _T_10366_16;
                                        end else begin
                                          if (_T_14104) begin
                                            _T_18065_40 <= _T_10366_17;
                                          end else begin
                                            if (_T_14102) begin
                                              _T_18065_40 <= _T_10366_18;
                                            end else begin
                                              if (_T_14100) begin
                                                _T_18065_40 <= _T_10366_19;
                                              end else begin
                                                if (_T_14098) begin
                                                  _T_18065_40 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14096) begin
                                                    _T_18065_40 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14094) begin
                                                      _T_18065_40 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14092) begin
                                                        _T_18065_40 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14090) begin
                                                          _T_18065_40 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14088) begin
                                                            _T_18065_40 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14086) begin
                                                              _T_18065_40 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14084) begin
                                                                _T_18065_40 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14082) begin
                                                                  _T_18065_40 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14080) begin
                                                                    _T_18065_40 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14078) begin
                                                                      _T_18065_40 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14076) begin
                                                                        _T_18065_40 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14074) begin
                                                                          _T_18065_40 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14072) begin
                                                                            _T_18065_40 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14070) begin
                                                                              _T_18065_40 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14068) begin
                                                                                _T_18065_40 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14066) begin
                                                                                  _T_18065_40 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14064) begin
                                                                                    _T_18065_40 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14062) begin
                                                                                      _T_18065_40 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14060) begin
                                                                                        _T_18065_40 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14058) begin
                                                                                          _T_18065_40 <= _T_10366_40;
                                                                                        end else begin
                                                                                          _T_18065_40 <= 8'h0;
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_40 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_41) begin
        if (_T_14265) begin
          _T_18065_41 <= _T_10366_0;
        end else begin
          if (_T_14263) begin
            _T_18065_41 <= _T_10366_1;
          end else begin
            if (_T_14261) begin
              _T_18065_41 <= _T_10366_2;
            end else begin
              if (_T_14259) begin
                _T_18065_41 <= _T_10366_3;
              end else begin
                if (_T_14257) begin
                  _T_18065_41 <= _T_10366_4;
                end else begin
                  if (_T_14255) begin
                    _T_18065_41 <= _T_10366_5;
                  end else begin
                    if (_T_14253) begin
                      _T_18065_41 <= _T_10366_6;
                    end else begin
                      if (_T_14251) begin
                        _T_18065_41 <= _T_10366_7;
                      end else begin
                        if (_T_14249) begin
                          _T_18065_41 <= _T_10366_8;
                        end else begin
                          if (_T_14247) begin
                            _T_18065_41 <= _T_10366_9;
                          end else begin
                            if (_T_14245) begin
                              _T_18065_41 <= _T_10366_10;
                            end else begin
                              if (_T_14243) begin
                                _T_18065_41 <= _T_10366_11;
                              end else begin
                                if (_T_14241) begin
                                  _T_18065_41 <= _T_10366_12;
                                end else begin
                                  if (_T_14239) begin
                                    _T_18065_41 <= _T_10366_13;
                                  end else begin
                                    if (_T_14237) begin
                                      _T_18065_41 <= _T_10366_14;
                                    end else begin
                                      if (_T_14235) begin
                                        _T_18065_41 <= _T_10366_15;
                                      end else begin
                                        if (_T_14233) begin
                                          _T_18065_41 <= _T_10366_16;
                                        end else begin
                                          if (_T_14231) begin
                                            _T_18065_41 <= _T_10366_17;
                                          end else begin
                                            if (_T_14229) begin
                                              _T_18065_41 <= _T_10366_18;
                                            end else begin
                                              if (_T_14227) begin
                                                _T_18065_41 <= _T_10366_19;
                                              end else begin
                                                if (_T_14225) begin
                                                  _T_18065_41 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14223) begin
                                                    _T_18065_41 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14221) begin
                                                      _T_18065_41 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14219) begin
                                                        _T_18065_41 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14217) begin
                                                          _T_18065_41 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14215) begin
                                                            _T_18065_41 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14213) begin
                                                              _T_18065_41 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14211) begin
                                                                _T_18065_41 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14209) begin
                                                                  _T_18065_41 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14207) begin
                                                                    _T_18065_41 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14205) begin
                                                                      _T_18065_41 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14203) begin
                                                                        _T_18065_41 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14201) begin
                                                                          _T_18065_41 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14199) begin
                                                                            _T_18065_41 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14197) begin
                                                                              _T_18065_41 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14195) begin
                                                                                _T_18065_41 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14193) begin
                                                                                  _T_18065_41 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14191) begin
                                                                                    _T_18065_41 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14189) begin
                                                                                      _T_18065_41 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14187) begin
                                                                                        _T_18065_41 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14185) begin
                                                                                          _T_18065_41 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14183) begin
                                                                                            _T_18065_41 <= _T_10366_41;
                                                                                          end else begin
                                                                                            _T_18065_41 <= 8'h0;
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_41 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_42) begin
        if (_T_14395) begin
          _T_18065_42 <= _T_10366_0;
        end else begin
          if (_T_14393) begin
            _T_18065_42 <= _T_10366_1;
          end else begin
            if (_T_14391) begin
              _T_18065_42 <= _T_10366_2;
            end else begin
              if (_T_14389) begin
                _T_18065_42 <= _T_10366_3;
              end else begin
                if (_T_14387) begin
                  _T_18065_42 <= _T_10366_4;
                end else begin
                  if (_T_14385) begin
                    _T_18065_42 <= _T_10366_5;
                  end else begin
                    if (_T_14383) begin
                      _T_18065_42 <= _T_10366_6;
                    end else begin
                      if (_T_14381) begin
                        _T_18065_42 <= _T_10366_7;
                      end else begin
                        if (_T_14379) begin
                          _T_18065_42 <= _T_10366_8;
                        end else begin
                          if (_T_14377) begin
                            _T_18065_42 <= _T_10366_9;
                          end else begin
                            if (_T_14375) begin
                              _T_18065_42 <= _T_10366_10;
                            end else begin
                              if (_T_14373) begin
                                _T_18065_42 <= _T_10366_11;
                              end else begin
                                if (_T_14371) begin
                                  _T_18065_42 <= _T_10366_12;
                                end else begin
                                  if (_T_14369) begin
                                    _T_18065_42 <= _T_10366_13;
                                  end else begin
                                    if (_T_14367) begin
                                      _T_18065_42 <= _T_10366_14;
                                    end else begin
                                      if (_T_14365) begin
                                        _T_18065_42 <= _T_10366_15;
                                      end else begin
                                        if (_T_14363) begin
                                          _T_18065_42 <= _T_10366_16;
                                        end else begin
                                          if (_T_14361) begin
                                            _T_18065_42 <= _T_10366_17;
                                          end else begin
                                            if (_T_14359) begin
                                              _T_18065_42 <= _T_10366_18;
                                            end else begin
                                              if (_T_14357) begin
                                                _T_18065_42 <= _T_10366_19;
                                              end else begin
                                                if (_T_14355) begin
                                                  _T_18065_42 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14353) begin
                                                    _T_18065_42 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14351) begin
                                                      _T_18065_42 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14349) begin
                                                        _T_18065_42 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14347) begin
                                                          _T_18065_42 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14345) begin
                                                            _T_18065_42 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14343) begin
                                                              _T_18065_42 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14341) begin
                                                                _T_18065_42 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14339) begin
                                                                  _T_18065_42 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14337) begin
                                                                    _T_18065_42 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14335) begin
                                                                      _T_18065_42 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14333) begin
                                                                        _T_18065_42 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14331) begin
                                                                          _T_18065_42 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14329) begin
                                                                            _T_18065_42 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14327) begin
                                                                              _T_18065_42 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14325) begin
                                                                                _T_18065_42 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14323) begin
                                                                                  _T_18065_42 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14321) begin
                                                                                    _T_18065_42 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14319) begin
                                                                                      _T_18065_42 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14317) begin
                                                                                        _T_18065_42 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14315) begin
                                                                                          _T_18065_42 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14313) begin
                                                                                            _T_18065_42 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14311) begin
                                                                                              _T_18065_42 <= _T_10366_42;
                                                                                            end else begin
                                                                                              _T_18065_42 <= 8'h0;
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_42 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_43) begin
        if (_T_14528) begin
          _T_18065_43 <= _T_10366_0;
        end else begin
          if (_T_14526) begin
            _T_18065_43 <= _T_10366_1;
          end else begin
            if (_T_14524) begin
              _T_18065_43 <= _T_10366_2;
            end else begin
              if (_T_14522) begin
                _T_18065_43 <= _T_10366_3;
              end else begin
                if (_T_14520) begin
                  _T_18065_43 <= _T_10366_4;
                end else begin
                  if (_T_14518) begin
                    _T_18065_43 <= _T_10366_5;
                  end else begin
                    if (_T_14516) begin
                      _T_18065_43 <= _T_10366_6;
                    end else begin
                      if (_T_14514) begin
                        _T_18065_43 <= _T_10366_7;
                      end else begin
                        if (_T_14512) begin
                          _T_18065_43 <= _T_10366_8;
                        end else begin
                          if (_T_14510) begin
                            _T_18065_43 <= _T_10366_9;
                          end else begin
                            if (_T_14508) begin
                              _T_18065_43 <= _T_10366_10;
                            end else begin
                              if (_T_14506) begin
                                _T_18065_43 <= _T_10366_11;
                              end else begin
                                if (_T_14504) begin
                                  _T_18065_43 <= _T_10366_12;
                                end else begin
                                  if (_T_14502) begin
                                    _T_18065_43 <= _T_10366_13;
                                  end else begin
                                    if (_T_14500) begin
                                      _T_18065_43 <= _T_10366_14;
                                    end else begin
                                      if (_T_14498) begin
                                        _T_18065_43 <= _T_10366_15;
                                      end else begin
                                        if (_T_14496) begin
                                          _T_18065_43 <= _T_10366_16;
                                        end else begin
                                          if (_T_14494) begin
                                            _T_18065_43 <= _T_10366_17;
                                          end else begin
                                            if (_T_14492) begin
                                              _T_18065_43 <= _T_10366_18;
                                            end else begin
                                              if (_T_14490) begin
                                                _T_18065_43 <= _T_10366_19;
                                              end else begin
                                                if (_T_14488) begin
                                                  _T_18065_43 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14486) begin
                                                    _T_18065_43 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14484) begin
                                                      _T_18065_43 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14482) begin
                                                        _T_18065_43 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14480) begin
                                                          _T_18065_43 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14478) begin
                                                            _T_18065_43 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14476) begin
                                                              _T_18065_43 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14474) begin
                                                                _T_18065_43 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14472) begin
                                                                  _T_18065_43 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14470) begin
                                                                    _T_18065_43 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14468) begin
                                                                      _T_18065_43 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14466) begin
                                                                        _T_18065_43 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14464) begin
                                                                          _T_18065_43 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14462) begin
                                                                            _T_18065_43 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14460) begin
                                                                              _T_18065_43 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14458) begin
                                                                                _T_18065_43 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14456) begin
                                                                                  _T_18065_43 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14454) begin
                                                                                    _T_18065_43 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14452) begin
                                                                                      _T_18065_43 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14450) begin
                                                                                        _T_18065_43 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14448) begin
                                                                                          _T_18065_43 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14446) begin
                                                                                            _T_18065_43 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14444) begin
                                                                                              _T_18065_43 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14442) begin
                                                                                                _T_18065_43 <= _T_10366_43;
                                                                                              end else begin
                                                                                                _T_18065_43 <= 8'h0;
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_43 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_44) begin
        if (_T_14664) begin
          _T_18065_44 <= _T_10366_0;
        end else begin
          if (_T_14662) begin
            _T_18065_44 <= _T_10366_1;
          end else begin
            if (_T_14660) begin
              _T_18065_44 <= _T_10366_2;
            end else begin
              if (_T_14658) begin
                _T_18065_44 <= _T_10366_3;
              end else begin
                if (_T_14656) begin
                  _T_18065_44 <= _T_10366_4;
                end else begin
                  if (_T_14654) begin
                    _T_18065_44 <= _T_10366_5;
                  end else begin
                    if (_T_14652) begin
                      _T_18065_44 <= _T_10366_6;
                    end else begin
                      if (_T_14650) begin
                        _T_18065_44 <= _T_10366_7;
                      end else begin
                        if (_T_14648) begin
                          _T_18065_44 <= _T_10366_8;
                        end else begin
                          if (_T_14646) begin
                            _T_18065_44 <= _T_10366_9;
                          end else begin
                            if (_T_14644) begin
                              _T_18065_44 <= _T_10366_10;
                            end else begin
                              if (_T_14642) begin
                                _T_18065_44 <= _T_10366_11;
                              end else begin
                                if (_T_14640) begin
                                  _T_18065_44 <= _T_10366_12;
                                end else begin
                                  if (_T_14638) begin
                                    _T_18065_44 <= _T_10366_13;
                                  end else begin
                                    if (_T_14636) begin
                                      _T_18065_44 <= _T_10366_14;
                                    end else begin
                                      if (_T_14634) begin
                                        _T_18065_44 <= _T_10366_15;
                                      end else begin
                                        if (_T_14632) begin
                                          _T_18065_44 <= _T_10366_16;
                                        end else begin
                                          if (_T_14630) begin
                                            _T_18065_44 <= _T_10366_17;
                                          end else begin
                                            if (_T_14628) begin
                                              _T_18065_44 <= _T_10366_18;
                                            end else begin
                                              if (_T_14626) begin
                                                _T_18065_44 <= _T_10366_19;
                                              end else begin
                                                if (_T_14624) begin
                                                  _T_18065_44 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14622) begin
                                                    _T_18065_44 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14620) begin
                                                      _T_18065_44 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14618) begin
                                                        _T_18065_44 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14616) begin
                                                          _T_18065_44 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14614) begin
                                                            _T_18065_44 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14612) begin
                                                              _T_18065_44 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14610) begin
                                                                _T_18065_44 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14608) begin
                                                                  _T_18065_44 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14606) begin
                                                                    _T_18065_44 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14604) begin
                                                                      _T_18065_44 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14602) begin
                                                                        _T_18065_44 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14600) begin
                                                                          _T_18065_44 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14598) begin
                                                                            _T_18065_44 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14596) begin
                                                                              _T_18065_44 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14594) begin
                                                                                _T_18065_44 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14592) begin
                                                                                  _T_18065_44 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14590) begin
                                                                                    _T_18065_44 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14588) begin
                                                                                      _T_18065_44 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14586) begin
                                                                                        _T_18065_44 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14584) begin
                                                                                          _T_18065_44 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14582) begin
                                                                                            _T_18065_44 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14580) begin
                                                                                              _T_18065_44 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14578) begin
                                                                                                _T_18065_44 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14576) begin
                                                                                                  _T_18065_44 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  _T_18065_44 <= 8'h0;
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_44 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_45) begin
        if (_T_14803) begin
          _T_18065_45 <= _T_10366_0;
        end else begin
          if (_T_14801) begin
            _T_18065_45 <= _T_10366_1;
          end else begin
            if (_T_14799) begin
              _T_18065_45 <= _T_10366_2;
            end else begin
              if (_T_14797) begin
                _T_18065_45 <= _T_10366_3;
              end else begin
                if (_T_14795) begin
                  _T_18065_45 <= _T_10366_4;
                end else begin
                  if (_T_14793) begin
                    _T_18065_45 <= _T_10366_5;
                  end else begin
                    if (_T_14791) begin
                      _T_18065_45 <= _T_10366_6;
                    end else begin
                      if (_T_14789) begin
                        _T_18065_45 <= _T_10366_7;
                      end else begin
                        if (_T_14787) begin
                          _T_18065_45 <= _T_10366_8;
                        end else begin
                          if (_T_14785) begin
                            _T_18065_45 <= _T_10366_9;
                          end else begin
                            if (_T_14783) begin
                              _T_18065_45 <= _T_10366_10;
                            end else begin
                              if (_T_14781) begin
                                _T_18065_45 <= _T_10366_11;
                              end else begin
                                if (_T_14779) begin
                                  _T_18065_45 <= _T_10366_12;
                                end else begin
                                  if (_T_14777) begin
                                    _T_18065_45 <= _T_10366_13;
                                  end else begin
                                    if (_T_14775) begin
                                      _T_18065_45 <= _T_10366_14;
                                    end else begin
                                      if (_T_14773) begin
                                        _T_18065_45 <= _T_10366_15;
                                      end else begin
                                        if (_T_14771) begin
                                          _T_18065_45 <= _T_10366_16;
                                        end else begin
                                          if (_T_14769) begin
                                            _T_18065_45 <= _T_10366_17;
                                          end else begin
                                            if (_T_14767) begin
                                              _T_18065_45 <= _T_10366_18;
                                            end else begin
                                              if (_T_14765) begin
                                                _T_18065_45 <= _T_10366_19;
                                              end else begin
                                                if (_T_14763) begin
                                                  _T_18065_45 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14761) begin
                                                    _T_18065_45 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14759) begin
                                                      _T_18065_45 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14757) begin
                                                        _T_18065_45 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14755) begin
                                                          _T_18065_45 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14753) begin
                                                            _T_18065_45 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14751) begin
                                                              _T_18065_45 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14749) begin
                                                                _T_18065_45 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14747) begin
                                                                  _T_18065_45 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14745) begin
                                                                    _T_18065_45 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14743) begin
                                                                      _T_18065_45 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14741) begin
                                                                        _T_18065_45 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14739) begin
                                                                          _T_18065_45 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14737) begin
                                                                            _T_18065_45 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14735) begin
                                                                              _T_18065_45 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14733) begin
                                                                                _T_18065_45 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14731) begin
                                                                                  _T_18065_45 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14729) begin
                                                                                    _T_18065_45 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14727) begin
                                                                                      _T_18065_45 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14725) begin
                                                                                        _T_18065_45 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14723) begin
                                                                                          _T_18065_45 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14721) begin
                                                                                            _T_18065_45 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14719) begin
                                                                                              _T_18065_45 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14717) begin
                                                                                                _T_18065_45 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14715) begin
                                                                                                  _T_18065_45 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_14713) begin
                                                                                                    _T_18065_45 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    _T_18065_45 <= 8'h0;
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_45 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_46) begin
        if (_T_14945) begin
          _T_18065_46 <= _T_10366_0;
        end else begin
          if (_T_14943) begin
            _T_18065_46 <= _T_10366_1;
          end else begin
            if (_T_14941) begin
              _T_18065_46 <= _T_10366_2;
            end else begin
              if (_T_14939) begin
                _T_18065_46 <= _T_10366_3;
              end else begin
                if (_T_14937) begin
                  _T_18065_46 <= _T_10366_4;
                end else begin
                  if (_T_14935) begin
                    _T_18065_46 <= _T_10366_5;
                  end else begin
                    if (_T_14933) begin
                      _T_18065_46 <= _T_10366_6;
                    end else begin
                      if (_T_14931) begin
                        _T_18065_46 <= _T_10366_7;
                      end else begin
                        if (_T_14929) begin
                          _T_18065_46 <= _T_10366_8;
                        end else begin
                          if (_T_14927) begin
                            _T_18065_46 <= _T_10366_9;
                          end else begin
                            if (_T_14925) begin
                              _T_18065_46 <= _T_10366_10;
                            end else begin
                              if (_T_14923) begin
                                _T_18065_46 <= _T_10366_11;
                              end else begin
                                if (_T_14921) begin
                                  _T_18065_46 <= _T_10366_12;
                                end else begin
                                  if (_T_14919) begin
                                    _T_18065_46 <= _T_10366_13;
                                  end else begin
                                    if (_T_14917) begin
                                      _T_18065_46 <= _T_10366_14;
                                    end else begin
                                      if (_T_14915) begin
                                        _T_18065_46 <= _T_10366_15;
                                      end else begin
                                        if (_T_14913) begin
                                          _T_18065_46 <= _T_10366_16;
                                        end else begin
                                          if (_T_14911) begin
                                            _T_18065_46 <= _T_10366_17;
                                          end else begin
                                            if (_T_14909) begin
                                              _T_18065_46 <= _T_10366_18;
                                            end else begin
                                              if (_T_14907) begin
                                                _T_18065_46 <= _T_10366_19;
                                              end else begin
                                                if (_T_14905) begin
                                                  _T_18065_46 <= _T_10366_20;
                                                end else begin
                                                  if (_T_14903) begin
                                                    _T_18065_46 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_14901) begin
                                                      _T_18065_46 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_14899) begin
                                                        _T_18065_46 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_14897) begin
                                                          _T_18065_46 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_14895) begin
                                                            _T_18065_46 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_14893) begin
                                                              _T_18065_46 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_14891) begin
                                                                _T_18065_46 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_14889) begin
                                                                  _T_18065_46 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_14887) begin
                                                                    _T_18065_46 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_14885) begin
                                                                      _T_18065_46 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_14883) begin
                                                                        _T_18065_46 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_14881) begin
                                                                          _T_18065_46 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_14879) begin
                                                                            _T_18065_46 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_14877) begin
                                                                              _T_18065_46 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_14875) begin
                                                                                _T_18065_46 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_14873) begin
                                                                                  _T_18065_46 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_14871) begin
                                                                                    _T_18065_46 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_14869) begin
                                                                                      _T_18065_46 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_14867) begin
                                                                                        _T_18065_46 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_14865) begin
                                                                                          _T_18065_46 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_14863) begin
                                                                                            _T_18065_46 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_14861) begin
                                                                                              _T_18065_46 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_14859) begin
                                                                                                _T_18065_46 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_14857) begin
                                                                                                  _T_18065_46 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_14855) begin
                                                                                                    _T_18065_46 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_14853) begin
                                                                                                      _T_18065_46 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      _T_18065_46 <= 8'h0;
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_46 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_47) begin
        if (_T_15090) begin
          _T_18065_47 <= _T_10366_0;
        end else begin
          if (_T_15088) begin
            _T_18065_47 <= _T_10366_1;
          end else begin
            if (_T_15086) begin
              _T_18065_47 <= _T_10366_2;
            end else begin
              if (_T_15084) begin
                _T_18065_47 <= _T_10366_3;
              end else begin
                if (_T_15082) begin
                  _T_18065_47 <= _T_10366_4;
                end else begin
                  if (_T_15080) begin
                    _T_18065_47 <= _T_10366_5;
                  end else begin
                    if (_T_15078) begin
                      _T_18065_47 <= _T_10366_6;
                    end else begin
                      if (_T_15076) begin
                        _T_18065_47 <= _T_10366_7;
                      end else begin
                        if (_T_15074) begin
                          _T_18065_47 <= _T_10366_8;
                        end else begin
                          if (_T_15072) begin
                            _T_18065_47 <= _T_10366_9;
                          end else begin
                            if (_T_15070) begin
                              _T_18065_47 <= _T_10366_10;
                            end else begin
                              if (_T_15068) begin
                                _T_18065_47 <= _T_10366_11;
                              end else begin
                                if (_T_15066) begin
                                  _T_18065_47 <= _T_10366_12;
                                end else begin
                                  if (_T_15064) begin
                                    _T_18065_47 <= _T_10366_13;
                                  end else begin
                                    if (_T_15062) begin
                                      _T_18065_47 <= _T_10366_14;
                                    end else begin
                                      if (_T_15060) begin
                                        _T_18065_47 <= _T_10366_15;
                                      end else begin
                                        if (_T_15058) begin
                                          _T_18065_47 <= _T_10366_16;
                                        end else begin
                                          if (_T_15056) begin
                                            _T_18065_47 <= _T_10366_17;
                                          end else begin
                                            if (_T_15054) begin
                                              _T_18065_47 <= _T_10366_18;
                                            end else begin
                                              if (_T_15052) begin
                                                _T_18065_47 <= _T_10366_19;
                                              end else begin
                                                if (_T_15050) begin
                                                  _T_18065_47 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15048) begin
                                                    _T_18065_47 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15046) begin
                                                      _T_18065_47 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15044) begin
                                                        _T_18065_47 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15042) begin
                                                          _T_18065_47 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15040) begin
                                                            _T_18065_47 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15038) begin
                                                              _T_18065_47 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15036) begin
                                                                _T_18065_47 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15034) begin
                                                                  _T_18065_47 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15032) begin
                                                                    _T_18065_47 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15030) begin
                                                                      _T_18065_47 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15028) begin
                                                                        _T_18065_47 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15026) begin
                                                                          _T_18065_47 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15024) begin
                                                                            _T_18065_47 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15022) begin
                                                                              _T_18065_47 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15020) begin
                                                                                _T_18065_47 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15018) begin
                                                                                  _T_18065_47 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15016) begin
                                                                                    _T_18065_47 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15014) begin
                                                                                      _T_18065_47 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15012) begin
                                                                                        _T_18065_47 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15010) begin
                                                                                          _T_18065_47 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15008) begin
                                                                                            _T_18065_47 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15006) begin
                                                                                              _T_18065_47 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15004) begin
                                                                                                _T_18065_47 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15002) begin
                                                                                                  _T_18065_47 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15000) begin
                                                                                                    _T_18065_47 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_14998) begin
                                                                                                      _T_18065_47 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_14996) begin
                                                                                                        _T_18065_47 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        _T_18065_47 <= 8'h0;
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_47 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_48) begin
        if (_T_15238) begin
          _T_18065_48 <= _T_10366_0;
        end else begin
          if (_T_15236) begin
            _T_18065_48 <= _T_10366_1;
          end else begin
            if (_T_15234) begin
              _T_18065_48 <= _T_10366_2;
            end else begin
              if (_T_15232) begin
                _T_18065_48 <= _T_10366_3;
              end else begin
                if (_T_15230) begin
                  _T_18065_48 <= _T_10366_4;
                end else begin
                  if (_T_15228) begin
                    _T_18065_48 <= _T_10366_5;
                  end else begin
                    if (_T_15226) begin
                      _T_18065_48 <= _T_10366_6;
                    end else begin
                      if (_T_15224) begin
                        _T_18065_48 <= _T_10366_7;
                      end else begin
                        if (_T_15222) begin
                          _T_18065_48 <= _T_10366_8;
                        end else begin
                          if (_T_15220) begin
                            _T_18065_48 <= _T_10366_9;
                          end else begin
                            if (_T_15218) begin
                              _T_18065_48 <= _T_10366_10;
                            end else begin
                              if (_T_15216) begin
                                _T_18065_48 <= _T_10366_11;
                              end else begin
                                if (_T_15214) begin
                                  _T_18065_48 <= _T_10366_12;
                                end else begin
                                  if (_T_15212) begin
                                    _T_18065_48 <= _T_10366_13;
                                  end else begin
                                    if (_T_15210) begin
                                      _T_18065_48 <= _T_10366_14;
                                    end else begin
                                      if (_T_15208) begin
                                        _T_18065_48 <= _T_10366_15;
                                      end else begin
                                        if (_T_15206) begin
                                          _T_18065_48 <= _T_10366_16;
                                        end else begin
                                          if (_T_15204) begin
                                            _T_18065_48 <= _T_10366_17;
                                          end else begin
                                            if (_T_15202) begin
                                              _T_18065_48 <= _T_10366_18;
                                            end else begin
                                              if (_T_15200) begin
                                                _T_18065_48 <= _T_10366_19;
                                              end else begin
                                                if (_T_15198) begin
                                                  _T_18065_48 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15196) begin
                                                    _T_18065_48 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15194) begin
                                                      _T_18065_48 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15192) begin
                                                        _T_18065_48 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15190) begin
                                                          _T_18065_48 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15188) begin
                                                            _T_18065_48 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15186) begin
                                                              _T_18065_48 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15184) begin
                                                                _T_18065_48 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15182) begin
                                                                  _T_18065_48 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15180) begin
                                                                    _T_18065_48 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15178) begin
                                                                      _T_18065_48 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15176) begin
                                                                        _T_18065_48 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15174) begin
                                                                          _T_18065_48 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15172) begin
                                                                            _T_18065_48 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15170) begin
                                                                              _T_18065_48 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15168) begin
                                                                                _T_18065_48 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15166) begin
                                                                                  _T_18065_48 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15164) begin
                                                                                    _T_18065_48 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15162) begin
                                                                                      _T_18065_48 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15160) begin
                                                                                        _T_18065_48 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15158) begin
                                                                                          _T_18065_48 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15156) begin
                                                                                            _T_18065_48 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15154) begin
                                                                                              _T_18065_48 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15152) begin
                                                                                                _T_18065_48 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15150) begin
                                                                                                  _T_18065_48 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15148) begin
                                                                                                    _T_18065_48 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15146) begin
                                                                                                      _T_18065_48 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15144) begin
                                                                                                        _T_18065_48 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15142) begin
                                                                                                          _T_18065_48 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          _T_18065_48 <= 8'h0;
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_48 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_49) begin
        if (_T_15389) begin
          _T_18065_49 <= _T_10366_0;
        end else begin
          if (_T_15387) begin
            _T_18065_49 <= _T_10366_1;
          end else begin
            if (_T_15385) begin
              _T_18065_49 <= _T_10366_2;
            end else begin
              if (_T_15383) begin
                _T_18065_49 <= _T_10366_3;
              end else begin
                if (_T_15381) begin
                  _T_18065_49 <= _T_10366_4;
                end else begin
                  if (_T_15379) begin
                    _T_18065_49 <= _T_10366_5;
                  end else begin
                    if (_T_15377) begin
                      _T_18065_49 <= _T_10366_6;
                    end else begin
                      if (_T_15375) begin
                        _T_18065_49 <= _T_10366_7;
                      end else begin
                        if (_T_15373) begin
                          _T_18065_49 <= _T_10366_8;
                        end else begin
                          if (_T_15371) begin
                            _T_18065_49 <= _T_10366_9;
                          end else begin
                            if (_T_15369) begin
                              _T_18065_49 <= _T_10366_10;
                            end else begin
                              if (_T_15367) begin
                                _T_18065_49 <= _T_10366_11;
                              end else begin
                                if (_T_15365) begin
                                  _T_18065_49 <= _T_10366_12;
                                end else begin
                                  if (_T_15363) begin
                                    _T_18065_49 <= _T_10366_13;
                                  end else begin
                                    if (_T_15361) begin
                                      _T_18065_49 <= _T_10366_14;
                                    end else begin
                                      if (_T_15359) begin
                                        _T_18065_49 <= _T_10366_15;
                                      end else begin
                                        if (_T_15357) begin
                                          _T_18065_49 <= _T_10366_16;
                                        end else begin
                                          if (_T_15355) begin
                                            _T_18065_49 <= _T_10366_17;
                                          end else begin
                                            if (_T_15353) begin
                                              _T_18065_49 <= _T_10366_18;
                                            end else begin
                                              if (_T_15351) begin
                                                _T_18065_49 <= _T_10366_19;
                                              end else begin
                                                if (_T_15349) begin
                                                  _T_18065_49 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15347) begin
                                                    _T_18065_49 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15345) begin
                                                      _T_18065_49 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15343) begin
                                                        _T_18065_49 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15341) begin
                                                          _T_18065_49 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15339) begin
                                                            _T_18065_49 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15337) begin
                                                              _T_18065_49 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15335) begin
                                                                _T_18065_49 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15333) begin
                                                                  _T_18065_49 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15331) begin
                                                                    _T_18065_49 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15329) begin
                                                                      _T_18065_49 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15327) begin
                                                                        _T_18065_49 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15325) begin
                                                                          _T_18065_49 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15323) begin
                                                                            _T_18065_49 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15321) begin
                                                                              _T_18065_49 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15319) begin
                                                                                _T_18065_49 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15317) begin
                                                                                  _T_18065_49 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15315) begin
                                                                                    _T_18065_49 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15313) begin
                                                                                      _T_18065_49 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15311) begin
                                                                                        _T_18065_49 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15309) begin
                                                                                          _T_18065_49 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15307) begin
                                                                                            _T_18065_49 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15305) begin
                                                                                              _T_18065_49 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15303) begin
                                                                                                _T_18065_49 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15301) begin
                                                                                                  _T_18065_49 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15299) begin
                                                                                                    _T_18065_49 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15297) begin
                                                                                                      _T_18065_49 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15295) begin
                                                                                                        _T_18065_49 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15293) begin
                                                                                                          _T_18065_49 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15291) begin
                                                                                                            _T_18065_49 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            _T_18065_49 <= 8'h0;
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_49 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_50) begin
        if (_T_15543) begin
          _T_18065_50 <= _T_10366_0;
        end else begin
          if (_T_15541) begin
            _T_18065_50 <= _T_10366_1;
          end else begin
            if (_T_15539) begin
              _T_18065_50 <= _T_10366_2;
            end else begin
              if (_T_15537) begin
                _T_18065_50 <= _T_10366_3;
              end else begin
                if (_T_15535) begin
                  _T_18065_50 <= _T_10366_4;
                end else begin
                  if (_T_15533) begin
                    _T_18065_50 <= _T_10366_5;
                  end else begin
                    if (_T_15531) begin
                      _T_18065_50 <= _T_10366_6;
                    end else begin
                      if (_T_15529) begin
                        _T_18065_50 <= _T_10366_7;
                      end else begin
                        if (_T_15527) begin
                          _T_18065_50 <= _T_10366_8;
                        end else begin
                          if (_T_15525) begin
                            _T_18065_50 <= _T_10366_9;
                          end else begin
                            if (_T_15523) begin
                              _T_18065_50 <= _T_10366_10;
                            end else begin
                              if (_T_15521) begin
                                _T_18065_50 <= _T_10366_11;
                              end else begin
                                if (_T_15519) begin
                                  _T_18065_50 <= _T_10366_12;
                                end else begin
                                  if (_T_15517) begin
                                    _T_18065_50 <= _T_10366_13;
                                  end else begin
                                    if (_T_15515) begin
                                      _T_18065_50 <= _T_10366_14;
                                    end else begin
                                      if (_T_15513) begin
                                        _T_18065_50 <= _T_10366_15;
                                      end else begin
                                        if (_T_15511) begin
                                          _T_18065_50 <= _T_10366_16;
                                        end else begin
                                          if (_T_15509) begin
                                            _T_18065_50 <= _T_10366_17;
                                          end else begin
                                            if (_T_15507) begin
                                              _T_18065_50 <= _T_10366_18;
                                            end else begin
                                              if (_T_15505) begin
                                                _T_18065_50 <= _T_10366_19;
                                              end else begin
                                                if (_T_15503) begin
                                                  _T_18065_50 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15501) begin
                                                    _T_18065_50 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15499) begin
                                                      _T_18065_50 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15497) begin
                                                        _T_18065_50 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15495) begin
                                                          _T_18065_50 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15493) begin
                                                            _T_18065_50 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15491) begin
                                                              _T_18065_50 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15489) begin
                                                                _T_18065_50 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15487) begin
                                                                  _T_18065_50 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15485) begin
                                                                    _T_18065_50 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15483) begin
                                                                      _T_18065_50 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15481) begin
                                                                        _T_18065_50 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15479) begin
                                                                          _T_18065_50 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15477) begin
                                                                            _T_18065_50 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15475) begin
                                                                              _T_18065_50 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15473) begin
                                                                                _T_18065_50 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15471) begin
                                                                                  _T_18065_50 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15469) begin
                                                                                    _T_18065_50 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15467) begin
                                                                                      _T_18065_50 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15465) begin
                                                                                        _T_18065_50 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15463) begin
                                                                                          _T_18065_50 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15461) begin
                                                                                            _T_18065_50 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15459) begin
                                                                                              _T_18065_50 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15457) begin
                                                                                                _T_18065_50 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15455) begin
                                                                                                  _T_18065_50 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15453) begin
                                                                                                    _T_18065_50 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15451) begin
                                                                                                      _T_18065_50 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15449) begin
                                                                                                        _T_18065_50 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15447) begin
                                                                                                          _T_18065_50 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15445) begin
                                                                                                            _T_18065_50 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15443) begin
                                                                                                              _T_18065_50 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              _T_18065_50 <= 8'h0;
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_50 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_51) begin
        if (_T_15700) begin
          _T_18065_51 <= _T_10366_0;
        end else begin
          if (_T_15698) begin
            _T_18065_51 <= _T_10366_1;
          end else begin
            if (_T_15696) begin
              _T_18065_51 <= _T_10366_2;
            end else begin
              if (_T_15694) begin
                _T_18065_51 <= _T_10366_3;
              end else begin
                if (_T_15692) begin
                  _T_18065_51 <= _T_10366_4;
                end else begin
                  if (_T_15690) begin
                    _T_18065_51 <= _T_10366_5;
                  end else begin
                    if (_T_15688) begin
                      _T_18065_51 <= _T_10366_6;
                    end else begin
                      if (_T_15686) begin
                        _T_18065_51 <= _T_10366_7;
                      end else begin
                        if (_T_15684) begin
                          _T_18065_51 <= _T_10366_8;
                        end else begin
                          if (_T_15682) begin
                            _T_18065_51 <= _T_10366_9;
                          end else begin
                            if (_T_15680) begin
                              _T_18065_51 <= _T_10366_10;
                            end else begin
                              if (_T_15678) begin
                                _T_18065_51 <= _T_10366_11;
                              end else begin
                                if (_T_15676) begin
                                  _T_18065_51 <= _T_10366_12;
                                end else begin
                                  if (_T_15674) begin
                                    _T_18065_51 <= _T_10366_13;
                                  end else begin
                                    if (_T_15672) begin
                                      _T_18065_51 <= _T_10366_14;
                                    end else begin
                                      if (_T_15670) begin
                                        _T_18065_51 <= _T_10366_15;
                                      end else begin
                                        if (_T_15668) begin
                                          _T_18065_51 <= _T_10366_16;
                                        end else begin
                                          if (_T_15666) begin
                                            _T_18065_51 <= _T_10366_17;
                                          end else begin
                                            if (_T_15664) begin
                                              _T_18065_51 <= _T_10366_18;
                                            end else begin
                                              if (_T_15662) begin
                                                _T_18065_51 <= _T_10366_19;
                                              end else begin
                                                if (_T_15660) begin
                                                  _T_18065_51 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15658) begin
                                                    _T_18065_51 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15656) begin
                                                      _T_18065_51 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15654) begin
                                                        _T_18065_51 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15652) begin
                                                          _T_18065_51 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15650) begin
                                                            _T_18065_51 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15648) begin
                                                              _T_18065_51 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15646) begin
                                                                _T_18065_51 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15644) begin
                                                                  _T_18065_51 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15642) begin
                                                                    _T_18065_51 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15640) begin
                                                                      _T_18065_51 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15638) begin
                                                                        _T_18065_51 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15636) begin
                                                                          _T_18065_51 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15634) begin
                                                                            _T_18065_51 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15632) begin
                                                                              _T_18065_51 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15630) begin
                                                                                _T_18065_51 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15628) begin
                                                                                  _T_18065_51 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15626) begin
                                                                                    _T_18065_51 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15624) begin
                                                                                      _T_18065_51 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15622) begin
                                                                                        _T_18065_51 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15620) begin
                                                                                          _T_18065_51 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15618) begin
                                                                                            _T_18065_51 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15616) begin
                                                                                              _T_18065_51 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15614) begin
                                                                                                _T_18065_51 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15612) begin
                                                                                                  _T_18065_51 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15610) begin
                                                                                                    _T_18065_51 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15608) begin
                                                                                                      _T_18065_51 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15606) begin
                                                                                                        _T_18065_51 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15604) begin
                                                                                                          _T_18065_51 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15602) begin
                                                                                                            _T_18065_51 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15600) begin
                                                                                                              _T_18065_51 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15598) begin
                                                                                                                _T_18065_51 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                _T_18065_51 <= 8'h0;
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_51 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_52) begin
        if (_T_15860) begin
          _T_18065_52 <= _T_10366_0;
        end else begin
          if (_T_15858) begin
            _T_18065_52 <= _T_10366_1;
          end else begin
            if (_T_15856) begin
              _T_18065_52 <= _T_10366_2;
            end else begin
              if (_T_15854) begin
                _T_18065_52 <= _T_10366_3;
              end else begin
                if (_T_15852) begin
                  _T_18065_52 <= _T_10366_4;
                end else begin
                  if (_T_15850) begin
                    _T_18065_52 <= _T_10366_5;
                  end else begin
                    if (_T_15848) begin
                      _T_18065_52 <= _T_10366_6;
                    end else begin
                      if (_T_15846) begin
                        _T_18065_52 <= _T_10366_7;
                      end else begin
                        if (_T_15844) begin
                          _T_18065_52 <= _T_10366_8;
                        end else begin
                          if (_T_15842) begin
                            _T_18065_52 <= _T_10366_9;
                          end else begin
                            if (_T_15840) begin
                              _T_18065_52 <= _T_10366_10;
                            end else begin
                              if (_T_15838) begin
                                _T_18065_52 <= _T_10366_11;
                              end else begin
                                if (_T_15836) begin
                                  _T_18065_52 <= _T_10366_12;
                                end else begin
                                  if (_T_15834) begin
                                    _T_18065_52 <= _T_10366_13;
                                  end else begin
                                    if (_T_15832) begin
                                      _T_18065_52 <= _T_10366_14;
                                    end else begin
                                      if (_T_15830) begin
                                        _T_18065_52 <= _T_10366_15;
                                      end else begin
                                        if (_T_15828) begin
                                          _T_18065_52 <= _T_10366_16;
                                        end else begin
                                          if (_T_15826) begin
                                            _T_18065_52 <= _T_10366_17;
                                          end else begin
                                            if (_T_15824) begin
                                              _T_18065_52 <= _T_10366_18;
                                            end else begin
                                              if (_T_15822) begin
                                                _T_18065_52 <= _T_10366_19;
                                              end else begin
                                                if (_T_15820) begin
                                                  _T_18065_52 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15818) begin
                                                    _T_18065_52 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15816) begin
                                                      _T_18065_52 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15814) begin
                                                        _T_18065_52 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15812) begin
                                                          _T_18065_52 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15810) begin
                                                            _T_18065_52 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15808) begin
                                                              _T_18065_52 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15806) begin
                                                                _T_18065_52 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15804) begin
                                                                  _T_18065_52 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15802) begin
                                                                    _T_18065_52 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15800) begin
                                                                      _T_18065_52 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15798) begin
                                                                        _T_18065_52 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15796) begin
                                                                          _T_18065_52 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15794) begin
                                                                            _T_18065_52 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15792) begin
                                                                              _T_18065_52 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15790) begin
                                                                                _T_18065_52 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15788) begin
                                                                                  _T_18065_52 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15786) begin
                                                                                    _T_18065_52 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15784) begin
                                                                                      _T_18065_52 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15782) begin
                                                                                        _T_18065_52 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15780) begin
                                                                                          _T_18065_52 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15778) begin
                                                                                            _T_18065_52 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15776) begin
                                                                                              _T_18065_52 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15774) begin
                                                                                                _T_18065_52 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15772) begin
                                                                                                  _T_18065_52 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15770) begin
                                                                                                    _T_18065_52 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15768) begin
                                                                                                      _T_18065_52 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15766) begin
                                                                                                        _T_18065_52 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15764) begin
                                                                                                          _T_18065_52 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15762) begin
                                                                                                            _T_18065_52 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15760) begin
                                                                                                              _T_18065_52 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15758) begin
                                                                                                                _T_18065_52 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_15756) begin
                                                                                                                  _T_18065_52 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  _T_18065_52 <= 8'h0;
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_52 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_53) begin
        if (_T_16023) begin
          _T_18065_53 <= _T_10366_0;
        end else begin
          if (_T_16021) begin
            _T_18065_53 <= _T_10366_1;
          end else begin
            if (_T_16019) begin
              _T_18065_53 <= _T_10366_2;
            end else begin
              if (_T_16017) begin
                _T_18065_53 <= _T_10366_3;
              end else begin
                if (_T_16015) begin
                  _T_18065_53 <= _T_10366_4;
                end else begin
                  if (_T_16013) begin
                    _T_18065_53 <= _T_10366_5;
                  end else begin
                    if (_T_16011) begin
                      _T_18065_53 <= _T_10366_6;
                    end else begin
                      if (_T_16009) begin
                        _T_18065_53 <= _T_10366_7;
                      end else begin
                        if (_T_16007) begin
                          _T_18065_53 <= _T_10366_8;
                        end else begin
                          if (_T_16005) begin
                            _T_18065_53 <= _T_10366_9;
                          end else begin
                            if (_T_16003) begin
                              _T_18065_53 <= _T_10366_10;
                            end else begin
                              if (_T_16001) begin
                                _T_18065_53 <= _T_10366_11;
                              end else begin
                                if (_T_15999) begin
                                  _T_18065_53 <= _T_10366_12;
                                end else begin
                                  if (_T_15997) begin
                                    _T_18065_53 <= _T_10366_13;
                                  end else begin
                                    if (_T_15995) begin
                                      _T_18065_53 <= _T_10366_14;
                                    end else begin
                                      if (_T_15993) begin
                                        _T_18065_53 <= _T_10366_15;
                                      end else begin
                                        if (_T_15991) begin
                                          _T_18065_53 <= _T_10366_16;
                                        end else begin
                                          if (_T_15989) begin
                                            _T_18065_53 <= _T_10366_17;
                                          end else begin
                                            if (_T_15987) begin
                                              _T_18065_53 <= _T_10366_18;
                                            end else begin
                                              if (_T_15985) begin
                                                _T_18065_53 <= _T_10366_19;
                                              end else begin
                                                if (_T_15983) begin
                                                  _T_18065_53 <= _T_10366_20;
                                                end else begin
                                                  if (_T_15981) begin
                                                    _T_18065_53 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_15979) begin
                                                      _T_18065_53 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_15977) begin
                                                        _T_18065_53 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_15975) begin
                                                          _T_18065_53 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_15973) begin
                                                            _T_18065_53 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_15971) begin
                                                              _T_18065_53 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_15969) begin
                                                                _T_18065_53 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_15967) begin
                                                                  _T_18065_53 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_15965) begin
                                                                    _T_18065_53 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_15963) begin
                                                                      _T_18065_53 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_15961) begin
                                                                        _T_18065_53 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_15959) begin
                                                                          _T_18065_53 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_15957) begin
                                                                            _T_18065_53 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_15955) begin
                                                                              _T_18065_53 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_15953) begin
                                                                                _T_18065_53 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_15951) begin
                                                                                  _T_18065_53 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_15949) begin
                                                                                    _T_18065_53 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_15947) begin
                                                                                      _T_18065_53 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_15945) begin
                                                                                        _T_18065_53 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_15943) begin
                                                                                          _T_18065_53 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_15941) begin
                                                                                            _T_18065_53 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_15939) begin
                                                                                              _T_18065_53 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_15937) begin
                                                                                                _T_18065_53 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_15935) begin
                                                                                                  _T_18065_53 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_15933) begin
                                                                                                    _T_18065_53 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_15931) begin
                                                                                                      _T_18065_53 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_15929) begin
                                                                                                        _T_18065_53 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_15927) begin
                                                                                                          _T_18065_53 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_15925) begin
                                                                                                            _T_18065_53 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_15923) begin
                                                                                                              _T_18065_53 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_15921) begin
                                                                                                                _T_18065_53 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_15919) begin
                                                                                                                  _T_18065_53 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_15917) begin
                                                                                                                    _T_18065_53 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    _T_18065_53 <= 8'h0;
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_53 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_54) begin
        if (_T_16189) begin
          _T_18065_54 <= _T_10366_0;
        end else begin
          if (_T_16187) begin
            _T_18065_54 <= _T_10366_1;
          end else begin
            if (_T_16185) begin
              _T_18065_54 <= _T_10366_2;
            end else begin
              if (_T_16183) begin
                _T_18065_54 <= _T_10366_3;
              end else begin
                if (_T_16181) begin
                  _T_18065_54 <= _T_10366_4;
                end else begin
                  if (_T_16179) begin
                    _T_18065_54 <= _T_10366_5;
                  end else begin
                    if (_T_16177) begin
                      _T_18065_54 <= _T_10366_6;
                    end else begin
                      if (_T_16175) begin
                        _T_18065_54 <= _T_10366_7;
                      end else begin
                        if (_T_16173) begin
                          _T_18065_54 <= _T_10366_8;
                        end else begin
                          if (_T_16171) begin
                            _T_18065_54 <= _T_10366_9;
                          end else begin
                            if (_T_16169) begin
                              _T_18065_54 <= _T_10366_10;
                            end else begin
                              if (_T_16167) begin
                                _T_18065_54 <= _T_10366_11;
                              end else begin
                                if (_T_16165) begin
                                  _T_18065_54 <= _T_10366_12;
                                end else begin
                                  if (_T_16163) begin
                                    _T_18065_54 <= _T_10366_13;
                                  end else begin
                                    if (_T_16161) begin
                                      _T_18065_54 <= _T_10366_14;
                                    end else begin
                                      if (_T_16159) begin
                                        _T_18065_54 <= _T_10366_15;
                                      end else begin
                                        if (_T_16157) begin
                                          _T_18065_54 <= _T_10366_16;
                                        end else begin
                                          if (_T_16155) begin
                                            _T_18065_54 <= _T_10366_17;
                                          end else begin
                                            if (_T_16153) begin
                                              _T_18065_54 <= _T_10366_18;
                                            end else begin
                                              if (_T_16151) begin
                                                _T_18065_54 <= _T_10366_19;
                                              end else begin
                                                if (_T_16149) begin
                                                  _T_18065_54 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16147) begin
                                                    _T_18065_54 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16145) begin
                                                      _T_18065_54 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16143) begin
                                                        _T_18065_54 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16141) begin
                                                          _T_18065_54 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16139) begin
                                                            _T_18065_54 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16137) begin
                                                              _T_18065_54 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16135) begin
                                                                _T_18065_54 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16133) begin
                                                                  _T_18065_54 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16131) begin
                                                                    _T_18065_54 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16129) begin
                                                                      _T_18065_54 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16127) begin
                                                                        _T_18065_54 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16125) begin
                                                                          _T_18065_54 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16123) begin
                                                                            _T_18065_54 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16121) begin
                                                                              _T_18065_54 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16119) begin
                                                                                _T_18065_54 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16117) begin
                                                                                  _T_18065_54 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16115) begin
                                                                                    _T_18065_54 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16113) begin
                                                                                      _T_18065_54 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16111) begin
                                                                                        _T_18065_54 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16109) begin
                                                                                          _T_18065_54 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16107) begin
                                                                                            _T_18065_54 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16105) begin
                                                                                              _T_18065_54 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16103) begin
                                                                                                _T_18065_54 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16101) begin
                                                                                                  _T_18065_54 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16099) begin
                                                                                                    _T_18065_54 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16097) begin
                                                                                                      _T_18065_54 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16095) begin
                                                                                                        _T_18065_54 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16093) begin
                                                                                                          _T_18065_54 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16091) begin
                                                                                                            _T_18065_54 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16089) begin
                                                                                                              _T_18065_54 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16087) begin
                                                                                                                _T_18065_54 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16085) begin
                                                                                                                  _T_18065_54 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16083) begin
                                                                                                                    _T_18065_54 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16081) begin
                                                                                                                      _T_18065_54 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      _T_18065_54 <= 8'h0;
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_54 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_55) begin
        if (_T_16358) begin
          _T_18065_55 <= _T_10366_0;
        end else begin
          if (_T_16356) begin
            _T_18065_55 <= _T_10366_1;
          end else begin
            if (_T_16354) begin
              _T_18065_55 <= _T_10366_2;
            end else begin
              if (_T_16352) begin
                _T_18065_55 <= _T_10366_3;
              end else begin
                if (_T_16350) begin
                  _T_18065_55 <= _T_10366_4;
                end else begin
                  if (_T_16348) begin
                    _T_18065_55 <= _T_10366_5;
                  end else begin
                    if (_T_16346) begin
                      _T_18065_55 <= _T_10366_6;
                    end else begin
                      if (_T_16344) begin
                        _T_18065_55 <= _T_10366_7;
                      end else begin
                        if (_T_16342) begin
                          _T_18065_55 <= _T_10366_8;
                        end else begin
                          if (_T_16340) begin
                            _T_18065_55 <= _T_10366_9;
                          end else begin
                            if (_T_16338) begin
                              _T_18065_55 <= _T_10366_10;
                            end else begin
                              if (_T_16336) begin
                                _T_18065_55 <= _T_10366_11;
                              end else begin
                                if (_T_16334) begin
                                  _T_18065_55 <= _T_10366_12;
                                end else begin
                                  if (_T_16332) begin
                                    _T_18065_55 <= _T_10366_13;
                                  end else begin
                                    if (_T_16330) begin
                                      _T_18065_55 <= _T_10366_14;
                                    end else begin
                                      if (_T_16328) begin
                                        _T_18065_55 <= _T_10366_15;
                                      end else begin
                                        if (_T_16326) begin
                                          _T_18065_55 <= _T_10366_16;
                                        end else begin
                                          if (_T_16324) begin
                                            _T_18065_55 <= _T_10366_17;
                                          end else begin
                                            if (_T_16322) begin
                                              _T_18065_55 <= _T_10366_18;
                                            end else begin
                                              if (_T_16320) begin
                                                _T_18065_55 <= _T_10366_19;
                                              end else begin
                                                if (_T_16318) begin
                                                  _T_18065_55 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16316) begin
                                                    _T_18065_55 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16314) begin
                                                      _T_18065_55 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16312) begin
                                                        _T_18065_55 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16310) begin
                                                          _T_18065_55 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16308) begin
                                                            _T_18065_55 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16306) begin
                                                              _T_18065_55 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16304) begin
                                                                _T_18065_55 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16302) begin
                                                                  _T_18065_55 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16300) begin
                                                                    _T_18065_55 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16298) begin
                                                                      _T_18065_55 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16296) begin
                                                                        _T_18065_55 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16294) begin
                                                                          _T_18065_55 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16292) begin
                                                                            _T_18065_55 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16290) begin
                                                                              _T_18065_55 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16288) begin
                                                                                _T_18065_55 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16286) begin
                                                                                  _T_18065_55 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16284) begin
                                                                                    _T_18065_55 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16282) begin
                                                                                      _T_18065_55 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16280) begin
                                                                                        _T_18065_55 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16278) begin
                                                                                          _T_18065_55 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16276) begin
                                                                                            _T_18065_55 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16274) begin
                                                                                              _T_18065_55 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16272) begin
                                                                                                _T_18065_55 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16270) begin
                                                                                                  _T_18065_55 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16268) begin
                                                                                                    _T_18065_55 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16266) begin
                                                                                                      _T_18065_55 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16264) begin
                                                                                                        _T_18065_55 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16262) begin
                                                                                                          _T_18065_55 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16260) begin
                                                                                                            _T_18065_55 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16258) begin
                                                                                                              _T_18065_55 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16256) begin
                                                                                                                _T_18065_55 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16254) begin
                                                                                                                  _T_18065_55 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16252) begin
                                                                                                                    _T_18065_55 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16250) begin
                                                                                                                      _T_18065_55 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16248) begin
                                                                                                                        _T_18065_55 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        _T_18065_55 <= 8'h0;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_55 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_56) begin
        if (_T_16530) begin
          _T_18065_56 <= _T_10366_0;
        end else begin
          if (_T_16528) begin
            _T_18065_56 <= _T_10366_1;
          end else begin
            if (_T_16526) begin
              _T_18065_56 <= _T_10366_2;
            end else begin
              if (_T_16524) begin
                _T_18065_56 <= _T_10366_3;
              end else begin
                if (_T_16522) begin
                  _T_18065_56 <= _T_10366_4;
                end else begin
                  if (_T_16520) begin
                    _T_18065_56 <= _T_10366_5;
                  end else begin
                    if (_T_16518) begin
                      _T_18065_56 <= _T_10366_6;
                    end else begin
                      if (_T_16516) begin
                        _T_18065_56 <= _T_10366_7;
                      end else begin
                        if (_T_16514) begin
                          _T_18065_56 <= _T_10366_8;
                        end else begin
                          if (_T_16512) begin
                            _T_18065_56 <= _T_10366_9;
                          end else begin
                            if (_T_16510) begin
                              _T_18065_56 <= _T_10366_10;
                            end else begin
                              if (_T_16508) begin
                                _T_18065_56 <= _T_10366_11;
                              end else begin
                                if (_T_16506) begin
                                  _T_18065_56 <= _T_10366_12;
                                end else begin
                                  if (_T_16504) begin
                                    _T_18065_56 <= _T_10366_13;
                                  end else begin
                                    if (_T_16502) begin
                                      _T_18065_56 <= _T_10366_14;
                                    end else begin
                                      if (_T_16500) begin
                                        _T_18065_56 <= _T_10366_15;
                                      end else begin
                                        if (_T_16498) begin
                                          _T_18065_56 <= _T_10366_16;
                                        end else begin
                                          if (_T_16496) begin
                                            _T_18065_56 <= _T_10366_17;
                                          end else begin
                                            if (_T_16494) begin
                                              _T_18065_56 <= _T_10366_18;
                                            end else begin
                                              if (_T_16492) begin
                                                _T_18065_56 <= _T_10366_19;
                                              end else begin
                                                if (_T_16490) begin
                                                  _T_18065_56 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16488) begin
                                                    _T_18065_56 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16486) begin
                                                      _T_18065_56 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16484) begin
                                                        _T_18065_56 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16482) begin
                                                          _T_18065_56 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16480) begin
                                                            _T_18065_56 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16478) begin
                                                              _T_18065_56 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16476) begin
                                                                _T_18065_56 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16474) begin
                                                                  _T_18065_56 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16472) begin
                                                                    _T_18065_56 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16470) begin
                                                                      _T_18065_56 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16468) begin
                                                                        _T_18065_56 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16466) begin
                                                                          _T_18065_56 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16464) begin
                                                                            _T_18065_56 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16462) begin
                                                                              _T_18065_56 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16460) begin
                                                                                _T_18065_56 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16458) begin
                                                                                  _T_18065_56 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16456) begin
                                                                                    _T_18065_56 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16454) begin
                                                                                      _T_18065_56 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16452) begin
                                                                                        _T_18065_56 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16450) begin
                                                                                          _T_18065_56 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16448) begin
                                                                                            _T_18065_56 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16446) begin
                                                                                              _T_18065_56 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16444) begin
                                                                                                _T_18065_56 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16442) begin
                                                                                                  _T_18065_56 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16440) begin
                                                                                                    _T_18065_56 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16438) begin
                                                                                                      _T_18065_56 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16436) begin
                                                                                                        _T_18065_56 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16434) begin
                                                                                                          _T_18065_56 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16432) begin
                                                                                                            _T_18065_56 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16430) begin
                                                                                                              _T_18065_56 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16428) begin
                                                                                                                _T_18065_56 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16426) begin
                                                                                                                  _T_18065_56 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16424) begin
                                                                                                                    _T_18065_56 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16422) begin
                                                                                                                      _T_18065_56 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16420) begin
                                                                                                                        _T_18065_56 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16418) begin
                                                                                                                          _T_18065_56 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          _T_18065_56 <= 8'h0;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_56 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_57) begin
        if (_T_16705) begin
          _T_18065_57 <= _T_10366_0;
        end else begin
          if (_T_16703) begin
            _T_18065_57 <= _T_10366_1;
          end else begin
            if (_T_16701) begin
              _T_18065_57 <= _T_10366_2;
            end else begin
              if (_T_16699) begin
                _T_18065_57 <= _T_10366_3;
              end else begin
                if (_T_16697) begin
                  _T_18065_57 <= _T_10366_4;
                end else begin
                  if (_T_16695) begin
                    _T_18065_57 <= _T_10366_5;
                  end else begin
                    if (_T_16693) begin
                      _T_18065_57 <= _T_10366_6;
                    end else begin
                      if (_T_16691) begin
                        _T_18065_57 <= _T_10366_7;
                      end else begin
                        if (_T_16689) begin
                          _T_18065_57 <= _T_10366_8;
                        end else begin
                          if (_T_16687) begin
                            _T_18065_57 <= _T_10366_9;
                          end else begin
                            if (_T_16685) begin
                              _T_18065_57 <= _T_10366_10;
                            end else begin
                              if (_T_16683) begin
                                _T_18065_57 <= _T_10366_11;
                              end else begin
                                if (_T_16681) begin
                                  _T_18065_57 <= _T_10366_12;
                                end else begin
                                  if (_T_16679) begin
                                    _T_18065_57 <= _T_10366_13;
                                  end else begin
                                    if (_T_16677) begin
                                      _T_18065_57 <= _T_10366_14;
                                    end else begin
                                      if (_T_16675) begin
                                        _T_18065_57 <= _T_10366_15;
                                      end else begin
                                        if (_T_16673) begin
                                          _T_18065_57 <= _T_10366_16;
                                        end else begin
                                          if (_T_16671) begin
                                            _T_18065_57 <= _T_10366_17;
                                          end else begin
                                            if (_T_16669) begin
                                              _T_18065_57 <= _T_10366_18;
                                            end else begin
                                              if (_T_16667) begin
                                                _T_18065_57 <= _T_10366_19;
                                              end else begin
                                                if (_T_16665) begin
                                                  _T_18065_57 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16663) begin
                                                    _T_18065_57 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16661) begin
                                                      _T_18065_57 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16659) begin
                                                        _T_18065_57 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16657) begin
                                                          _T_18065_57 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16655) begin
                                                            _T_18065_57 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16653) begin
                                                              _T_18065_57 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16651) begin
                                                                _T_18065_57 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16649) begin
                                                                  _T_18065_57 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16647) begin
                                                                    _T_18065_57 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16645) begin
                                                                      _T_18065_57 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16643) begin
                                                                        _T_18065_57 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16641) begin
                                                                          _T_18065_57 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16639) begin
                                                                            _T_18065_57 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16637) begin
                                                                              _T_18065_57 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16635) begin
                                                                                _T_18065_57 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16633) begin
                                                                                  _T_18065_57 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16631) begin
                                                                                    _T_18065_57 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16629) begin
                                                                                      _T_18065_57 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16627) begin
                                                                                        _T_18065_57 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16625) begin
                                                                                          _T_18065_57 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16623) begin
                                                                                            _T_18065_57 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16621) begin
                                                                                              _T_18065_57 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16619) begin
                                                                                                _T_18065_57 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16617) begin
                                                                                                  _T_18065_57 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16615) begin
                                                                                                    _T_18065_57 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16613) begin
                                                                                                      _T_18065_57 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16611) begin
                                                                                                        _T_18065_57 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16609) begin
                                                                                                          _T_18065_57 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16607) begin
                                                                                                            _T_18065_57 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16605) begin
                                                                                                              _T_18065_57 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16603) begin
                                                                                                                _T_18065_57 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16601) begin
                                                                                                                  _T_18065_57 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16599) begin
                                                                                                                    _T_18065_57 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16597) begin
                                                                                                                      _T_18065_57 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16595) begin
                                                                                                                        _T_18065_57 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16593) begin
                                                                                                                          _T_18065_57 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16591) begin
                                                                                                                            _T_18065_57 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            _T_18065_57 <= 8'h0;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_57 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_58) begin
        if (_T_16883) begin
          _T_18065_58 <= _T_10366_0;
        end else begin
          if (_T_16881) begin
            _T_18065_58 <= _T_10366_1;
          end else begin
            if (_T_16879) begin
              _T_18065_58 <= _T_10366_2;
            end else begin
              if (_T_16877) begin
                _T_18065_58 <= _T_10366_3;
              end else begin
                if (_T_16875) begin
                  _T_18065_58 <= _T_10366_4;
                end else begin
                  if (_T_16873) begin
                    _T_18065_58 <= _T_10366_5;
                  end else begin
                    if (_T_16871) begin
                      _T_18065_58 <= _T_10366_6;
                    end else begin
                      if (_T_16869) begin
                        _T_18065_58 <= _T_10366_7;
                      end else begin
                        if (_T_16867) begin
                          _T_18065_58 <= _T_10366_8;
                        end else begin
                          if (_T_16865) begin
                            _T_18065_58 <= _T_10366_9;
                          end else begin
                            if (_T_16863) begin
                              _T_18065_58 <= _T_10366_10;
                            end else begin
                              if (_T_16861) begin
                                _T_18065_58 <= _T_10366_11;
                              end else begin
                                if (_T_16859) begin
                                  _T_18065_58 <= _T_10366_12;
                                end else begin
                                  if (_T_16857) begin
                                    _T_18065_58 <= _T_10366_13;
                                  end else begin
                                    if (_T_16855) begin
                                      _T_18065_58 <= _T_10366_14;
                                    end else begin
                                      if (_T_16853) begin
                                        _T_18065_58 <= _T_10366_15;
                                      end else begin
                                        if (_T_16851) begin
                                          _T_18065_58 <= _T_10366_16;
                                        end else begin
                                          if (_T_16849) begin
                                            _T_18065_58 <= _T_10366_17;
                                          end else begin
                                            if (_T_16847) begin
                                              _T_18065_58 <= _T_10366_18;
                                            end else begin
                                              if (_T_16845) begin
                                                _T_18065_58 <= _T_10366_19;
                                              end else begin
                                                if (_T_16843) begin
                                                  _T_18065_58 <= _T_10366_20;
                                                end else begin
                                                  if (_T_16841) begin
                                                    _T_18065_58 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_16839) begin
                                                      _T_18065_58 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_16837) begin
                                                        _T_18065_58 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_16835) begin
                                                          _T_18065_58 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_16833) begin
                                                            _T_18065_58 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_16831) begin
                                                              _T_18065_58 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_16829) begin
                                                                _T_18065_58 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_16827) begin
                                                                  _T_18065_58 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_16825) begin
                                                                    _T_18065_58 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_16823) begin
                                                                      _T_18065_58 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_16821) begin
                                                                        _T_18065_58 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_16819) begin
                                                                          _T_18065_58 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16817) begin
                                                                            _T_18065_58 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16815) begin
                                                                              _T_18065_58 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16813) begin
                                                                                _T_18065_58 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16811) begin
                                                                                  _T_18065_58 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16809) begin
                                                                                    _T_18065_58 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16807) begin
                                                                                      _T_18065_58 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16805) begin
                                                                                        _T_18065_58 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16803) begin
                                                                                          _T_18065_58 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16801) begin
                                                                                            _T_18065_58 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16799) begin
                                                                                              _T_18065_58 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16797) begin
                                                                                                _T_18065_58 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16795) begin
                                                                                                  _T_18065_58 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16793) begin
                                                                                                    _T_18065_58 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16791) begin
                                                                                                      _T_18065_58 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16789) begin
                                                                                                        _T_18065_58 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16787) begin
                                                                                                          _T_18065_58 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16785) begin
                                                                                                            _T_18065_58 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16783) begin
                                                                                                              _T_18065_58 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16781) begin
                                                                                                                _T_18065_58 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16779) begin
                                                                                                                  _T_18065_58 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16777) begin
                                                                                                                    _T_18065_58 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16775) begin
                                                                                                                      _T_18065_58 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16773) begin
                                                                                                                        _T_18065_58 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16771) begin
                                                                                                                          _T_18065_58 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16769) begin
                                                                                                                            _T_18065_58 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16767) begin
                                                                                                                              _T_18065_58 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              _T_18065_58 <= 8'h0;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_58 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_59) begin
        if (_T_17064) begin
          _T_18065_59 <= _T_10366_0;
        end else begin
          if (_T_17062) begin
            _T_18065_59 <= _T_10366_1;
          end else begin
            if (_T_17060) begin
              _T_18065_59 <= _T_10366_2;
            end else begin
              if (_T_17058) begin
                _T_18065_59 <= _T_10366_3;
              end else begin
                if (_T_17056) begin
                  _T_18065_59 <= _T_10366_4;
                end else begin
                  if (_T_17054) begin
                    _T_18065_59 <= _T_10366_5;
                  end else begin
                    if (_T_17052) begin
                      _T_18065_59 <= _T_10366_6;
                    end else begin
                      if (_T_17050) begin
                        _T_18065_59 <= _T_10366_7;
                      end else begin
                        if (_T_17048) begin
                          _T_18065_59 <= _T_10366_8;
                        end else begin
                          if (_T_17046) begin
                            _T_18065_59 <= _T_10366_9;
                          end else begin
                            if (_T_17044) begin
                              _T_18065_59 <= _T_10366_10;
                            end else begin
                              if (_T_17042) begin
                                _T_18065_59 <= _T_10366_11;
                              end else begin
                                if (_T_17040) begin
                                  _T_18065_59 <= _T_10366_12;
                                end else begin
                                  if (_T_17038) begin
                                    _T_18065_59 <= _T_10366_13;
                                  end else begin
                                    if (_T_17036) begin
                                      _T_18065_59 <= _T_10366_14;
                                    end else begin
                                      if (_T_17034) begin
                                        _T_18065_59 <= _T_10366_15;
                                      end else begin
                                        if (_T_17032) begin
                                          _T_18065_59 <= _T_10366_16;
                                        end else begin
                                          if (_T_17030) begin
                                            _T_18065_59 <= _T_10366_17;
                                          end else begin
                                            if (_T_17028) begin
                                              _T_18065_59 <= _T_10366_18;
                                            end else begin
                                              if (_T_17026) begin
                                                _T_18065_59 <= _T_10366_19;
                                              end else begin
                                                if (_T_17024) begin
                                                  _T_18065_59 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17022) begin
                                                    _T_18065_59 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17020) begin
                                                      _T_18065_59 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17018) begin
                                                        _T_18065_59 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17016) begin
                                                          _T_18065_59 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17014) begin
                                                            _T_18065_59 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17012) begin
                                                              _T_18065_59 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17010) begin
                                                                _T_18065_59 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17008) begin
                                                                  _T_18065_59 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17006) begin
                                                                    _T_18065_59 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17004) begin
                                                                      _T_18065_59 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17002) begin
                                                                        _T_18065_59 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17000) begin
                                                                          _T_18065_59 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_16998) begin
                                                                            _T_18065_59 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_16996) begin
                                                                              _T_18065_59 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_16994) begin
                                                                                _T_18065_59 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_16992) begin
                                                                                  _T_18065_59 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_16990) begin
                                                                                    _T_18065_59 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_16988) begin
                                                                                      _T_18065_59 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_16986) begin
                                                                                        _T_18065_59 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_16984) begin
                                                                                          _T_18065_59 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_16982) begin
                                                                                            _T_18065_59 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_16980) begin
                                                                                              _T_18065_59 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_16978) begin
                                                                                                _T_18065_59 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_16976) begin
                                                                                                  _T_18065_59 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_16974) begin
                                                                                                    _T_18065_59 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_16972) begin
                                                                                                      _T_18065_59 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_16970) begin
                                                                                                        _T_18065_59 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_16968) begin
                                                                                                          _T_18065_59 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_16966) begin
                                                                                                            _T_18065_59 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_16964) begin
                                                                                                              _T_18065_59 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_16962) begin
                                                                                                                _T_18065_59 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_16960) begin
                                                                                                                  _T_18065_59 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_16958) begin
                                                                                                                    _T_18065_59 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_16956) begin
                                                                                                                      _T_18065_59 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_16954) begin
                                                                                                                        _T_18065_59 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_16952) begin
                                                                                                                          _T_18065_59 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_16950) begin
                                                                                                                            _T_18065_59 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_16948) begin
                                                                                                                              _T_18065_59 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_16946) begin
                                                                                                                                _T_18065_59 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                _T_18065_59 <= 8'h0;
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_59 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_60) begin
        if (_T_17248) begin
          _T_18065_60 <= _T_10366_0;
        end else begin
          if (_T_17246) begin
            _T_18065_60 <= _T_10366_1;
          end else begin
            if (_T_17244) begin
              _T_18065_60 <= _T_10366_2;
            end else begin
              if (_T_17242) begin
                _T_18065_60 <= _T_10366_3;
              end else begin
                if (_T_17240) begin
                  _T_18065_60 <= _T_10366_4;
                end else begin
                  if (_T_17238) begin
                    _T_18065_60 <= _T_10366_5;
                  end else begin
                    if (_T_17236) begin
                      _T_18065_60 <= _T_10366_6;
                    end else begin
                      if (_T_17234) begin
                        _T_18065_60 <= _T_10366_7;
                      end else begin
                        if (_T_17232) begin
                          _T_18065_60 <= _T_10366_8;
                        end else begin
                          if (_T_17230) begin
                            _T_18065_60 <= _T_10366_9;
                          end else begin
                            if (_T_17228) begin
                              _T_18065_60 <= _T_10366_10;
                            end else begin
                              if (_T_17226) begin
                                _T_18065_60 <= _T_10366_11;
                              end else begin
                                if (_T_17224) begin
                                  _T_18065_60 <= _T_10366_12;
                                end else begin
                                  if (_T_17222) begin
                                    _T_18065_60 <= _T_10366_13;
                                  end else begin
                                    if (_T_17220) begin
                                      _T_18065_60 <= _T_10366_14;
                                    end else begin
                                      if (_T_17218) begin
                                        _T_18065_60 <= _T_10366_15;
                                      end else begin
                                        if (_T_17216) begin
                                          _T_18065_60 <= _T_10366_16;
                                        end else begin
                                          if (_T_17214) begin
                                            _T_18065_60 <= _T_10366_17;
                                          end else begin
                                            if (_T_17212) begin
                                              _T_18065_60 <= _T_10366_18;
                                            end else begin
                                              if (_T_17210) begin
                                                _T_18065_60 <= _T_10366_19;
                                              end else begin
                                                if (_T_17208) begin
                                                  _T_18065_60 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17206) begin
                                                    _T_18065_60 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17204) begin
                                                      _T_18065_60 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17202) begin
                                                        _T_18065_60 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17200) begin
                                                          _T_18065_60 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17198) begin
                                                            _T_18065_60 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17196) begin
                                                              _T_18065_60 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17194) begin
                                                                _T_18065_60 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17192) begin
                                                                  _T_18065_60 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17190) begin
                                                                    _T_18065_60 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17188) begin
                                                                      _T_18065_60 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17186) begin
                                                                        _T_18065_60 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17184) begin
                                                                          _T_18065_60 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17182) begin
                                                                            _T_18065_60 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17180) begin
                                                                              _T_18065_60 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17178) begin
                                                                                _T_18065_60 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17176) begin
                                                                                  _T_18065_60 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17174) begin
                                                                                    _T_18065_60 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17172) begin
                                                                                      _T_18065_60 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17170) begin
                                                                                        _T_18065_60 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17168) begin
                                                                                          _T_18065_60 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17166) begin
                                                                                            _T_18065_60 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17164) begin
                                                                                              _T_18065_60 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17162) begin
                                                                                                _T_18065_60 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17160) begin
                                                                                                  _T_18065_60 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17158) begin
                                                                                                    _T_18065_60 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17156) begin
                                                                                                      _T_18065_60 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17154) begin
                                                                                                        _T_18065_60 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17152) begin
                                                                                                          _T_18065_60 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17150) begin
                                                                                                            _T_18065_60 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17148) begin
                                                                                                              _T_18065_60 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17146) begin
                                                                                                                _T_18065_60 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17144) begin
                                                                                                                  _T_18065_60 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17142) begin
                                                                                                                    _T_18065_60 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17140) begin
                                                                                                                      _T_18065_60 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17138) begin
                                                                                                                        _T_18065_60 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17136) begin
                                                                                                                          _T_18065_60 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17134) begin
                                                                                                                            _T_18065_60 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17132) begin
                                                                                                                              _T_18065_60 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17130) begin
                                                                                                                                _T_18065_60 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17128) begin
                                                                                                                                  _T_18065_60 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  _T_18065_60 <= 8'h0;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_60 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_61) begin
        if (_T_17435) begin
          _T_18065_61 <= _T_10366_0;
        end else begin
          if (_T_17433) begin
            _T_18065_61 <= _T_10366_1;
          end else begin
            if (_T_17431) begin
              _T_18065_61 <= _T_10366_2;
            end else begin
              if (_T_17429) begin
                _T_18065_61 <= _T_10366_3;
              end else begin
                if (_T_17427) begin
                  _T_18065_61 <= _T_10366_4;
                end else begin
                  if (_T_17425) begin
                    _T_18065_61 <= _T_10366_5;
                  end else begin
                    if (_T_17423) begin
                      _T_18065_61 <= _T_10366_6;
                    end else begin
                      if (_T_17421) begin
                        _T_18065_61 <= _T_10366_7;
                      end else begin
                        if (_T_17419) begin
                          _T_18065_61 <= _T_10366_8;
                        end else begin
                          if (_T_17417) begin
                            _T_18065_61 <= _T_10366_9;
                          end else begin
                            if (_T_17415) begin
                              _T_18065_61 <= _T_10366_10;
                            end else begin
                              if (_T_17413) begin
                                _T_18065_61 <= _T_10366_11;
                              end else begin
                                if (_T_17411) begin
                                  _T_18065_61 <= _T_10366_12;
                                end else begin
                                  if (_T_17409) begin
                                    _T_18065_61 <= _T_10366_13;
                                  end else begin
                                    if (_T_17407) begin
                                      _T_18065_61 <= _T_10366_14;
                                    end else begin
                                      if (_T_17405) begin
                                        _T_18065_61 <= _T_10366_15;
                                      end else begin
                                        if (_T_17403) begin
                                          _T_18065_61 <= _T_10366_16;
                                        end else begin
                                          if (_T_17401) begin
                                            _T_18065_61 <= _T_10366_17;
                                          end else begin
                                            if (_T_17399) begin
                                              _T_18065_61 <= _T_10366_18;
                                            end else begin
                                              if (_T_17397) begin
                                                _T_18065_61 <= _T_10366_19;
                                              end else begin
                                                if (_T_17395) begin
                                                  _T_18065_61 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17393) begin
                                                    _T_18065_61 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17391) begin
                                                      _T_18065_61 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17389) begin
                                                        _T_18065_61 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17387) begin
                                                          _T_18065_61 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17385) begin
                                                            _T_18065_61 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17383) begin
                                                              _T_18065_61 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17381) begin
                                                                _T_18065_61 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17379) begin
                                                                  _T_18065_61 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17377) begin
                                                                    _T_18065_61 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17375) begin
                                                                      _T_18065_61 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17373) begin
                                                                        _T_18065_61 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17371) begin
                                                                          _T_18065_61 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17369) begin
                                                                            _T_18065_61 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17367) begin
                                                                              _T_18065_61 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17365) begin
                                                                                _T_18065_61 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17363) begin
                                                                                  _T_18065_61 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17361) begin
                                                                                    _T_18065_61 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17359) begin
                                                                                      _T_18065_61 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17357) begin
                                                                                        _T_18065_61 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17355) begin
                                                                                          _T_18065_61 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17353) begin
                                                                                            _T_18065_61 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17351) begin
                                                                                              _T_18065_61 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17349) begin
                                                                                                _T_18065_61 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17347) begin
                                                                                                  _T_18065_61 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17345) begin
                                                                                                    _T_18065_61 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17343) begin
                                                                                                      _T_18065_61 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17341) begin
                                                                                                        _T_18065_61 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17339) begin
                                                                                                          _T_18065_61 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17337) begin
                                                                                                            _T_18065_61 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17335) begin
                                                                                                              _T_18065_61 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17333) begin
                                                                                                                _T_18065_61 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17331) begin
                                                                                                                  _T_18065_61 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17329) begin
                                                                                                                    _T_18065_61 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17327) begin
                                                                                                                      _T_18065_61 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17325) begin
                                                                                                                        _T_18065_61 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17323) begin
                                                                                                                          _T_18065_61 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17321) begin
                                                                                                                            _T_18065_61 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17319) begin
                                                                                                                              _T_18065_61 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17317) begin
                                                                                                                                _T_18065_61 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17315) begin
                                                                                                                                  _T_18065_61 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17313) begin
                                                                                                                                    _T_18065_61 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    _T_18065_61 <= 8'h0;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_61 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_62) begin
        if (_T_17625) begin
          _T_18065_62 <= _T_10366_0;
        end else begin
          if (_T_17623) begin
            _T_18065_62 <= _T_10366_1;
          end else begin
            if (_T_17621) begin
              _T_18065_62 <= _T_10366_2;
            end else begin
              if (_T_17619) begin
                _T_18065_62 <= _T_10366_3;
              end else begin
                if (_T_17617) begin
                  _T_18065_62 <= _T_10366_4;
                end else begin
                  if (_T_17615) begin
                    _T_18065_62 <= _T_10366_5;
                  end else begin
                    if (_T_17613) begin
                      _T_18065_62 <= _T_10366_6;
                    end else begin
                      if (_T_17611) begin
                        _T_18065_62 <= _T_10366_7;
                      end else begin
                        if (_T_17609) begin
                          _T_18065_62 <= _T_10366_8;
                        end else begin
                          if (_T_17607) begin
                            _T_18065_62 <= _T_10366_9;
                          end else begin
                            if (_T_17605) begin
                              _T_18065_62 <= _T_10366_10;
                            end else begin
                              if (_T_17603) begin
                                _T_18065_62 <= _T_10366_11;
                              end else begin
                                if (_T_17601) begin
                                  _T_18065_62 <= _T_10366_12;
                                end else begin
                                  if (_T_17599) begin
                                    _T_18065_62 <= _T_10366_13;
                                  end else begin
                                    if (_T_17597) begin
                                      _T_18065_62 <= _T_10366_14;
                                    end else begin
                                      if (_T_17595) begin
                                        _T_18065_62 <= _T_10366_15;
                                      end else begin
                                        if (_T_17593) begin
                                          _T_18065_62 <= _T_10366_16;
                                        end else begin
                                          if (_T_17591) begin
                                            _T_18065_62 <= _T_10366_17;
                                          end else begin
                                            if (_T_17589) begin
                                              _T_18065_62 <= _T_10366_18;
                                            end else begin
                                              if (_T_17587) begin
                                                _T_18065_62 <= _T_10366_19;
                                              end else begin
                                                if (_T_17585) begin
                                                  _T_18065_62 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17583) begin
                                                    _T_18065_62 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17581) begin
                                                      _T_18065_62 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17579) begin
                                                        _T_18065_62 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17577) begin
                                                          _T_18065_62 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17575) begin
                                                            _T_18065_62 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17573) begin
                                                              _T_18065_62 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17571) begin
                                                                _T_18065_62 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17569) begin
                                                                  _T_18065_62 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17567) begin
                                                                    _T_18065_62 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17565) begin
                                                                      _T_18065_62 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17563) begin
                                                                        _T_18065_62 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17561) begin
                                                                          _T_18065_62 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17559) begin
                                                                            _T_18065_62 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17557) begin
                                                                              _T_18065_62 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17555) begin
                                                                                _T_18065_62 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17553) begin
                                                                                  _T_18065_62 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17551) begin
                                                                                    _T_18065_62 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17549) begin
                                                                                      _T_18065_62 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17547) begin
                                                                                        _T_18065_62 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17545) begin
                                                                                          _T_18065_62 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17543) begin
                                                                                            _T_18065_62 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17541) begin
                                                                                              _T_18065_62 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17539) begin
                                                                                                _T_18065_62 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17537) begin
                                                                                                  _T_18065_62 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17535) begin
                                                                                                    _T_18065_62 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17533) begin
                                                                                                      _T_18065_62 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17531) begin
                                                                                                        _T_18065_62 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17529) begin
                                                                                                          _T_18065_62 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17527) begin
                                                                                                            _T_18065_62 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17525) begin
                                                                                                              _T_18065_62 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17523) begin
                                                                                                                _T_18065_62 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17521) begin
                                                                                                                  _T_18065_62 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17519) begin
                                                                                                                    _T_18065_62 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17517) begin
                                                                                                                      _T_18065_62 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17515) begin
                                                                                                                        _T_18065_62 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17513) begin
                                                                                                                          _T_18065_62 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17511) begin
                                                                                                                            _T_18065_62 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17509) begin
                                                                                                                              _T_18065_62 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17507) begin
                                                                                                                                _T_18065_62 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17505) begin
                                                                                                                                  _T_18065_62 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17503) begin
                                                                                                                                    _T_18065_62 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_17501) begin
                                                                                                                                      _T_18065_62 <= _T_10366_62;
                                                                                                                                    end else begin
                                                                                                                                      _T_18065_62 <= 8'h0;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_62 <= 8'h0;
      end
    end
    if (_T_10362) begin
      if (_T_10436_63) begin
        if (_T_17818) begin
          _T_18065_63 <= _T_10366_0;
        end else begin
          if (_T_17816) begin
            _T_18065_63 <= _T_10366_1;
          end else begin
            if (_T_17814) begin
              _T_18065_63 <= _T_10366_2;
            end else begin
              if (_T_17812) begin
                _T_18065_63 <= _T_10366_3;
              end else begin
                if (_T_17810) begin
                  _T_18065_63 <= _T_10366_4;
                end else begin
                  if (_T_17808) begin
                    _T_18065_63 <= _T_10366_5;
                  end else begin
                    if (_T_17806) begin
                      _T_18065_63 <= _T_10366_6;
                    end else begin
                      if (_T_17804) begin
                        _T_18065_63 <= _T_10366_7;
                      end else begin
                        if (_T_17802) begin
                          _T_18065_63 <= _T_10366_8;
                        end else begin
                          if (_T_17800) begin
                            _T_18065_63 <= _T_10366_9;
                          end else begin
                            if (_T_17798) begin
                              _T_18065_63 <= _T_10366_10;
                            end else begin
                              if (_T_17796) begin
                                _T_18065_63 <= _T_10366_11;
                              end else begin
                                if (_T_17794) begin
                                  _T_18065_63 <= _T_10366_12;
                                end else begin
                                  if (_T_17792) begin
                                    _T_18065_63 <= _T_10366_13;
                                  end else begin
                                    if (_T_17790) begin
                                      _T_18065_63 <= _T_10366_14;
                                    end else begin
                                      if (_T_17788) begin
                                        _T_18065_63 <= _T_10366_15;
                                      end else begin
                                        if (_T_17786) begin
                                          _T_18065_63 <= _T_10366_16;
                                        end else begin
                                          if (_T_17784) begin
                                            _T_18065_63 <= _T_10366_17;
                                          end else begin
                                            if (_T_17782) begin
                                              _T_18065_63 <= _T_10366_18;
                                            end else begin
                                              if (_T_17780) begin
                                                _T_18065_63 <= _T_10366_19;
                                              end else begin
                                                if (_T_17778) begin
                                                  _T_18065_63 <= _T_10366_20;
                                                end else begin
                                                  if (_T_17776) begin
                                                    _T_18065_63 <= _T_10366_21;
                                                  end else begin
                                                    if (_T_17774) begin
                                                      _T_18065_63 <= _T_10366_22;
                                                    end else begin
                                                      if (_T_17772) begin
                                                        _T_18065_63 <= _T_10366_23;
                                                      end else begin
                                                        if (_T_17770) begin
                                                          _T_18065_63 <= _T_10366_24;
                                                        end else begin
                                                          if (_T_17768) begin
                                                            _T_18065_63 <= _T_10366_25;
                                                          end else begin
                                                            if (_T_17766) begin
                                                              _T_18065_63 <= _T_10366_26;
                                                            end else begin
                                                              if (_T_17764) begin
                                                                _T_18065_63 <= _T_10366_27;
                                                              end else begin
                                                                if (_T_17762) begin
                                                                  _T_18065_63 <= _T_10366_28;
                                                                end else begin
                                                                  if (_T_17760) begin
                                                                    _T_18065_63 <= _T_10366_29;
                                                                  end else begin
                                                                    if (_T_17758) begin
                                                                      _T_18065_63 <= _T_10366_30;
                                                                    end else begin
                                                                      if (_T_17756) begin
                                                                        _T_18065_63 <= _T_10366_31;
                                                                      end else begin
                                                                        if (_T_17754) begin
                                                                          _T_18065_63 <= _T_10366_32;
                                                                        end else begin
                                                                          if (_T_17752) begin
                                                                            _T_18065_63 <= _T_10366_33;
                                                                          end else begin
                                                                            if (_T_17750) begin
                                                                              _T_18065_63 <= _T_10366_34;
                                                                            end else begin
                                                                              if (_T_17748) begin
                                                                                _T_18065_63 <= _T_10366_35;
                                                                              end else begin
                                                                                if (_T_17746) begin
                                                                                  _T_18065_63 <= _T_10366_36;
                                                                                end else begin
                                                                                  if (_T_17744) begin
                                                                                    _T_18065_63 <= _T_10366_37;
                                                                                  end else begin
                                                                                    if (_T_17742) begin
                                                                                      _T_18065_63 <= _T_10366_38;
                                                                                    end else begin
                                                                                      if (_T_17740) begin
                                                                                        _T_18065_63 <= _T_10366_39;
                                                                                      end else begin
                                                                                        if (_T_17738) begin
                                                                                          _T_18065_63 <= _T_10366_40;
                                                                                        end else begin
                                                                                          if (_T_17736) begin
                                                                                            _T_18065_63 <= _T_10366_41;
                                                                                          end else begin
                                                                                            if (_T_17734) begin
                                                                                              _T_18065_63 <= _T_10366_42;
                                                                                            end else begin
                                                                                              if (_T_17732) begin
                                                                                                _T_18065_63 <= _T_10366_43;
                                                                                              end else begin
                                                                                                if (_T_17730) begin
                                                                                                  _T_18065_63 <= _T_10366_44;
                                                                                                end else begin
                                                                                                  if (_T_17728) begin
                                                                                                    _T_18065_63 <= _T_10366_45;
                                                                                                  end else begin
                                                                                                    if (_T_17726) begin
                                                                                                      _T_18065_63 <= _T_10366_46;
                                                                                                    end else begin
                                                                                                      if (_T_17724) begin
                                                                                                        _T_18065_63 <= _T_10366_47;
                                                                                                      end else begin
                                                                                                        if (_T_17722) begin
                                                                                                          _T_18065_63 <= _T_10366_48;
                                                                                                        end else begin
                                                                                                          if (_T_17720) begin
                                                                                                            _T_18065_63 <= _T_10366_49;
                                                                                                          end else begin
                                                                                                            if (_T_17718) begin
                                                                                                              _T_18065_63 <= _T_10366_50;
                                                                                                            end else begin
                                                                                                              if (_T_17716) begin
                                                                                                                _T_18065_63 <= _T_10366_51;
                                                                                                              end else begin
                                                                                                                if (_T_17714) begin
                                                                                                                  _T_18065_63 <= _T_10366_52;
                                                                                                                end else begin
                                                                                                                  if (_T_17712) begin
                                                                                                                    _T_18065_63 <= _T_10366_53;
                                                                                                                  end else begin
                                                                                                                    if (_T_17710) begin
                                                                                                                      _T_18065_63 <= _T_10366_54;
                                                                                                                    end else begin
                                                                                                                      if (_T_17708) begin
                                                                                                                        _T_18065_63 <= _T_10366_55;
                                                                                                                      end else begin
                                                                                                                        if (_T_17706) begin
                                                                                                                          _T_18065_63 <= _T_10366_56;
                                                                                                                        end else begin
                                                                                                                          if (_T_17704) begin
                                                                                                                            _T_18065_63 <= _T_10366_57;
                                                                                                                          end else begin
                                                                                                                            if (_T_17702) begin
                                                                                                                              _T_18065_63 <= _T_10366_58;
                                                                                                                            end else begin
                                                                                                                              if (_T_17700) begin
                                                                                                                                _T_18065_63 <= _T_10366_59;
                                                                                                                              end else begin
                                                                                                                                if (_T_17698) begin
                                                                                                                                  _T_18065_63 <= _T_10366_60;
                                                                                                                                end else begin
                                                                                                                                  if (_T_17696) begin
                                                                                                                                    _T_18065_63 <= _T_10366_61;
                                                                                                                                  end else begin
                                                                                                                                    if (_T_17694) begin
                                                                                                                                      _T_18065_63 <= _T_10366_62;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_17692) begin
                                                                                                                                        _T_18065_63 <= _T_10366_63;
                                                                                                                                      end else begin
                                                                                                                                        _T_18065_63 <= 8'h0;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        _T_18065_63 <= 8'h0;
      end
    end
    if (reset) begin
      _T_18396 <= 1'h0;
    end else begin
      _T_18396 <= _T_17822;
    end
    if (_T_17822) begin
      _T_18400_0 <= _T_18267;
    end
    if (_T_17822) begin
      _T_18400_1 <= _T_18269;
    end
    if (_T_17822) begin
      _T_18400_2 <= _T_18271;
    end
    if (_T_17822) begin
      _T_18400_3 <= _T_18273;
    end
    if (_T_17822) begin
      _T_18400_4 <= _T_18275;
    end
    if (_T_17822) begin
      _T_18400_5 <= _T_18277;
    end
    if (_T_17822) begin
      _T_18400_6 <= _T_18279;
    end
    if (_T_17822) begin
      _T_18400_7 <= _T_18281;
    end
    if (_T_17822) begin
      _T_18400_8 <= _T_18283;
    end
    if (_T_17822) begin
      _T_18400_9 <= _T_18285;
    end
    if (_T_17822) begin
      _T_18400_10 <= _T_18287;
    end
    if (_T_17822) begin
      _T_18400_11 <= _T_18289;
    end
    if (_T_17822) begin
      _T_18400_12 <= _T_18291;
    end
    if (_T_17822) begin
      _T_18400_13 <= _T_18293;
    end
    if (_T_17822) begin
      _T_18400_14 <= _T_18295;
    end
    if (_T_17822) begin
      _T_18400_15 <= _T_18297;
    end
    if (_T_17822) begin
      _T_18400_16 <= _T_18299;
    end
    if (_T_17822) begin
      _T_18400_17 <= _T_18301;
    end
    if (_T_17822) begin
      _T_18400_18 <= _T_18303;
    end
    if (_T_17822) begin
      _T_18400_19 <= _T_18305;
    end
    if (_T_17822) begin
      _T_18400_20 <= _T_18307;
    end
    if (_T_17822) begin
      _T_18400_21 <= _T_18309;
    end
    if (_T_17822) begin
      _T_18400_22 <= _T_18311;
    end
    if (_T_17822) begin
      _T_18400_23 <= _T_18313;
    end
    if (_T_17822) begin
      _T_18400_24 <= _T_18315;
    end
    if (_T_17822) begin
      _T_18400_25 <= _T_18317;
    end
    if (_T_17822) begin
      _T_18400_26 <= _T_18319;
    end
    if (_T_17822) begin
      _T_18400_27 <= _T_18321;
    end
    if (_T_17822) begin
      _T_18400_28 <= _T_18323;
    end
    if (_T_17822) begin
      _T_18400_29 <= _T_18325;
    end
    if (_T_17822) begin
      _T_18400_30 <= _T_18327;
    end
    if (_T_17822) begin
      _T_18400_31 <= _T_18329;
    end
    if (_T_17822) begin
      _T_18400_32 <= _T_18331;
    end
    if (_T_17822) begin
      _T_18400_33 <= _T_18333;
    end
    if (_T_17822) begin
      _T_18400_34 <= _T_18335;
    end
    if (_T_17822) begin
      _T_18400_35 <= _T_18337;
    end
    if (_T_17822) begin
      _T_18400_36 <= _T_18339;
    end
    if (_T_17822) begin
      _T_18400_37 <= _T_18341;
    end
    if (_T_17822) begin
      _T_18400_38 <= _T_18343;
    end
    if (_T_17822) begin
      _T_18400_39 <= _T_18345;
    end
    if (_T_17822) begin
      _T_18400_40 <= _T_18347;
    end
    if (_T_17822) begin
      _T_18400_41 <= _T_18349;
    end
    if (_T_17822) begin
      _T_18400_42 <= _T_18351;
    end
    if (_T_17822) begin
      _T_18400_43 <= _T_18353;
    end
    if (_T_17822) begin
      _T_18400_44 <= _T_18355;
    end
    if (_T_17822) begin
      _T_18400_45 <= _T_18357;
    end
    if (_T_17822) begin
      _T_18400_46 <= _T_18359;
    end
    if (_T_17822) begin
      _T_18400_47 <= _T_18361;
    end
    if (_T_17822) begin
      _T_18400_48 <= _T_18363;
    end
    if (_T_17822) begin
      _T_18400_49 <= _T_18365;
    end
    if (_T_17822) begin
      _T_18400_50 <= _T_18367;
    end
    if (_T_17822) begin
      _T_18400_51 <= _T_18369;
    end
    if (_T_17822) begin
      _T_18400_52 <= _T_18371;
    end
    if (_T_17822) begin
      _T_18400_53 <= _T_18373;
    end
    if (_T_17822) begin
      _T_18400_54 <= _T_18375;
    end
    if (_T_17822) begin
      _T_18400_55 <= _T_18377;
    end
    if (_T_17822) begin
      _T_18400_56 <= _T_18379;
    end
    if (_T_17822) begin
      _T_18400_57 <= _T_18381;
    end
    if (_T_17822) begin
      _T_18400_58 <= _T_18383;
    end
    if (_T_17822) begin
      _T_18400_59 <= _T_18385;
    end
    if (_T_17822) begin
      _T_18400_60 <= _T_18387;
    end
    if (_T_17822) begin
      _T_18400_61 <= _T_18389;
    end
    if (_T_17822) begin
      _T_18400_62 <= _T_18391;
    end
    if (_T_17822) begin
      _T_18400_63 <= _T_18393;
    end
    if (reset) begin
      _T_18605_0 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_0 <= _T_17961_0;
      end
    end
    if (reset) begin
      _T_18605_1 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_1 <= _T_17961_1;
      end
    end
    if (reset) begin
      _T_18605_2 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_2 <= _T_17961_2;
      end
    end
    if (reset) begin
      _T_18605_3 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_3 <= _T_17961_3;
      end
    end
    if (reset) begin
      _T_18605_4 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_4 <= _T_17961_4;
      end
    end
    if (reset) begin
      _T_18605_5 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_5 <= _T_17961_5;
      end
    end
    if (reset) begin
      _T_18605_6 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_6 <= _T_17961_6;
      end
    end
    if (reset) begin
      _T_18605_7 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_7 <= _T_17961_7;
      end
    end
    if (reset) begin
      _T_18605_8 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_8 <= _T_17961_8;
      end
    end
    if (reset) begin
      _T_18605_9 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_9 <= _T_17961_9;
      end
    end
    if (reset) begin
      _T_18605_10 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_10 <= _T_17961_10;
      end
    end
    if (reset) begin
      _T_18605_11 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_11 <= _T_17961_11;
      end
    end
    if (reset) begin
      _T_18605_12 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_12 <= _T_17961_12;
      end
    end
    if (reset) begin
      _T_18605_13 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_13 <= _T_17961_13;
      end
    end
    if (reset) begin
      _T_18605_14 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_14 <= _T_17961_14;
      end
    end
    if (reset) begin
      _T_18605_15 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_15 <= _T_17961_15;
      end
    end
    if (reset) begin
      _T_18605_16 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_16 <= _T_17961_16;
      end
    end
    if (reset) begin
      _T_18605_17 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_17 <= _T_17961_17;
      end
    end
    if (reset) begin
      _T_18605_18 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_18 <= _T_17961_18;
      end
    end
    if (reset) begin
      _T_18605_19 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_19 <= _T_17961_19;
      end
    end
    if (reset) begin
      _T_18605_20 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_20 <= _T_17961_20;
      end
    end
    if (reset) begin
      _T_18605_21 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_21 <= _T_17961_21;
      end
    end
    if (reset) begin
      _T_18605_22 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_22 <= _T_17961_22;
      end
    end
    if (reset) begin
      _T_18605_23 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_23 <= _T_17961_23;
      end
    end
    if (reset) begin
      _T_18605_24 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_24 <= _T_17961_24;
      end
    end
    if (reset) begin
      _T_18605_25 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_25 <= _T_17961_25;
      end
    end
    if (reset) begin
      _T_18605_26 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_26 <= _T_17961_26;
      end
    end
    if (reset) begin
      _T_18605_27 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_27 <= _T_17961_27;
      end
    end
    if (reset) begin
      _T_18605_28 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_28 <= _T_17961_28;
      end
    end
    if (reset) begin
      _T_18605_29 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_29 <= _T_17961_29;
      end
    end
    if (reset) begin
      _T_18605_30 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_30 <= _T_17961_30;
      end
    end
    if (reset) begin
      _T_18605_31 <= 1'h0;
    end else begin
      if (_T_17822) begin
        _T_18605_31 <= _T_17961_31;
      end
    end
    if (_T_17822) begin
      _T_18709_0 <= _T_18065_0;
    end
    if (_T_17822) begin
      _T_18709_1 <= _T_18065_1;
    end
    if (_T_17822) begin
      _T_18709_2 <= _T_18065_2;
    end
    if (_T_17822) begin
      _T_18709_3 <= _T_18065_3;
    end
    if (_T_17822) begin
      _T_18709_4 <= _T_18065_4;
    end
    if (_T_17822) begin
      _T_18709_5 <= _T_18065_5;
    end
    if (_T_17822) begin
      _T_18709_6 <= _T_18065_6;
    end
    if (_T_17822) begin
      _T_18709_7 <= _T_18065_7;
    end
    if (_T_17822) begin
      _T_18709_8 <= _T_18065_8;
    end
    if (_T_17822) begin
      _T_18709_9 <= _T_18065_9;
    end
    if (_T_17822) begin
      _T_18709_10 <= _T_18065_10;
    end
    if (_T_17822) begin
      _T_18709_11 <= _T_18065_11;
    end
    if (_T_17822) begin
      _T_18709_12 <= _T_18065_12;
    end
    if (_T_17822) begin
      _T_18709_13 <= _T_18065_13;
    end
    if (_T_17822) begin
      _T_18709_14 <= _T_18065_14;
    end
    if (_T_17822) begin
      _T_18709_15 <= _T_18065_15;
    end
    if (_T_17822) begin
      _T_18709_16 <= _T_18065_16;
    end
    if (_T_17822) begin
      _T_18709_17 <= _T_18065_17;
    end
    if (_T_17822) begin
      _T_18709_18 <= _T_18065_18;
    end
    if (_T_17822) begin
      _T_18709_19 <= _T_18065_19;
    end
    if (_T_17822) begin
      _T_18709_20 <= _T_18065_20;
    end
    if (_T_17822) begin
      _T_18709_21 <= _T_18065_21;
    end
    if (_T_17822) begin
      _T_18709_22 <= _T_18065_22;
    end
    if (_T_17822) begin
      _T_18709_23 <= _T_18065_23;
    end
    if (_T_17822) begin
      _T_18709_24 <= _T_18065_24;
    end
    if (_T_17822) begin
      _T_18709_25 <= _T_18065_25;
    end
    if (_T_17822) begin
      _T_18709_26 <= _T_18065_26;
    end
    if (_T_17822) begin
      _T_18709_27 <= _T_18065_27;
    end
    if (_T_17822) begin
      _T_18709_28 <= _T_18065_28;
    end
    if (_T_17822) begin
      _T_18709_29 <= _T_18065_29;
    end
    if (_T_17822) begin
      _T_18709_30 <= _T_18065_30;
    end
    if (_T_17822) begin
      _T_18709_31 <= _T_18065_31;
    end
    if (_T_17822) begin
      _T_18709_32 <= _T_18065_32;
    end
    if (_T_17822) begin
      _T_18709_33 <= _T_18065_33;
    end
    if (_T_17822) begin
      _T_18709_34 <= _T_18065_34;
    end
    if (_T_17822) begin
      _T_18709_35 <= _T_18065_35;
    end
    if (_T_17822) begin
      _T_18709_36 <= _T_18065_36;
    end
    if (_T_17822) begin
      _T_18709_37 <= _T_18065_37;
    end
    if (_T_17822) begin
      _T_18709_38 <= _T_18065_38;
    end
    if (_T_17822) begin
      _T_18709_39 <= _T_18065_39;
    end
    if (_T_17822) begin
      _T_18709_40 <= _T_18065_40;
    end
    if (_T_17822) begin
      _T_18709_41 <= _T_18065_41;
    end
    if (_T_17822) begin
      _T_18709_42 <= _T_18065_42;
    end
    if (_T_17822) begin
      _T_18709_43 <= _T_18065_43;
    end
    if (_T_17822) begin
      _T_18709_44 <= _T_18065_44;
    end
    if (_T_17822) begin
      _T_18709_45 <= _T_18065_45;
    end
    if (_T_17822) begin
      _T_18709_46 <= _T_18065_46;
    end
    if (_T_17822) begin
      _T_18709_47 <= _T_18065_47;
    end
    if (_T_17822) begin
      _T_18709_48 <= _T_18065_48;
    end
    if (_T_17822) begin
      _T_18709_49 <= _T_18065_49;
    end
    if (_T_17822) begin
      _T_18709_50 <= _T_18065_50;
    end
    if (_T_17822) begin
      _T_18709_51 <= _T_18065_51;
    end
    if (_T_17822) begin
      _T_18709_52 <= _T_18065_52;
    end
    if (_T_17822) begin
      _T_18709_53 <= _T_18065_53;
    end
    if (_T_17822) begin
      _T_18709_54 <= _T_18065_54;
    end
    if (_T_17822) begin
      _T_18709_55 <= _T_18065_55;
    end
    if (_T_17822) begin
      _T_18709_56 <= _T_18065_56;
    end
    if (_T_17822) begin
      _T_18709_57 <= _T_18065_57;
    end
    if (_T_17822) begin
      _T_18709_58 <= _T_18065_58;
    end
    if (_T_17822) begin
      _T_18709_59 <= _T_18065_59;
    end
    if (_T_17822) begin
      _T_18709_60 <= _T_18065_60;
    end
    if (_T_17822) begin
      _T_18709_61 <= _T_18065_61;
    end
    if (_T_17822) begin
      _T_18709_62 <= _T_18065_62;
    end
    if (_T_17822) begin
      _T_18709_63 <= _T_18065_63;
    end
  end
endmodule
module NV_soDLA_CSC_wl( // @[:@14280.2]
  input          clock, // @[:@14281.4]
  input          reset, // @[:@14282.4]
  input          io_nvdla_core_clk, // @[:@14283.4]
  input          io_nvdla_core_ng_clk, // @[:@14283.4]
  input          io_sg2wl_pd_valid, // @[:@14283.4]
  input  [17:0]  io_sg2wl_pd_bits, // @[:@14283.4]
  input          io_sg2wl_reuse_rls, // @[:@14283.4]
  input  [1:0]   io_sc_state, // @[:@14283.4]
  input          io_sc2cdma_wt_pending_req, // @[:@14283.4]
  input          io_cdma2sc_wt_updt_valid, // @[:@14283.4]
  input  [14:0]  io_cdma2sc_wt_updt_bits_entries, // @[:@14283.4]
  input  [13:0]  io_cdma2sc_wt_updt_bits_kernels, // @[:@14283.4]
  input  [8:0]   io_cdma2sc_wmb_entries, // @[:@14283.4]
  output         io_sc2cdma_wt_updt_valid, // @[:@14283.4]
  output [14:0]  io_sc2cdma_wt_updt_bits_entries, // @[:@14283.4]
  output [13:0]  io_sc2cdma_wt_updt_bits_kernels, // @[:@14283.4]
  output [8:0]   io_sc2cdma_wmb_entries, // @[:@14283.4]
  output         io_sc2buf_wt_rd_addr_valid, // @[:@14283.4]
  output [12:0]  io_sc2buf_wt_rd_addr_bits, // @[:@14283.4]
  input          io_sc2buf_wt_rd_data_valid, // @[:@14283.4]
  input  [511:0] io_sc2buf_wt_rd_data_bits, // @[:@14283.4]
  output         io_sc2mac_wt_a_valid, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_0, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_1, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_2, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_3, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_4, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_5, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_6, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_7, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_8, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_9, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_10, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_11, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_12, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_13, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_14, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_sel_15, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_0, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_1, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_2, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_3, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_4, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_5, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_6, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_7, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_8, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_9, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_10, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_11, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_12, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_13, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_14, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_15, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_16, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_17, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_18, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_19, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_20, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_21, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_22, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_23, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_24, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_25, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_26, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_27, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_28, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_29, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_30, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_31, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_32, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_33, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_34, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_35, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_36, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_37, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_38, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_39, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_40, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_41, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_42, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_43, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_44, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_45, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_46, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_47, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_48, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_49, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_50, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_51, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_52, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_53, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_54, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_55, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_56, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_57, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_58, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_59, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_60, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_61, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_62, // @[:@14283.4]
  output         io_sc2mac_wt_a_bits_mask_63, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_0, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_1, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_2, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_3, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_4, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_5, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_6, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_7, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_8, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_9, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_10, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_11, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_12, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_13, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_14, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_15, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_16, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_17, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_18, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_19, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_20, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_21, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_22, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_23, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_24, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_25, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_26, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_27, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_28, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_29, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_30, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_31, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_32, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_33, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_34, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_35, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_36, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_37, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_38, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_39, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_40, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_41, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_42, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_43, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_44, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_45, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_46, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_47, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_48, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_49, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_50, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_51, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_52, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_53, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_54, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_55, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_56, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_57, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_58, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_59, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_60, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_61, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_62, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_a_bits_data_63, // @[:@14283.4]
  output         io_sc2mac_wt_b_valid, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_0, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_1, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_2, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_3, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_4, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_5, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_6, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_7, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_8, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_9, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_10, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_11, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_12, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_13, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_14, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_sel_15, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_0, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_1, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_2, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_3, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_4, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_5, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_6, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_7, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_8, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_9, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_10, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_11, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_12, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_13, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_14, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_15, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_16, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_17, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_18, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_19, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_20, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_21, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_22, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_23, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_24, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_25, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_26, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_27, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_28, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_29, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_30, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_31, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_32, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_33, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_34, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_35, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_36, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_37, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_38, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_39, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_40, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_41, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_42, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_43, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_44, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_45, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_46, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_47, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_48, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_49, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_50, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_51, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_52, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_53, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_54, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_55, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_56, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_57, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_58, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_59, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_60, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_61, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_62, // @[:@14283.4]
  output         io_sc2mac_wt_b_bits_mask_63, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_0, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_1, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_2, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_3, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_4, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_5, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_6, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_7, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_8, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_9, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_10, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_11, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_12, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_13, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_14, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_15, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_16, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_17, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_18, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_19, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_20, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_21, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_22, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_23, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_24, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_25, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_26, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_27, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_28, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_29, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_30, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_31, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_32, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_33, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_34, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_35, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_36, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_37, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_38, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_39, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_40, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_41, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_42, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_43, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_44, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_45, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_46, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_47, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_48, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_49, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_50, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_51, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_52, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_53, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_54, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_55, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_56, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_57, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_58, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_59, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_60, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_61, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_62, // @[:@14283.4]
  output [7:0]   io_sc2mac_wt_b_bits_data_63, // @[:@14283.4]
  input          io_reg2dp_op_en, // @[:@14283.4]
  input  [1:0]   io_reg2dp_in_precision, // @[:@14283.4]
  input  [1:0]   io_reg2dp_proc_precision, // @[:@14283.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@14283.4]
  input          io_reg2dp_weight_reuse, // @[:@14283.4]
  input          io_reg2dp_skip_weight_rls, // @[:@14283.4]
  input          io_reg2dp_weight_format, // @[:@14283.4]
  input  [31:0]  io_reg2dp_weight_bytes, // @[:@14283.4]
  input  [27:0]  io_reg2dp_wmb_bytes, // @[:@14283.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@14283.4]
  input  [4:0]   io_reg2dp_weight_bank // @[:@14283.4]
);
  wire  NV_NVDLA_CSC_WL_dec_reset; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_valid; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_input_bits_data_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [9:0] NV_NVDLA_CSC_WL_dec_io_input_mask_en; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_valid; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_32; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_33; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_34; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_35; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_36; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_37; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_38; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_39; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_40; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_41; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_42; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_43; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_44; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_45; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_46; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_47; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_48; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_49; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_50; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_51; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_52; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_53; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_54; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_55; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_56; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_57; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_58; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_59; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_60; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_61; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_62; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire [7:0] NV_NVDLA_CSC_WL_dec_io_output_bits_data_63; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  wire  NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31; // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
  reg  _T_698; // @[NV_NVDLA_CSC_wl.scala 95:35:@14286.4]
  reg [31:0] _RAND_0;
  wire  _T_700; // @[NV_NVDLA_CSC_wl.scala 97:35:@14287.4]
  wire  _T_704; // @[NV_NVDLA_CSC_wl.scala 99:38:@14289.4]
  wire  _T_706; // @[NV_NVDLA_CSC_wl.scala 100:35:@14290.4]
  wire  _T_707; // @[NV_NVDLA_CSC_wl.scala 101:37:@14291.4]
  wire  _T_708; // @[NV_NVDLA_CSC_wl.scala 101:35:@14292.4]
  reg [4:0] _T_715; // @[NV_NVDLA_CSC_wl.scala 108:28:@14295.4]
  reg [31:0] _RAND_1;
  reg [4:0] _T_722; // @[NV_NVDLA_CSC_wl.scala 109:30:@14297.4]
  reg [31:0] _RAND_2;
  reg [14:0] _T_729; // @[NV_NVDLA_CSC_wl.scala 110:38:@14299.4]
  reg [31:0] _RAND_3;
  reg [8:0] _T_736; // @[NV_NVDLA_CSC_wl.scala 111:35:@14301.4]
  reg [31:0] _RAND_4;
  reg [2:0] _T_739; // @[NV_NVDLA_CSC_wl.scala 112:30:@14302.4]
  reg [31:0] _RAND_5;
  reg  _T_742; // @[NV_NVDLA_CSC_wl.scala 113:35:@14303.4]
  reg [31:0] _RAND_6;
  wire  _T_743; // @[NV_NVDLA_CSC_wl.scala 115:36:@14304.4]
  wire [5:0] _T_749; // @[NV_NVDLA_CSC_wl.scala 120:42:@14308.6]
  wire [4:0] _T_750; // @[NV_NVDLA_CSC_wl.scala 120:42:@14309.6]
  wire [5:0] _T_752; // @[NV_NVDLA_CSC_wl.scala 121:46:@14311.6]
  wire [4:0] _T_753; // @[NV_NVDLA_CSC_wl.scala 121:46:@14312.6]
  wire [8:0] _T_755; // @[NV_NVDLA_CSC_wl.scala 122:42:@14314.6]
  wire [2:0] _T_756; // @[NV_NVDLA_CSC_wl.scala 122:67:@14315.6]
  wire [4:0] _GEN_0; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  wire [4:0] _GEN_1; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  wire [2:0] _GEN_2; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  wire  _GEN_3; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  wire  _T_757; // @[NV_NVDLA_CSC_wl.scala 125:21:@14319.4]
  wire [14:0] _T_758; // @[NV_NVDLA_CSC_wl.scala 126:54:@14321.6]
  wire [8:0] _T_759; // @[NV_NVDLA_CSC_wl.scala 127:70:@14323.6]
  wire [8:0] _T_761; // @[NV_NVDLA_CSC_wl.scala 127:32:@14324.6]
  wire [14:0] _GEN_4; // @[NV_NVDLA_CSC_wl.scala 125:49:@14320.4]
  wire [8:0] _GEN_5; // @[NV_NVDLA_CSC_wl.scala 125:49:@14320.4]
  reg  _T_1692; // @[NV_NVDLA_CSC_wl.scala 654:76:@15119.4]
  reg [31:0] _RAND_7;
  reg [35:0] _T_1712; // @[NV_NVDLA_CSC_wl.scala 656:75:@15126.4]
  reg [63:0] _RAND_8;
  wire  _T_1759; // @[NV_NVDLA_CSC_wl.scala 693:34:@15202.4]
  wire  _T_857; // @[NV_NVDLA_CSC_wl.scala 203:36:@14402.4]
  wire  _T_858; // @[NV_NVDLA_CSC_wl.scala 207:25:@14403.4]
  wire [14:0] _T_1755; // @[NV_NVDLA_CSC_wl.scala 689:44:@15197.4]
  wire [14:0] _T_859; // @[NV_NVDLA_CSC_wl.scala 208:29:@14405.4]
  wire [8:0] _T_1754; // @[NV_NVDLA_CSC_wl.scala 688:45:@15195.4]
  wire [8:0] _T_860; // @[NV_NVDLA_CSC_wl.scala 209:30:@14407.4]
  reg [14:0] _T_798; // @[NV_NVDLA_CSC_wl.scala 153:62:@14348.4]
  reg [31:0] _RAND_9;
  wire [15:0] _T_799; // @[NV_NVDLA_CSC_wl.scala 155:39:@14349.4]
  wire [14:0] _T_800; // @[NV_NVDLA_CSC_wl.scala 155:39:@14350.4]
  wire [13:0] _T_802; // @[Cat.scala 30:58:@14351.4]
  wire [14:0] _GEN_497; // @[NV_NVDLA_CSC_wl.scala 156:48:@14352.4]
  wire [15:0] _T_803; // @[NV_NVDLA_CSC_wl.scala 156:48:@14352.4]
  wire [15:0] _T_804; // @[NV_NVDLA_CSC_wl.scala 156:48:@14353.4]
  wire [14:0] _T_805; // @[NV_NVDLA_CSC_wl.scala 156:48:@14354.4]
  wire  _T_808; // @[NV_NVDLA_CSC_wl.scala 157:48:@14356.4]
  wire  _T_810; // @[NV_NVDLA_CSC_wl.scala 158:88:@14357.4]
  wire [14:0] _T_811; // @[NV_NVDLA_CSC_wl.scala 158:113:@14358.4]
  wire [14:0] _T_812; // @[NV_NVDLA_CSC_wl.scala 158:87:@14359.4]
  wire [14:0] _T_813; // @[NV_NVDLA_CSC_wl.scala 158:28:@14360.4]
  wire  _T_847; // @[NV_NVDLA_CSC_wl.scala 184:21:@14388.4]
  wire [14:0] _GEN_8; // @[NV_NVDLA_CSC_wl.scala 184:30:@14389.4]
  reg  _T_863; // @[NV_NVDLA_CSC_wl.scala 212:40:@14409.4]
  reg [31:0] _RAND_10;
  reg [14:0] _T_867; // @[Reg.scala 19:20:@14413.4]
  reg [31:0] _RAND_11;
  wire [14:0] _GEN_12; // @[Reg.scala 20:19:@14414.4]
  reg [8:0] _T_871; // @[Reg.scala 19:20:@14419.4]
  reg [31:0] _RAND_12;
  wire [8:0] _GEN_13; // @[Reg.scala 20:19:@14420.4]
  reg  _T_877; // @[NV_NVDLA_CSC_wl.scala 223:71:@14426.4]
  reg [31:0] _RAND_13;
  reg [17:0] _T_882; // @[NV_NVDLA_CSC_wl.scala 225:67:@14428.4]
  reg [31:0] _RAND_14;
  wire  _T_879; // @[NV_NVDLA_CSC_wl.scala 224:26:@14427.4 NV_NVDLA_CSC_wl.scala 228:19:@14430.4]
  wire [17:0] _GEN_14; // @[NV_NVDLA_CSC_wl.scala 232:30:@14432.4]
  wire [6:0] _T_883; // @[NV_NVDLA_CSC_wl.scala 241:31:@14435.4]
  wire [5:0] _T_884; // @[NV_NVDLA_CSC_wl.scala 242:31:@14436.4]
  wire [1:0] _T_885; // @[NV_NVDLA_CSC_wl.scala 243:29:@14437.4]
  wire  _T_886; // @[NV_NVDLA_CSC_wl.scala 244:31:@14438.4]
  wire  _T_887; // @[NV_NVDLA_CSC_wl.scala 245:29:@14439.4]
  wire  _T_888; // @[NV_NVDLA_CSC_wl.scala 246:30:@14440.4]
  reg [4:0] _T_893; // @[NV_NVDLA_CSC_wl.scala 254:29:@14442.4]
  reg [31:0] _RAND_15;
  reg  _T_896; // @[NV_NVDLA_CSC_wl.scala 255:36:@14443.4]
  reg [31:0] _RAND_16;
  wire [5:0] _T_898; // @[NV_NVDLA_CSC_wl.scala 257:37:@14444.4]
  wire [4:0] _T_899; // @[NV_NVDLA_CSC_wl.scala 257:37:@14445.4]
  wire [4:0] _T_904; // @[NV_NVDLA_CSC_wl.scala 259:39:@14448.4]
  wire  _T_905; // @[NV_NVDLA_CSC_wl.scala 260:38:@14449.4]
  wire [4:0] _T_902; // @[NV_NVDLA_CSC_wl.scala 258:59:@14446.4]
  wire [4:0] _T_903; // @[NV_NVDLA_CSC_wl.scala 258:27:@14447.4]
  wire  _T_908; // @[NV_NVDLA_CSC_wl.scala 262:64:@14451.4]
  wire  _T_909; // @[NV_NVDLA_CSC_wl.scala 262:51:@14452.4]
  wire  _T_911; // @[NV_NVDLA_CSC_wl.scala 262:50:@14453.4]
  wire  _T_912; // @[NV_NVDLA_CSC_wl.scala 262:29:@14454.4]
  wire  _T_913; // @[NV_NVDLA_CSC_wl.scala 263:38:@14455.4]
  wire [4:0] _GEN_15; // @[NV_NVDLA_CSC_wl.scala 265:28:@14456.4]
  reg [10:0] _T_920; // @[NV_NVDLA_CSC_wl.scala 272:34:@14461.4]
  reg [31:0] _RAND_17;
  reg [10:0] _T_923; // @[NV_NVDLA_CSC_wl.scala 273:39:@14462.4]
  reg [31:0] _RAND_18;
  wire  _T_966; // @[NV_NVDLA_CSC_wl.scala 289:37:@14493.4]
  wire  _T_964; // @[Mux.scala 46:19:@14490.4]
  wire [7:0] _T_942; // @[Cat.scala 30:58:@14476.4]
  wire  _T_962; // @[Mux.scala 46:19:@14488.4]
  wire [6:0] _T_951; // @[NV_NVDLA_CSC_wl.scala 285:101:@14480.4]
  wire [8:0] _T_954; // @[Cat.scala 30:58:@14482.4]
  wire  _T_960; // @[Mux.scala 46:19:@14486.4]
  wire [7:0] _T_958; // @[Cat.scala 30:58:@14484.4]
  wire [8:0] _T_959; // @[NV_NVDLA_CSC_wl.scala 286:109:@14485.4]
  wire [5:0] _T_944; // @[NV_NVDLA_CSC_wl.scala 282:92:@14477.4]
  wire [8:0] _T_947; // @[Cat.scala 30:58:@14479.4]
  wire [8:0] _T_961; // @[Mux.scala 46:16:@14487.4]
  wire [8:0] _T_963; // @[Mux.scala 46:16:@14489.4]
  wire [8:0] _T_965; // @[Mux.scala 46:16:@14491.4]
  wire [7:0] _T_917; // @[NV_NVDLA_CSC_wl.scala 271:31:@14460.4 NV_NVDLA_CSC_wl.scala 282:21:@14492.4]
  wire [10:0] _T_968; // @[Cat.scala 30:58:@14494.4]
  wire  _T_969; // @[NV_NVDLA_CSC_wl.scala 289:75:@14495.4]
  wire  _T_970; // @[NV_NVDLA_CSC_wl.scala 289:56:@14496.4]
  wire  _T_924; // @[NV_NVDLA_CSC_wl.scala 275:35:@14463.4]
  wire [10:0] _T_927; // @[NV_NVDLA_CSC_wl.scala 275:34:@14464.4]
  wire [7:0] _T_929; // @[NV_NVDLA_CSC_wl.scala 276:34:@14465.4]
  wire [11:0] _T_930; // @[NV_NVDLA_CSC_wl.scala 277:47:@14466.4]
  wire [10:0] _T_931; // @[NV_NVDLA_CSC_wl.scala 277:47:@14467.4]
  wire [10:0] _GEN_501; // @[NV_NVDLA_CSC_wl.scala 277:69:@14468.4]
  wire [11:0] _T_932; // @[NV_NVDLA_CSC_wl.scala 277:69:@14468.4]
  wire [11:0] _T_933; // @[NV_NVDLA_CSC_wl.scala 277:69:@14469.4]
  wire [10:0] _T_934; // @[NV_NVDLA_CSC_wl.scala 277:69:@14470.4]
  wire  _T_936; // @[NV_NVDLA_CSC_wl.scala 278:82:@14471.4]
  wire  _T_937; // @[NV_NVDLA_CSC_wl.scala 278:80:@14472.4]
  wire  _T_938; // @[NV_NVDLA_CSC_wl.scala 278:96:@14473.4]
  wire [10:0] _T_939; // @[NV_NVDLA_CSC_wl.scala 278:65:@14474.4]
  wire [10:0] _T_940; // @[NV_NVDLA_CSC_wl.scala 278:32:@14475.4]
  wire  _T_972; // @[NV_NVDLA_CSC_wl.scala 290:43:@14499.4]
  wire  _T_974; // @[NV_NVDLA_CSC_wl.scala 291:85:@14501.4]
  wire  _T_975; // @[NV_NVDLA_CSC_wl.scala 291:101:@14502.4]
  wire  _T_976; // @[NV_NVDLA_CSC_wl.scala 291:48:@14503.4]
  wire [10:0] _GEN_16; // @[NV_NVDLA_CSC_wl.scala 293:33:@14504.4]
  wire [10:0] _GEN_17; // @[NV_NVDLA_CSC_wl.scala 296:38:@14507.4]
  reg  _T_1003; // @[NV_NVDLA_CSC_wl.scala 318:34:@14535.4]
  reg [31:0] _RAND_19;
  reg [8:0] _T_1006; // @[NV_NVDLA_CSC_wl.scala 319:30:@14536.4]
  reg [31:0] _RAND_20;
  wire  _T_1007; // @[NV_NVDLA_CSC_wl.scala 321:58:@14537.4]
  wire  _T_1008; // @[NV_NVDLA_CSC_wl.scala 321:42:@14538.4]
  wire  _T_1010; // @[NV_NVDLA_CSC_wl.scala 322:48:@14539.4]
  wire  _T_1012; // @[NV_NVDLA_CSC_wl.scala 322:32:@14540.4]
  wire  _T_1013; // @[NV_NVDLA_CSC_wl.scala 321:32:@14541.4]
  wire [9:0] _T_1015; // @[NV_NVDLA_CSC_wl.scala 323:39:@14542.4]
  wire [8:0] _T_1016; // @[NV_NVDLA_CSC_wl.scala 323:39:@14543.4]
  wire  _T_1018; // @[NV_NVDLA_CSC_wl.scala 325:43:@14544.4]
  wire [8:0] _T_1020; // @[NV_NVDLA_CSC_wl.scala 325:28:@14545.4]
  wire [8:0] _T_1021; // @[NV_NVDLA_CSC_wl.scala 324:28:@14546.4]
  wire  _T_1022; // @[NV_NVDLA_CSC_wl.scala 326:58:@14547.4]
  wire  _T_1023; // @[NV_NVDLA_CSC_wl.scala 326:75:@14548.4]
  wire  _T_1024; // @[NV_NVDLA_CSC_wl.scala 326:91:@14549.4]
  wire  _T_1025; // @[NV_NVDLA_CSC_wl.scala 326:39:@14550.4]
  wire  _T_1026; // @[NV_NVDLA_CSC_wl.scala 326:126:@14551.4]
  wire  _T_1027; // @[NV_NVDLA_CSC_wl.scala 326:144:@14552.4]
  wire  _T_1028; // @[NV_NVDLA_CSC_wl.scala 326:142:@14553.4]
  wire  _T_1029; // @[NV_NVDLA_CSC_wl.scala 326:107:@14554.4]
  wire  _T_1031; // @[NV_NVDLA_CSC_wl.scala 327:47:@14556.4]
  wire [8:0] _T_1032; // @[NV_NVDLA_CSC_wl.scala 327:30:@14557.4]
  wire [8:0] _GEN_20; // @[NV_NVDLA_CSC_wl.scala 330:29:@14559.4]
  reg [6:0] _T_1041; // @[NV_NVDLA_CSC_wl.scala 337:41:@14564.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_1044; // @[NV_NVDLA_CSC_wl.scala 338:37:@14565.4]
  reg [31:0] _RAND_22;
  reg [8:0] _T_1047; // @[NV_NVDLA_CSC_wl.scala 339:41:@14566.4]
  reg [31:0] _RAND_23;
  reg  _T_1050; // @[NV_NVDLA_CSC_wl.scala 340:40:@14567.4]
  reg [31:0] _RAND_24;
  reg  _T_1053; // @[NV_NVDLA_CSC_wl.scala 341:41:@14568.4]
  reg [31:0] _RAND_25;
  reg  _T_1056; // @[NV_NVDLA_CSC_wl.scala 342:39:@14569.4]
  reg [31:0] _RAND_26;
  reg  _T_1059; // @[NV_NVDLA_CSC_wl.scala 343:33:@14570.4]
  reg [31:0] _RAND_27;
  reg [1:0] _T_1062; // @[NV_NVDLA_CSC_wl.scala 344:39:@14571.4]
  reg [31:0] _RAND_28;
  wire [6:0] _GEN_22; // @[NV_NVDLA_CSC_wl.scala 351:25:@14577.4]
  wire [7:0] _GEN_23; // @[NV_NVDLA_CSC_wl.scala 351:25:@14577.4]
  wire  _T_1063; // @[NV_NVDLA_CSC_wl.scala 355:25:@14581.4]
  wire  _T_1064; // @[NV_NVDLA_CSC_wl.scala 355:41:@14582.4]
  wire [8:0] _GEN_24; // @[NV_NVDLA_CSC_wl.scala 355:57:@14583.4]
  wire  _T_1067; // @[NV_NVDLA_CSC_wl.scala 362:41:@14592.6]
  wire  _GEN_25; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  wire  _GEN_26; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  wire  _GEN_27; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  wire  _GEN_28; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  wire [1:0] _GEN_29; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  wire [30:0] _T_1076; // @[Cat.scala 30:58:@14603.4]
  reg  _T_1081; // @[NV_NVDLA_CSC_wl.scala 385:77:@14605.4]
  reg [31:0] _RAND_29;
  reg  _T_1084; // @[NV_NVDLA_CSC_wl.scala 385:77:@14606.4]
  reg [31:0] _RAND_30;
  reg  _T_1087; // @[NV_NVDLA_CSC_wl.scala 385:77:@14607.4]
  reg [31:0] _RAND_31;
  reg  _T_1090; // @[NV_NVDLA_CSC_wl.scala 385:77:@14608.4]
  reg [31:0] _RAND_32;
  reg  _T_1093; // @[NV_NVDLA_CSC_wl.scala 385:77:@14609.4]
  reg [31:0] _RAND_33;
  reg  _T_1096; // @[NV_NVDLA_CSC_wl.scala 385:77:@14610.4]
  reg [31:0] _RAND_34;
  reg [30:0] _T_1101; // @[NV_NVDLA_CSC_wl.scala 387:75:@14612.4]
  reg [31:0] _RAND_35;
  reg [30:0] _T_1104; // @[NV_NVDLA_CSC_wl.scala 387:75:@14613.4]
  reg [31:0] _RAND_36;
  reg [30:0] _T_1107; // @[NV_NVDLA_CSC_wl.scala 387:75:@14614.4]
  reg [31:0] _RAND_37;
  reg [30:0] _T_1110; // @[NV_NVDLA_CSC_wl.scala 387:75:@14615.4]
  reg [31:0] _RAND_38;
  reg [30:0] _T_1113; // @[NV_NVDLA_CSC_wl.scala 387:75:@14616.4]
  reg [31:0] _RAND_39;
  reg [30:0] _T_1116; // @[NV_NVDLA_CSC_wl.scala 387:75:@14617.4]
  reg [31:0] _RAND_40;
  wire [30:0] _GEN_30; // @[NV_NVDLA_CSC_wl.scala 394:37:@14621.4]
  wire [30:0] _GEN_31; // @[NV_NVDLA_CSC_wl.scala 394:37:@14625.4]
  wire [30:0] _GEN_32; // @[NV_NVDLA_CSC_wl.scala 394:37:@14629.4]
  wire [30:0] _GEN_33; // @[NV_NVDLA_CSC_wl.scala 394:37:@14633.4]
  wire [30:0] _GEN_34; // @[NV_NVDLA_CSC_wl.scala 394:37:@14637.4]
  wire [30:0] _GEN_35; // @[NV_NVDLA_CSC_wl.scala 394:37:@14641.4]
  wire [6:0] _T_1117; // @[NV_NVDLA_CSC_wl.scala 404:46:@14644.4]
  wire [7:0] _T_1118; // @[NV_NVDLA_CSC_wl.scala 405:42:@14645.4]
  wire [8:0] _T_1119; // @[NV_NVDLA_CSC_wl.scala 406:46:@14646.4]
  wire  _T_1120; // @[NV_NVDLA_CSC_wl.scala 407:45:@14647.4]
  wire  _T_1121; // @[NV_NVDLA_CSC_wl.scala 408:46:@14648.4]
  wire  _T_1122; // @[NV_NVDLA_CSC_wl.scala 409:44:@14649.4]
  wire  _T_1123; // @[NV_NVDLA_CSC_wl.scala 410:38:@14650.4]
  wire [1:0] _T_1124; // @[NV_NVDLA_CSC_wl.scala 411:44:@14651.4]
  wire  _T_1137; // @[NV_NVDLA_CSC_wl.scala 421:91:@14656.4]
  wire  _T_1138; // @[NV_NVDLA_CSC_wl.scala 421:89:@14657.4]
  wire  _T_1145; // @[NV_NVDLA_CSC_wl.scala 422:72:@14664.4]
  wire  _T_1146; // @[NV_NVDLA_CSC_wl.scala 422:92:@14665.4]
  wire  _T_1147; // @[NV_NVDLA_CSC_wl.scala 422:51:@14666.4]
  wire  _T_1148; // @[NV_NVDLA_CSC_wl.scala 424:40:@14667.4]
  wire  _T_1149; // @[NV_NVDLA_CSC_wl.scala 424:19:@14668.4]
  reg [318:0] _T_1156; // @[NV_NVDLA_CSC_wl.scala 433:31:@14676.4]
  reg [319:0] _RAND_41;
  reg [511:0] _T_1163; // @[NV_NVDLA_CSC_wl.scala 434:35:@14678.4]
  reg [511:0] _RAND_42;
  wire [63:0] _T_1170; // @[NV_NVDLA_CSC_wl.scala 437:63:@14684.4]
  wire [190:0] _T_1171; // @[NV_NVDLA_CSC_wl.scala 437:45:@14685.4]
  wire  _T_1172; // @[NV_NVDLA_CSC_wl.scala 437:108:@14686.4]
  wire [63:0] _T_1176; // @[Bitwise.scala 72:12:@14688.4]
  wire [190:0] _GEN_503; // @[NV_NVDLA_CSC_wl.scala 437:85:@14689.4]
  wire [190:0] _T_1177; // @[NV_NVDLA_CSC_wl.scala 437:85:@14689.4]
  wire [318:0] _T_1183; // @[NV_NVDLA_CSC_wl.scala 438:56:@14691.4]
  wire [318:0] _T_1184; // @[NV_NVDLA_CSC_wl.scala 438:25:@14692.4]
  wire [63:0] _T_1185; // @[NV_NVDLA_CSC_wl.scala 439:41:@14693.4]
  wire [318:0] _GEN_504; // @[NV_NVDLA_CSC_wl.scala 439:63:@14694.4]
  wire [318:0] _T_1186; // @[NV_NVDLA_CSC_wl.scala 439:63:@14694.4]
  wire [318:0] _GEN_38; // @[NV_NVDLA_CSC_wl.scala 441:28:@14695.4]
  reg [511:0] _T_1193; // @[NV_NVDLA_CSC_wl.scala 447:40:@14699.4]
  reg [511:0] _RAND_43;
  wire [511:0] _T_1199; // @[NV_NVDLA_CSC_wl.scala 450:49:@14705.4]
  wire [511:0] _T_1208; // @[NV_NVDLA_CSC_wl.scala 453:84:@14710.4]
  wire [511:0] _T_1209; // @[NV_NVDLA_CSC_wl.scala 453:33:@14711.4]
  wire [4:0] _T_1215; // @[NV_NVDLA_CSC_wl.scala 456:52:@14717.4]
  wire [5:0] _T_1217; // @[Cat.scala 30:58:@14718.4]
  wire [5:0] _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@14720.4]
  wire [6:0] _T_1219; // @[NV_NVDLA_CSC_wl.scala 456:69:@14720.4]
  wire [5:0] _T_1220; // @[NV_NVDLA_CSC_wl.scala 456:69:@14721.4]
  wire [511:0] _GEN_39; // @[NV_NVDLA_CSC_wl.scala 458:34:@14722.4]
  wire [511:0] _GEN_40; // @[NV_NVDLA_CSC_wl.scala 461:39:@14725.4]
  reg  _T_1223; // @[NV_NVDLA_CSC_wl.scala 466:36:@14728.4]
  reg [31:0] _RAND_44;
  reg [6:0] _T_1226; // @[NV_NVDLA_CSC_wl.scala 467:37:@14729.4]
  reg [31:0] _RAND_45;
  reg  _T_1229; // @[NV_NVDLA_CSC_wl.scala 468:36:@14730.4]
  reg [31:0] _RAND_46;
  reg  _T_1232; // @[NV_NVDLA_CSC_wl.scala 469:37:@14731.4]
  reg [31:0] _RAND_47;
  reg  _T_1235; // @[NV_NVDLA_CSC_wl.scala 470:35:@14732.4]
  reg [31:0] _RAND_48;
  reg  _T_1238; // @[NV_NVDLA_CSC_wl.scala 471:29:@14733.4]
  reg [31:0] _RAND_49;
  reg [8:0] _T_1241; // @[NV_NVDLA_CSC_wl.scala 472:41:@14734.4]
  reg [31:0] _RAND_50;
  reg [1:0] _T_1244; // @[NV_NVDLA_CSC_wl.scala 473:35:@14735.4]
  reg [31:0] _RAND_51;
  reg [6:0] _T_1247; // @[NV_NVDLA_CSC_wl.scala 474:35:@14736.4]
  reg [31:0] _RAND_52;
  wire [6:0] _GEN_41; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire  _GEN_42; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire  _GEN_43; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire  _GEN_44; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire  _GEN_45; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire [8:0] _GEN_46; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire [1:0] _GEN_47; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire [6:0] _GEN_48; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_wl.scala 497:40:@14749.4]
  wire  _T_1319; // @[NV_NVDLA_CSC_wl.scala 497:40:@14751.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_wl.scala 497:40:@14753.4]
  wire  _T_1321; // @[NV_NVDLA_CSC_wl.scala 497:40:@14755.4]
  wire  _T_1322; // @[NV_NVDLA_CSC_wl.scala 497:40:@14757.4]
  wire  _T_1323; // @[NV_NVDLA_CSC_wl.scala 497:40:@14759.4]
  wire  _T_1324; // @[NV_NVDLA_CSC_wl.scala 497:40:@14761.4]
  wire  _T_1325; // @[NV_NVDLA_CSC_wl.scala 497:40:@14763.4]
  wire  _T_1326; // @[NV_NVDLA_CSC_wl.scala 497:40:@14765.4]
  wire  _T_1327; // @[NV_NVDLA_CSC_wl.scala 497:40:@14767.4]
  wire  _T_1328; // @[NV_NVDLA_CSC_wl.scala 497:40:@14769.4]
  wire  _T_1329; // @[NV_NVDLA_CSC_wl.scala 497:40:@14771.4]
  wire  _T_1330; // @[NV_NVDLA_CSC_wl.scala 497:40:@14773.4]
  wire  _T_1331; // @[NV_NVDLA_CSC_wl.scala 497:40:@14775.4]
  wire  _T_1332; // @[NV_NVDLA_CSC_wl.scala 497:40:@14777.4]
  wire  _T_1333; // @[NV_NVDLA_CSC_wl.scala 497:40:@14779.4]
  wire  _T_1334; // @[NV_NVDLA_CSC_wl.scala 497:40:@14781.4]
  wire  _T_1335; // @[NV_NVDLA_CSC_wl.scala 497:40:@14783.4]
  wire  _T_1336; // @[NV_NVDLA_CSC_wl.scala 497:40:@14785.4]
  wire  _T_1337; // @[NV_NVDLA_CSC_wl.scala 497:40:@14787.4]
  wire  _T_1338; // @[NV_NVDLA_CSC_wl.scala 497:40:@14789.4]
  wire  _T_1339; // @[NV_NVDLA_CSC_wl.scala 497:40:@14791.4]
  wire  _T_1340; // @[NV_NVDLA_CSC_wl.scala 497:40:@14793.4]
  wire  _T_1341; // @[NV_NVDLA_CSC_wl.scala 497:40:@14795.4]
  wire  _T_1342; // @[NV_NVDLA_CSC_wl.scala 497:40:@14797.4]
  wire  _T_1343; // @[NV_NVDLA_CSC_wl.scala 497:40:@14799.4]
  wire  _T_1344; // @[NV_NVDLA_CSC_wl.scala 497:40:@14801.4]
  wire  _T_1345; // @[NV_NVDLA_CSC_wl.scala 497:40:@14803.4]
  wire  _T_1346; // @[NV_NVDLA_CSC_wl.scala 497:40:@14805.4]
  wire  _T_1347; // @[NV_NVDLA_CSC_wl.scala 497:40:@14807.4]
  wire  _T_1348; // @[NV_NVDLA_CSC_wl.scala 497:40:@14809.4]
  wire  _T_1349; // @[NV_NVDLA_CSC_wl.scala 497:40:@14811.4]
  wire  _T_1350; // @[NV_NVDLA_CSC_wl.scala 497:40:@14813.4]
  wire  _T_1351; // @[NV_NVDLA_CSC_wl.scala 497:40:@14815.4]
  wire  _T_1352; // @[NV_NVDLA_CSC_wl.scala 497:40:@14817.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_wl.scala 497:40:@14819.4]
  wire  _T_1354; // @[NV_NVDLA_CSC_wl.scala 497:40:@14821.4]
  wire  _T_1355; // @[NV_NVDLA_CSC_wl.scala 497:40:@14823.4]
  wire  _T_1356; // @[NV_NVDLA_CSC_wl.scala 497:40:@14825.4]
  wire  _T_1357; // @[NV_NVDLA_CSC_wl.scala 497:40:@14827.4]
  wire  _T_1358; // @[NV_NVDLA_CSC_wl.scala 497:40:@14829.4]
  wire  _T_1359; // @[NV_NVDLA_CSC_wl.scala 497:40:@14831.4]
  wire  _T_1360; // @[NV_NVDLA_CSC_wl.scala 497:40:@14833.4]
  wire  _T_1361; // @[NV_NVDLA_CSC_wl.scala 497:40:@14835.4]
  wire  _T_1362; // @[NV_NVDLA_CSC_wl.scala 497:40:@14837.4]
  wire  _T_1363; // @[NV_NVDLA_CSC_wl.scala 497:40:@14839.4]
  wire  _T_1364; // @[NV_NVDLA_CSC_wl.scala 497:40:@14841.4]
  wire  _T_1365; // @[NV_NVDLA_CSC_wl.scala 497:40:@14843.4]
  wire  _T_1366; // @[NV_NVDLA_CSC_wl.scala 497:40:@14845.4]
  wire  _T_1367; // @[NV_NVDLA_CSC_wl.scala 497:40:@14847.4]
  wire  _T_1368; // @[NV_NVDLA_CSC_wl.scala 497:40:@14849.4]
  wire  _T_1369; // @[NV_NVDLA_CSC_wl.scala 497:40:@14851.4]
  wire  _T_1370; // @[NV_NVDLA_CSC_wl.scala 497:40:@14853.4]
  wire  _T_1371; // @[NV_NVDLA_CSC_wl.scala 497:40:@14855.4]
  wire  _T_1372; // @[NV_NVDLA_CSC_wl.scala 497:40:@14857.4]
  wire  _T_1373; // @[NV_NVDLA_CSC_wl.scala 497:40:@14859.4]
  wire  _T_1374; // @[NV_NVDLA_CSC_wl.scala 497:40:@14861.4]
  wire  _T_1375; // @[NV_NVDLA_CSC_wl.scala 497:40:@14863.4]
  wire  _T_1376; // @[NV_NVDLA_CSC_wl.scala 497:40:@14865.4]
  wire  _T_1377; // @[NV_NVDLA_CSC_wl.scala 497:40:@14867.4]
  wire  _T_1378; // @[NV_NVDLA_CSC_wl.scala 497:40:@14869.4]
  wire  _T_1379; // @[NV_NVDLA_CSC_wl.scala 497:40:@14871.4]
  wire  _T_1380; // @[NV_NVDLA_CSC_wl.scala 497:40:@14873.4]
  wire  _T_1381; // @[NV_NVDLA_CSC_wl.scala 497:40:@14875.4]
  wire [1:0] _T_1382; // @[NV_NVDLA_CSC_wl.scala 499:46:@14877.4]
  wire [1:0] _GEN_507; // @[NV_NVDLA_CSC_wl.scala 499:46:@14878.4]
  wire [2:0] _T_1383; // @[NV_NVDLA_CSC_wl.scala 499:46:@14878.4]
  wire [2:0] _GEN_508; // @[NV_NVDLA_CSC_wl.scala 499:46:@14879.4]
  wire [3:0] _T_1384; // @[NV_NVDLA_CSC_wl.scala 499:46:@14879.4]
  wire [3:0] _GEN_509; // @[NV_NVDLA_CSC_wl.scala 499:46:@14880.4]
  wire [4:0] _T_1385; // @[NV_NVDLA_CSC_wl.scala 499:46:@14880.4]
  wire [4:0] _GEN_510; // @[NV_NVDLA_CSC_wl.scala 499:46:@14881.4]
  wire [5:0] _T_1386; // @[NV_NVDLA_CSC_wl.scala 499:46:@14881.4]
  wire [5:0] _GEN_511; // @[NV_NVDLA_CSC_wl.scala 499:46:@14882.4]
  wire [6:0] _T_1387; // @[NV_NVDLA_CSC_wl.scala 499:46:@14882.4]
  wire [6:0] _GEN_512; // @[NV_NVDLA_CSC_wl.scala 499:46:@14883.4]
  wire [7:0] _T_1388; // @[NV_NVDLA_CSC_wl.scala 499:46:@14883.4]
  wire [7:0] _GEN_513; // @[NV_NVDLA_CSC_wl.scala 499:46:@14884.4]
  wire [8:0] _T_1389; // @[NV_NVDLA_CSC_wl.scala 499:46:@14884.4]
  wire [8:0] _GEN_514; // @[NV_NVDLA_CSC_wl.scala 499:46:@14885.4]
  wire [9:0] _T_1390; // @[NV_NVDLA_CSC_wl.scala 499:46:@14885.4]
  wire [9:0] _GEN_515; // @[NV_NVDLA_CSC_wl.scala 499:46:@14886.4]
  wire [10:0] _T_1391; // @[NV_NVDLA_CSC_wl.scala 499:46:@14886.4]
  wire [10:0] _GEN_516; // @[NV_NVDLA_CSC_wl.scala 499:46:@14887.4]
  wire [11:0] _T_1392; // @[NV_NVDLA_CSC_wl.scala 499:46:@14887.4]
  wire [11:0] _GEN_517; // @[NV_NVDLA_CSC_wl.scala 499:46:@14888.4]
  wire [12:0] _T_1393; // @[NV_NVDLA_CSC_wl.scala 499:46:@14888.4]
  wire [12:0] _GEN_518; // @[NV_NVDLA_CSC_wl.scala 499:46:@14889.4]
  wire [13:0] _T_1394; // @[NV_NVDLA_CSC_wl.scala 499:46:@14889.4]
  wire [13:0] _GEN_519; // @[NV_NVDLA_CSC_wl.scala 499:46:@14890.4]
  wire [14:0] _T_1395; // @[NV_NVDLA_CSC_wl.scala 499:46:@14890.4]
  wire [14:0] _GEN_520; // @[NV_NVDLA_CSC_wl.scala 499:46:@14891.4]
  wire [15:0] _T_1396; // @[NV_NVDLA_CSC_wl.scala 499:46:@14891.4]
  wire [15:0] _GEN_521; // @[NV_NVDLA_CSC_wl.scala 499:46:@14892.4]
  wire [16:0] _T_1397; // @[NV_NVDLA_CSC_wl.scala 499:46:@14892.4]
  wire [16:0] _GEN_522; // @[NV_NVDLA_CSC_wl.scala 499:46:@14893.4]
  wire [17:0] _T_1398; // @[NV_NVDLA_CSC_wl.scala 499:46:@14893.4]
  wire [17:0] _GEN_523; // @[NV_NVDLA_CSC_wl.scala 499:46:@14894.4]
  wire [18:0] _T_1399; // @[NV_NVDLA_CSC_wl.scala 499:46:@14894.4]
  wire [18:0] _GEN_524; // @[NV_NVDLA_CSC_wl.scala 499:46:@14895.4]
  wire [19:0] _T_1400; // @[NV_NVDLA_CSC_wl.scala 499:46:@14895.4]
  wire [19:0] _GEN_525; // @[NV_NVDLA_CSC_wl.scala 499:46:@14896.4]
  wire [20:0] _T_1401; // @[NV_NVDLA_CSC_wl.scala 499:46:@14896.4]
  wire [20:0] _GEN_526; // @[NV_NVDLA_CSC_wl.scala 499:46:@14897.4]
  wire [21:0] _T_1402; // @[NV_NVDLA_CSC_wl.scala 499:46:@14897.4]
  wire [21:0] _GEN_527; // @[NV_NVDLA_CSC_wl.scala 499:46:@14898.4]
  wire [22:0] _T_1403; // @[NV_NVDLA_CSC_wl.scala 499:46:@14898.4]
  wire [22:0] _GEN_528; // @[NV_NVDLA_CSC_wl.scala 499:46:@14899.4]
  wire [23:0] _T_1404; // @[NV_NVDLA_CSC_wl.scala 499:46:@14899.4]
  wire [23:0] _GEN_529; // @[NV_NVDLA_CSC_wl.scala 499:46:@14900.4]
  wire [24:0] _T_1405; // @[NV_NVDLA_CSC_wl.scala 499:46:@14900.4]
  wire [24:0] _GEN_530; // @[NV_NVDLA_CSC_wl.scala 499:46:@14901.4]
  wire [25:0] _T_1406; // @[NV_NVDLA_CSC_wl.scala 499:46:@14901.4]
  wire [25:0] _GEN_531; // @[NV_NVDLA_CSC_wl.scala 499:46:@14902.4]
  wire [26:0] _T_1407; // @[NV_NVDLA_CSC_wl.scala 499:46:@14902.4]
  wire [26:0] _GEN_532; // @[NV_NVDLA_CSC_wl.scala 499:46:@14903.4]
  wire [27:0] _T_1408; // @[NV_NVDLA_CSC_wl.scala 499:46:@14903.4]
  wire [27:0] _GEN_533; // @[NV_NVDLA_CSC_wl.scala 499:46:@14904.4]
  wire [28:0] _T_1409; // @[NV_NVDLA_CSC_wl.scala 499:46:@14904.4]
  wire [28:0] _GEN_534; // @[NV_NVDLA_CSC_wl.scala 499:46:@14905.4]
  wire [29:0] _T_1410; // @[NV_NVDLA_CSC_wl.scala 499:46:@14905.4]
  wire [29:0] _GEN_535; // @[NV_NVDLA_CSC_wl.scala 499:46:@14906.4]
  wire [30:0] _T_1411; // @[NV_NVDLA_CSC_wl.scala 499:46:@14906.4]
  wire [30:0] _GEN_536; // @[NV_NVDLA_CSC_wl.scala 499:46:@14907.4]
  wire [31:0] _T_1412; // @[NV_NVDLA_CSC_wl.scala 499:46:@14907.4]
  wire [31:0] _GEN_537; // @[NV_NVDLA_CSC_wl.scala 499:46:@14908.4]
  wire [32:0] _T_1413; // @[NV_NVDLA_CSC_wl.scala 499:46:@14908.4]
  wire [32:0] _GEN_538; // @[NV_NVDLA_CSC_wl.scala 499:46:@14909.4]
  wire [33:0] _T_1414; // @[NV_NVDLA_CSC_wl.scala 499:46:@14909.4]
  wire [33:0] _GEN_539; // @[NV_NVDLA_CSC_wl.scala 499:46:@14910.4]
  wire [34:0] _T_1415; // @[NV_NVDLA_CSC_wl.scala 499:46:@14910.4]
  wire [34:0] _GEN_540; // @[NV_NVDLA_CSC_wl.scala 499:46:@14911.4]
  wire [35:0] _T_1416; // @[NV_NVDLA_CSC_wl.scala 499:46:@14911.4]
  wire [35:0] _GEN_541; // @[NV_NVDLA_CSC_wl.scala 499:46:@14912.4]
  wire [36:0] _T_1417; // @[NV_NVDLA_CSC_wl.scala 499:46:@14912.4]
  wire [36:0] _GEN_542; // @[NV_NVDLA_CSC_wl.scala 499:46:@14913.4]
  wire [37:0] _T_1418; // @[NV_NVDLA_CSC_wl.scala 499:46:@14913.4]
  wire [37:0] _GEN_543; // @[NV_NVDLA_CSC_wl.scala 499:46:@14914.4]
  wire [38:0] _T_1419; // @[NV_NVDLA_CSC_wl.scala 499:46:@14914.4]
  wire [38:0] _GEN_544; // @[NV_NVDLA_CSC_wl.scala 499:46:@14915.4]
  wire [39:0] _T_1420; // @[NV_NVDLA_CSC_wl.scala 499:46:@14915.4]
  wire [39:0] _GEN_545; // @[NV_NVDLA_CSC_wl.scala 499:46:@14916.4]
  wire [40:0] _T_1421; // @[NV_NVDLA_CSC_wl.scala 499:46:@14916.4]
  wire [40:0] _GEN_546; // @[NV_NVDLA_CSC_wl.scala 499:46:@14917.4]
  wire [41:0] _T_1422; // @[NV_NVDLA_CSC_wl.scala 499:46:@14917.4]
  wire [41:0] _GEN_547; // @[NV_NVDLA_CSC_wl.scala 499:46:@14918.4]
  wire [42:0] _T_1423; // @[NV_NVDLA_CSC_wl.scala 499:46:@14918.4]
  wire [42:0] _GEN_548; // @[NV_NVDLA_CSC_wl.scala 499:46:@14919.4]
  wire [43:0] _T_1424; // @[NV_NVDLA_CSC_wl.scala 499:46:@14919.4]
  wire [43:0] _GEN_549; // @[NV_NVDLA_CSC_wl.scala 499:46:@14920.4]
  wire [44:0] _T_1425; // @[NV_NVDLA_CSC_wl.scala 499:46:@14920.4]
  wire [44:0] _GEN_550; // @[NV_NVDLA_CSC_wl.scala 499:46:@14921.4]
  wire [45:0] _T_1426; // @[NV_NVDLA_CSC_wl.scala 499:46:@14921.4]
  wire [45:0] _GEN_551; // @[NV_NVDLA_CSC_wl.scala 499:46:@14922.4]
  wire [46:0] _T_1427; // @[NV_NVDLA_CSC_wl.scala 499:46:@14922.4]
  wire [46:0] _GEN_552; // @[NV_NVDLA_CSC_wl.scala 499:46:@14923.4]
  wire [47:0] _T_1428; // @[NV_NVDLA_CSC_wl.scala 499:46:@14923.4]
  wire [47:0] _GEN_553; // @[NV_NVDLA_CSC_wl.scala 499:46:@14924.4]
  wire [48:0] _T_1429; // @[NV_NVDLA_CSC_wl.scala 499:46:@14924.4]
  wire [48:0] _GEN_554; // @[NV_NVDLA_CSC_wl.scala 499:46:@14925.4]
  wire [49:0] _T_1430; // @[NV_NVDLA_CSC_wl.scala 499:46:@14925.4]
  wire [49:0] _GEN_555; // @[NV_NVDLA_CSC_wl.scala 499:46:@14926.4]
  wire [50:0] _T_1431; // @[NV_NVDLA_CSC_wl.scala 499:46:@14926.4]
  wire [50:0] _GEN_556; // @[NV_NVDLA_CSC_wl.scala 499:46:@14927.4]
  wire [51:0] _T_1432; // @[NV_NVDLA_CSC_wl.scala 499:46:@14927.4]
  wire [51:0] _GEN_557; // @[NV_NVDLA_CSC_wl.scala 499:46:@14928.4]
  wire [52:0] _T_1433; // @[NV_NVDLA_CSC_wl.scala 499:46:@14928.4]
  wire [52:0] _GEN_558; // @[NV_NVDLA_CSC_wl.scala 499:46:@14929.4]
  wire [53:0] _T_1434; // @[NV_NVDLA_CSC_wl.scala 499:46:@14929.4]
  wire [53:0] _GEN_559; // @[NV_NVDLA_CSC_wl.scala 499:46:@14930.4]
  wire [54:0] _T_1435; // @[NV_NVDLA_CSC_wl.scala 499:46:@14930.4]
  wire [54:0] _GEN_560; // @[NV_NVDLA_CSC_wl.scala 499:46:@14931.4]
  wire [55:0] _T_1436; // @[NV_NVDLA_CSC_wl.scala 499:46:@14931.4]
  wire [55:0] _GEN_561; // @[NV_NVDLA_CSC_wl.scala 499:46:@14932.4]
  wire [56:0] _T_1437; // @[NV_NVDLA_CSC_wl.scala 499:46:@14932.4]
  wire [56:0] _GEN_562; // @[NV_NVDLA_CSC_wl.scala 499:46:@14933.4]
  wire [57:0] _T_1438; // @[NV_NVDLA_CSC_wl.scala 499:46:@14933.4]
  wire [57:0] _GEN_563; // @[NV_NVDLA_CSC_wl.scala 499:46:@14934.4]
  wire [58:0] _T_1439; // @[NV_NVDLA_CSC_wl.scala 499:46:@14934.4]
  wire [58:0] _GEN_564; // @[NV_NVDLA_CSC_wl.scala 499:46:@14935.4]
  wire [59:0] _T_1440; // @[NV_NVDLA_CSC_wl.scala 499:46:@14935.4]
  wire [59:0] _GEN_565; // @[NV_NVDLA_CSC_wl.scala 499:46:@14936.4]
  wire [60:0] _T_1441; // @[NV_NVDLA_CSC_wl.scala 499:46:@14936.4]
  wire [60:0] _GEN_566; // @[NV_NVDLA_CSC_wl.scala 499:46:@14937.4]
  wire [61:0] _T_1442; // @[NV_NVDLA_CSC_wl.scala 499:46:@14937.4]
  wire [61:0] _GEN_567; // @[NV_NVDLA_CSC_wl.scala 499:46:@14938.4]
  wire [62:0] _T_1443; // @[NV_NVDLA_CSC_wl.scala 499:46:@14938.4]
  wire [62:0] _GEN_568; // @[NV_NVDLA_CSC_wl.scala 499:46:@14939.4]
  wire [63:0] _T_1444; // @[NV_NVDLA_CSC_wl.scala 499:46:@14939.4]
  reg [63:0] _T_1447; // @[NV_NVDLA_CSC_wl.scala 502:33:@14940.4]
  reg [63:0] _RAND_53;
  wire [190:0] _T_1453; // @[NV_NVDLA_CSC_wl.scala 505:57:@14942.4]
  wire [190:0] _T_1454; // @[NV_NVDLA_CSC_wl.scala 505:26:@14943.4]
  wire  _T_1456; // @[NV_NVDLA_CSC_wl.scala 508:45:@14944.4]
  wire [63:0] _T_1467; // @[NV_NVDLA_CSC_wl.scala 508:27:@14947.4]
  wire  _T_1469; // @[NV_NVDLA_CSC_wl.scala 509:45:@14948.4]
  wire [63:0] _T_1480; // @[NV_NVDLA_CSC_wl.scala 509:27:@14951.4]
  wire  _T_1482; // @[NV_NVDLA_CSC_wl.scala 510:45:@14952.4]
  wire [63:0] _T_1493; // @[NV_NVDLA_CSC_wl.scala 510:27:@14955.4]
  wire [5:0] _T_1494; // @[NV_NVDLA_CSC_wl.scala 514:50:@14956.4]
  wire [6:0] _T_1496; // @[Cat.scala 30:58:@14957.4]
  wire [63:0] _T_1497; // @[NV_NVDLA_CSC_wl.scala 515:39:@14958.4]
  wire [190:0] _GEN_569; // @[NV_NVDLA_CSC_wl.scala 515:61:@14959.4]
  wire [190:0] _T_1498; // @[NV_NVDLA_CSC_wl.scala 515:61:@14959.4]
  wire [63:0] _T_1500; // @[NV_NVDLA_CSC_wl.scala 516:62:@14961.4]
  wire [190:0] _GEN_570; // @[NV_NVDLA_CSC_wl.scala 516:83:@14962.4]
  wire [190:0] _T_1501; // @[NV_NVDLA_CSC_wl.scala 516:83:@14962.4]
  wire [190:0] _GEN_571; // @[NV_NVDLA_CSC_wl.scala 516:100:@14963.4]
  wire [190:0] _T_1502; // @[NV_NVDLA_CSC_wl.scala 516:100:@14963.4]
  wire [63:0] _T_1504; // @[NV_NVDLA_CSC_wl.scala 517:62:@14965.4]
  wire [190:0] _GEN_572; // @[NV_NVDLA_CSC_wl.scala 517:83:@14966.4]
  wire [190:0] _T_1505; // @[NV_NVDLA_CSC_wl.scala 517:83:@14966.4]
  wire [190:0] _GEN_573; // @[NV_NVDLA_CSC_wl.scala 517:100:@14967.4]
  wire [190:0] _T_1506; // @[NV_NVDLA_CSC_wl.scala 517:100:@14967.4]
  wire [63:0] _T_1508; // @[NV_NVDLA_CSC_wl.scala 518:62:@14969.4]
  wire [190:0] _GEN_574; // @[NV_NVDLA_CSC_wl.scala 518:83:@14970.4]
  wire [190:0] _T_1509; // @[NV_NVDLA_CSC_wl.scala 518:83:@14970.4]
  wire [190:0] _GEN_575; // @[NV_NVDLA_CSC_wl.scala 518:100:@14971.4]
  wire [190:0] _T_1510; // @[NV_NVDLA_CSC_wl.scala 518:100:@14971.4]
  wire  _T_1517; // @[NV_NVDLA_CSC_wl.scala 523:41:@14973.4]
  wire  _T_1519; // @[NV_NVDLA_CSC_wl.scala 524:41:@14974.4]
  wire [31:0] _T_1520; // @[NV_NVDLA_CSC_wl.scala 524:82:@14975.4]
  wire [31:0] _T_1521; // @[NV_NVDLA_CSC_wl.scala 524:122:@14976.4]
  wire [63:0] _T_1522; // @[Cat.scala 30:58:@14977.4]
  wire [15:0] _T_1523; // @[NV_NVDLA_CSC_wl.scala 525:44:@14978.4]
  wire [15:0] _T_1524; // @[NV_NVDLA_CSC_wl.scala 525:84:@14979.4]
  wire [15:0] _T_1525; // @[NV_NVDLA_CSC_wl.scala 525:124:@14980.4]
  wire [15:0] _T_1526; // @[NV_NVDLA_CSC_wl.scala 525:164:@14981.4]
  wire [63:0] _T_1529; // @[Cat.scala 30:58:@14984.4]
  wire [63:0] _T_1530; // @[NV_NVDLA_CSC_wl.scala 524:28:@14985.4]
  wire [190:0] _T_1531; // @[NV_NVDLA_CSC_wl.scala 523:28:@14986.4]
  wire [190:0] _T_1532; // @[NV_NVDLA_CSC_wl.scala 522:28:@14987.4]
  wire [190:0] _GEN_576; // @[NV_NVDLA_CSC_wl.scala 528:61:@14988.4]
  wire  _T_1533; // @[NV_NVDLA_CSC_wl.scala 528:61:@14988.4]
  wire  _T_1534; // @[NV_NVDLA_CSC_wl.scala 528:44:@14989.4]
  reg [7:0] _T_1537; // @[NV_NVDLA_CSC_wl.scala 531:30:@14990.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_1540; // @[NV_NVDLA_CSC_wl.scala 532:35:@14991.4]
  reg [31:0] _RAND_55;
  wire [63:0] _GEN_577; // @[NV_NVDLA_CSC_wl.scala 534:57:@14992.4]
  wire  _T_1541; // @[NV_NVDLA_CSC_wl.scala 534:57:@14992.4]
  wire  _T_1542; // @[NV_NVDLA_CSC_wl.scala 534:42:@14993.4]
  wire  _T_1543; // @[NV_NVDLA_CSC_wl.scala 536:31:@14994.4]
  wire [7:0] _T_1546; // @[NV_NVDLA_CSC_wl.scala 536:30:@14995.4]
  wire [8:0] _T_1547; // @[NV_NVDLA_CSC_wl.scala 538:39:@14996.4]
  wire [7:0] _T_1548; // @[NV_NVDLA_CSC_wl.scala 538:39:@14997.4]
  wire [63:0] _GEN_578; // @[NV_NVDLA_CSC_wl.scala 538:57:@14998.4]
  wire [64:0] _T_1549; // @[NV_NVDLA_CSC_wl.scala 538:57:@14998.4]
  wire [64:0] _T_1550; // @[NV_NVDLA_CSC_wl.scala 538:57:@14999.4]
  wire [63:0] _T_1551; // @[NV_NVDLA_CSC_wl.scala 538:57:@15000.4]
  wire  _T_1553; // @[NV_NVDLA_CSC_wl.scala 540:29:@15001.4]
  wire  _T_1554; // @[NV_NVDLA_CSC_wl.scala 540:47:@15002.4]
  wire [63:0] _T_1555; // @[NV_NVDLA_CSC_wl.scala 540:28:@15003.4]
  wire [63:0] _T_1556; // @[NV_NVDLA_CSC_wl.scala 539:28:@15004.4]
  wire  _T_1557; // @[NV_NVDLA_CSC_wl.scala 543:61:@15005.4]
  wire  _T_1558; // @[NV_NVDLA_CSC_wl.scala 543:81:@15006.4]
  wire  _T_1559; // @[NV_NVDLA_CSC_wl.scala 543:40:@15007.4]
  wire  _T_1560; // @[NV_NVDLA_CSC_wl.scala 545:19:@15008.4]
  wire [63:0] _GEN_49; // @[NV_NVDLA_CSC_wl.scala 545:39:@15009.4]
  wire [63:0] _GEN_50; // @[NV_NVDLA_CSC_wl.scala 548:30:@15012.4]
  reg [12:0] _T_1563; // @[NV_NVDLA_CSC_wl.scala 553:30:@15015.4]
  reg [31:0] _RAND_56;
  reg [12:0] _T_1566; // @[NV_NVDLA_CSC_wl.scala 554:35:@15016.4]
  reg [31:0] _RAND_57;
  wire [13:0] _T_1568; // @[NV_NVDLA_CSC_wl.scala 556:39:@15017.4]
  wire [12:0] _T_1569; // @[NV_NVDLA_CSC_wl.scala 556:39:@15018.4]
  wire [13:0] _GEN_579; // @[NV_NVDLA_CSC_wl.scala 557:48:@15021.4]
  wire  _T_1576; // @[NV_NVDLA_CSC_wl.scala 557:48:@15021.4]
  wire [12:0] _T_1582; // @[NV_NVDLA_CSC_wl.scala 558:35:@15023.4]
  wire [12:0] _T_1583; // @[NV_NVDLA_CSC_wl.scala 560:53:@15024.4]
  wire [12:0] _T_1586; // @[NV_NVDLA_CSC_wl.scala 562:28:@15027.4]
  wire [12:0] _T_1587; // @[NV_NVDLA_CSC_wl.scala 561:28:@15028.4]
  wire [12:0] _T_1588; // @[NV_NVDLA_CSC_wl.scala 560:28:@15029.4]
  wire  _T_1589; // @[NV_NVDLA_CSC_wl.scala 566:40:@15030.4]
  wire  _T_1590; // @[NV_NVDLA_CSC_wl.scala 566:76:@15031.4]
  wire  _T_1591; // @[NV_NVDLA_CSC_wl.scala 566:55:@15032.4]
  wire  _T_1592; // @[NV_NVDLA_CSC_wl.scala 567:66:@15033.4]
  wire  _T_1593; // @[NV_NVDLA_CSC_wl.scala 567:86:@15034.4]
  wire  _T_1594; // @[NV_NVDLA_CSC_wl.scala 567:45:@15035.4]
  wire [13:0] _T_1600; // @[Cat.scala 30:58:@15037.4]
  wire [13:0] _GEN_580; // @[NV_NVDLA_CSC_wl.scala 568:39:@15038.4]
  wire [14:0] _T_1601; // @[NV_NVDLA_CSC_wl.scala 568:39:@15038.4]
  wire [13:0] _T_1602; // @[NV_NVDLA_CSC_wl.scala 568:39:@15039.4]
  wire [12:0] _GEN_51; // @[NV_NVDLA_CSC_wl.scala 570:29:@15040.4]
  wire [12:0] _GEN_52; // @[NV_NVDLA_CSC_wl.scala 573:34:@15043.4]
  reg  _T_1605; // @[NV_NVDLA_CSC_wl.scala 578:33:@15046.4]
  reg [31:0] _RAND_58;
  reg [14:0] _T_1608; // @[NV_NVDLA_CSC_wl.scala 579:29:@15047.4]
  reg [31:0] _RAND_59;
  wire  _T_1609; // @[NV_NVDLA_CSC_wl.scala 581:42:@15048.4]
  wire  _T_1612; // @[NV_NVDLA_CSC_wl.scala 581:76:@15049.4]
  wire  _T_1613; // @[NV_NVDLA_CSC_wl.scala 581:31:@15050.4]
  wire [15:0] _T_1615; // @[NV_NVDLA_CSC_wl.scala 582:37:@15051.4]
  wire [14:0] _T_1616; // @[NV_NVDLA_CSC_wl.scala 582:37:@15052.4]
  wire [14:0] _T_1619; // @[NV_NVDLA_CSC_wl.scala 583:84:@15053.4]
  wire [14:0] _T_1620; // @[NV_NVDLA_CSC_wl.scala 583:27:@15054.4]
  wire  _T_1621; // @[NV_NVDLA_CSC_wl.scala 584:59:@15055.4]
  wire  _T_1622; // @[NV_NVDLA_CSC_wl.scala 584:38:@15056.4]
  wire  _T_1623; // @[NV_NVDLA_CSC_wl.scala 584:82:@15057.4]
  wire  _T_1624; // @[NV_NVDLA_CSC_wl.scala 584:98:@15058.4]
  wire  _T_1625; // @[NV_NVDLA_CSC_wl.scala 584:79:@15059.4]
  wire  _T_1627; // @[NV_NVDLA_CSC_wl.scala 585:45:@15061.4]
  wire [14:0] _T_1628; // @[NV_NVDLA_CSC_wl.scala 585:29:@15062.4]
  wire [14:0] _GEN_53; // @[NV_NVDLA_CSC_wl.scala 588:28:@15064.4]
  reg  _T_1631; // @[NV_NVDLA_CSC_wl.scala 593:38:@15067.4]
  reg [31:0] _RAND_60;
  reg [12:0] _T_1634; // @[NV_NVDLA_CSC_wl.scala 594:40:@15068.4]
  reg [31:0] _RAND_61;
  reg  _T_1637; // @[NV_NVDLA_CSC_wl.scala 596:39:@15069.4]
  reg [31:0] _RAND_62;
  reg  _T_1640; // @[NV_NVDLA_CSC_wl.scala 597:39:@15070.4]
  reg [31:0] _RAND_63;
  reg  _T_1643; // @[NV_NVDLA_CSC_wl.scala 598:40:@15071.4]
  reg [31:0] _RAND_64;
  reg  _T_1646; // @[NV_NVDLA_CSC_wl.scala 599:38:@15072.4]
  reg [31:0] _RAND_65;
  reg  _T_1649; // @[NV_NVDLA_CSC_wl.scala 600:32:@15073.4]
  reg [31:0] _RAND_66;
  reg [7:0] _T_1652; // @[NV_NVDLA_CSC_wl.scala 601:34:@15074.4]
  reg [31:0] _RAND_67;
  reg  _T_1655; // @[NV_NVDLA_CSC_wl.scala 603:36:@15075.4]
  reg [31:0] _RAND_68;
  reg [8:0] _T_1658; // @[NV_NVDLA_CSC_wl.scala 604:44:@15076.4]
  reg [31:0] _RAND_69;
  reg [14:0] _T_1661; // @[NV_NVDLA_CSC_wl.scala 605:43:@15077.4]
  reg [31:0] _RAND_70;
  wire [13:0] _GEN_54; // @[NV_NVDLA_CSC_wl.scala 609:23:@15079.4]
  wire  _GEN_55; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  wire  _GEN_56; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  wire  _GEN_57; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  wire  _GEN_58; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  wire [63:0] _GEN_59; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  wire [190:0] _GEN_60; // @[NV_NVDLA_CSC_wl.scala 621:39:@15091.4]
  wire [8:0] _GEN_61; // @[NV_NVDLA_CSC_wl.scala 625:28:@15095.4]
  wire  _T_1663; // @[NV_NVDLA_CSC_wl.scala 628:28:@15098.4]
  wire [14:0] _GEN_62; // @[NV_NVDLA_CSC_wl.scala 628:41:@15099.4]
  wire [35:0] _T_1672; // @[Cat.scala 30:58:@15112.4]
  reg  _T_1677; // @[NV_NVDLA_CSC_wl.scala 654:76:@15114.4]
  reg [31:0] _RAND_71;
  reg  _T_1680; // @[NV_NVDLA_CSC_wl.scala 654:76:@15115.4]
  reg [31:0] _RAND_72;
  reg  _T_1683; // @[NV_NVDLA_CSC_wl.scala 654:76:@15116.4]
  reg [31:0] _RAND_73;
  reg  _T_1686; // @[NV_NVDLA_CSC_wl.scala 654:76:@15117.4]
  reg [31:0] _RAND_74;
  reg  _T_1689; // @[NV_NVDLA_CSC_wl.scala 654:76:@15118.4]
  reg [31:0] _RAND_75;
  reg [35:0] _T_1697; // @[NV_NVDLA_CSC_wl.scala 656:75:@15121.4]
  reg [63:0] _RAND_76;
  reg [35:0] _T_1700; // @[NV_NVDLA_CSC_wl.scala 656:75:@15122.4]
  reg [63:0] _RAND_77;
  reg [35:0] _T_1703; // @[NV_NVDLA_CSC_wl.scala 656:75:@15123.4]
  reg [63:0] _RAND_78;
  reg [35:0] _T_1706; // @[NV_NVDLA_CSC_wl.scala 656:75:@15124.4]
  reg [63:0] _RAND_79;
  reg [35:0] _T_1709; // @[NV_NVDLA_CSC_wl.scala 656:75:@15125.4]
  reg [63:0] _RAND_80;
  reg  _T_1717; // @[NV_NVDLA_CSC_wl.scala 658:74:@15128.4]
  reg [31:0] _RAND_81;
  reg  _T_1720; // @[NV_NVDLA_CSC_wl.scala 658:74:@15129.4]
  reg [31:0] _RAND_82;
  reg  _T_1723; // @[NV_NVDLA_CSC_wl.scala 658:74:@15130.4]
  reg [31:0] _RAND_83;
  reg  _T_1726; // @[NV_NVDLA_CSC_wl.scala 658:74:@15131.4]
  reg [31:0] _RAND_84;
  reg  _T_1729; // @[NV_NVDLA_CSC_wl.scala 658:74:@15132.4]
  reg [31:0] _RAND_85;
  reg  _T_1732; // @[NV_NVDLA_CSC_wl.scala 658:74:@15133.4]
  reg [31:0] _RAND_86;
  reg [63:0] _T_1737; // @[NV_NVDLA_CSC_wl.scala 660:75:@15135.4]
  reg [63:0] _RAND_87;
  reg [63:0] _T_1740; // @[NV_NVDLA_CSC_wl.scala 660:75:@15136.4]
  reg [63:0] _RAND_88;
  reg [63:0] _T_1743; // @[NV_NVDLA_CSC_wl.scala 660:75:@15137.4]
  reg [63:0] _RAND_89;
  reg [63:0] _T_1746; // @[NV_NVDLA_CSC_wl.scala 660:75:@15138.4]
  reg [63:0] _RAND_90;
  reg [63:0] _T_1749; // @[NV_NVDLA_CSC_wl.scala 660:75:@15139.4]
  reg [63:0] _RAND_91;
  reg [63:0] _T_1752; // @[NV_NVDLA_CSC_wl.scala 660:75:@15140.4]
  reg [63:0] _RAND_92;
  wire [35:0] _GEN_63; // @[NV_NVDLA_CSC_wl.scala 669:36:@15146.4]
  wire [63:0] _GEN_64; // @[NV_NVDLA_CSC_wl.scala 673:34:@15150.4]
  wire [35:0] _GEN_65; // @[NV_NVDLA_CSC_wl.scala 669:36:@15154.4]
  wire [63:0] _GEN_66; // @[NV_NVDLA_CSC_wl.scala 673:34:@15158.4]
  wire [35:0] _GEN_67; // @[NV_NVDLA_CSC_wl.scala 669:36:@15162.4]
  wire [63:0] _GEN_68; // @[NV_NVDLA_CSC_wl.scala 673:34:@15166.4]
  wire [35:0] _GEN_69; // @[NV_NVDLA_CSC_wl.scala 669:36:@15170.4]
  wire [63:0] _GEN_70; // @[NV_NVDLA_CSC_wl.scala 673:34:@15174.4]
  wire [35:0] _GEN_71; // @[NV_NVDLA_CSC_wl.scala 669:36:@15178.4]
  wire [63:0] _GEN_72; // @[NV_NVDLA_CSC_wl.scala 673:34:@15182.4]
  wire [35:0] _GEN_73; // @[NV_NVDLA_CSC_wl.scala 669:36:@15186.4]
  wire [63:0] _GEN_74; // @[NV_NVDLA_CSC_wl.scala 673:34:@15190.4]
  wire [7:0] _T_1753; // @[NV_NVDLA_CSC_wl.scala 687:38:@15194.4]
  wire  _T_1756; // @[NV_NVDLA_CSC_wl.scala 690:44:@15199.4]
  wire  _T_1757; // @[NV_NVDLA_CSC_wl.scala 691:45:@15200.4]
  wire  _T_1758; // @[NV_NVDLA_CSC_wl.scala 692:43:@15201.4]
  reg [6:0] _T_1762; // @[NV_NVDLA_CSC_wl.scala 699:37:@15204.4]
  reg [31:0] _RAND_93;
  reg [6:0] _T_1765; // @[NV_NVDLA_CSC_wl.scala 700:42:@15205.4]
  reg [31:0] _RAND_94;
  wire [7:0] _T_1768; // @[NV_NVDLA_CSC_wl.scala 702:37:@15206.4]
  wire  _T_1770; // @[NV_NVDLA_CSC_wl.scala 704:55:@15207.4]
  wire  _T_1771; // @[NV_NVDLA_CSC_wl.scala 704:53:@15208.4]
  wire [8:0] _T_1773; // @[Cat.scala 30:58:@15209.4]
  wire [7:0] _GEN_581; // @[NV_NVDLA_CSC_wl.scala 704:141:@15210.4]
  wire [8:0] _T_1774; // @[NV_NVDLA_CSC_wl.scala 704:141:@15210.4]
  wire [7:0] _T_1775; // @[NV_NVDLA_CSC_wl.scala 704:141:@15211.4]
  wire [8:0] _T_1776; // @[NV_NVDLA_CSC_wl.scala 704:166:@15212.4]
  wire [8:0] _T_1777; // @[NV_NVDLA_CSC_wl.scala 704:166:@15213.4]
  wire [7:0] _T_1778; // @[NV_NVDLA_CSC_wl.scala 704:166:@15214.4]
  wire [8:0] _T_1779; // @[NV_NVDLA_CSC_wl.scala 704:33:@15215.4]
  wire [8:0] _T_1780; // @[NV_NVDLA_CSC_wl.scala 703:35:@15216.4]
  wire [6:0] _T_1781; // @[NV_NVDLA_CSC_wl.scala 704:182:@15217.4]
  wire  _T_1782; // @[NV_NVDLA_CSC_wl.scala 705:42:@15218.4]
  wire  _T_1783; // @[NV_NVDLA_CSC_wl.scala 706:67:@15219.4]
  wire  _T_1784; // @[NV_NVDLA_CSC_wl.scala 706:47:@15220.4]
  wire [6:0] _GEN_75; // @[NV_NVDLA_CSC_wl.scala 708:32:@15221.4]
  wire [6:0] _GEN_76; // @[NV_NVDLA_CSC_wl.scala 711:37:@15224.4]
  reg [511:0] _T_1786; // @[NV_NVDLA_CSC_wl.scala 716:29:@15227.4]
  reg [511:0] _RAND_95;
  reg [511:0] _T_1788; // @[NV_NVDLA_CSC_wl.scala 717:34:@15228.4]
  reg [511:0] _RAND_96;
  wire [8:0] _T_1790; // @[NV_NVDLA_CSC_wl.scala 719:40:@15230.4]
  wire [8:0] _T_1791; // @[NV_NVDLA_CSC_wl.scala 719:40:@15231.4]
  wire [7:0] _T_1792; // @[NV_NVDLA_CSC_wl.scala 719:40:@15232.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@15234.4]
  wire [511:0] _T_1796; // @[NV_NVDLA_CSC_wl.scala 720:82:@15235.4]
  wire  _T_1798; // @[NV_NVDLA_CSC_wl.scala 721:58:@15236.4]
  wire  _T_1799; // @[NV_NVDLA_CSC_wl.scala 721:38:@15237.4]
  wire [511:0] _T_1801; // @[NV_NVDLA_CSC_wl.scala 721:36:@15238.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@15239.4]
  wire [511:0] _T_1804; // @[NV_NVDLA_CSC_wl.scala 722:45:@15240.4]
  wire  _T_1809; // @[NV_NVDLA_CSC_wl.scala 725:98:@15243.4]
  wire  _T_1810; // @[NV_NVDLA_CSC_wl.scala 725:71:@15244.4]
  wire [511:0] _T_1811; // @[NV_NVDLA_CSC_wl.scala 726:31:@15245.4]
  wire [511:0] _T_1812; // @[NV_NVDLA_CSC_wl.scala 725:31:@15246.4]
  wire [511:0] _T_1813; // @[NV_NVDLA_CSC_wl.scala 724:31:@15247.4]
  wire  _T_1815; // @[NV_NVDLA_CSC_wl.scala 729:86:@15248.4]
  wire  _T_1816; // @[NV_NVDLA_CSC_wl.scala 729:62:@15249.4]
  wire  _T_1817; // @[NV_NVDLA_CSC_wl.scala 729:42:@15250.4]
  wire  _T_1821; // @[NV_NVDLA_CSC_wl.scala 730:86:@15253.4]
  wire  _T_1822; // @[NV_NVDLA_CSC_wl.scala 730:47:@15254.4]
  wire [9:0] _T_1825; // @[Cat.scala 30:58:@15256.4]
  wire [1534:0] _GEN_583; // @[NV_NVDLA_CSC_wl.scala 731:55:@15257.4]
  wire [1534:0] _T_1826; // @[NV_NVDLA_CSC_wl.scala 731:55:@15257.4]
  wire [1534:0] _T_1828; // @[NV_NVDLA_CSC_wl.scala 732:32:@15258.4]
  reg [7:0] _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_97;
  reg [7:0] _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_98;
  reg [7:0] _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_99;
  reg [7:0] _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_100;
  reg [7:0] _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_101;
  reg [7:0] _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_102;
  reg [7:0] _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_103;
  reg [7:0] _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_104;
  reg [7:0] _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_105;
  reg [7:0] _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_106;
  reg [7:0] _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_107;
  reg [7:0] _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_108;
  reg [7:0] _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_109;
  reg [7:0] _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_110;
  reg [7:0] _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_111;
  reg [7:0] _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_112;
  reg [7:0] _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_113;
  reg [7:0] _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_115;
  reg [7:0] _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_116;
  reg [7:0] _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_117;
  reg [7:0] _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_118;
  reg [7:0] _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_119;
  reg [7:0] _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_120;
  reg [7:0] _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_121;
  reg [7:0] _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_122;
  reg [7:0] _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_123;
  reg [7:0] _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_124;
  reg [7:0] _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_125;
  reg [7:0] _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_126;
  reg [7:0] _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_127;
  reg [7:0] _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_128;
  reg [7:0] _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_129;
  reg [7:0] _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_130;
  reg [7:0] _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_131;
  reg [7:0] _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_132;
  reg [7:0] _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_133;
  reg [7:0] _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_134;
  reg [7:0] _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_135;
  reg [7:0] _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_136;
  reg [7:0] _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_144;
  reg [7:0] _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_145;
  reg [7:0] _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_146;
  reg [7:0] _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_147;
  reg [7:0] _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_148;
  reg [7:0] _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_149;
  reg [7:0] _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_150;
  reg [7:0] _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_151;
  reg [7:0] _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_152;
  reg [7:0] _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_153;
  reg [7:0] _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_154;
  reg [7:0] _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_155;
  reg [7:0] _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_156;
  reg [7:0] _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_157;
  reg [7:0] _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_158;
  reg [7:0] _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_159;
  reg [7:0] _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 742:33:@15330.4]
  reg [31:0] _RAND_160;
  wire [1534:0] _GEN_584; // @[NV_NVDLA_CSC_wl.scala 744:42:@15331.4]
  wire [1534:0] _T_2292; // @[NV_NVDLA_CSC_wl.scala 744:42:@15331.4]
  wire [7:0] _T_2293; // @[NV_NVDLA_CSC_wl.scala 747:45:@15333.6]
  wire [7:0] _T_2294; // @[NV_NVDLA_CSC_wl.scala 747:45:@15335.6]
  wire [7:0] _T_2295; // @[NV_NVDLA_CSC_wl.scala 747:45:@15337.6]
  wire [7:0] _T_2296; // @[NV_NVDLA_CSC_wl.scala 747:45:@15339.6]
  wire [7:0] _T_2297; // @[NV_NVDLA_CSC_wl.scala 747:45:@15341.6]
  wire [7:0] _T_2298; // @[NV_NVDLA_CSC_wl.scala 747:45:@15343.6]
  wire [7:0] _T_2299; // @[NV_NVDLA_CSC_wl.scala 747:45:@15345.6]
  wire [7:0] _T_2300; // @[NV_NVDLA_CSC_wl.scala 747:45:@15347.6]
  wire [7:0] _T_2301; // @[NV_NVDLA_CSC_wl.scala 747:45:@15349.6]
  wire [7:0] _T_2302; // @[NV_NVDLA_CSC_wl.scala 747:45:@15351.6]
  wire [7:0] _T_2303; // @[NV_NVDLA_CSC_wl.scala 747:45:@15353.6]
  wire [7:0] _T_2304; // @[NV_NVDLA_CSC_wl.scala 747:45:@15355.6]
  wire [7:0] _T_2305; // @[NV_NVDLA_CSC_wl.scala 747:45:@15357.6]
  wire [7:0] _T_2306; // @[NV_NVDLA_CSC_wl.scala 747:45:@15359.6]
  wire [7:0] _T_2307; // @[NV_NVDLA_CSC_wl.scala 747:45:@15361.6]
  wire [7:0] _T_2308; // @[NV_NVDLA_CSC_wl.scala 747:45:@15363.6]
  wire [7:0] _T_2309; // @[NV_NVDLA_CSC_wl.scala 747:45:@15365.6]
  wire [7:0] _T_2310; // @[NV_NVDLA_CSC_wl.scala 747:45:@15367.6]
  wire [7:0] _T_2311; // @[NV_NVDLA_CSC_wl.scala 747:45:@15369.6]
  wire [7:0] _T_2312; // @[NV_NVDLA_CSC_wl.scala 747:45:@15371.6]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_wl.scala 747:45:@15373.6]
  wire [7:0] _T_2314; // @[NV_NVDLA_CSC_wl.scala 747:45:@15375.6]
  wire [7:0] _T_2315; // @[NV_NVDLA_CSC_wl.scala 747:45:@15377.6]
  wire [7:0] _T_2316; // @[NV_NVDLA_CSC_wl.scala 747:45:@15379.6]
  wire [7:0] _T_2317; // @[NV_NVDLA_CSC_wl.scala 747:45:@15381.6]
  wire [7:0] _T_2318; // @[NV_NVDLA_CSC_wl.scala 747:45:@15383.6]
  wire [7:0] _T_2319; // @[NV_NVDLA_CSC_wl.scala 747:45:@15385.6]
  wire [7:0] _T_2320; // @[NV_NVDLA_CSC_wl.scala 747:45:@15387.6]
  wire [7:0] _T_2321; // @[NV_NVDLA_CSC_wl.scala 747:45:@15389.6]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_wl.scala 747:45:@15391.6]
  wire [7:0] _T_2323; // @[NV_NVDLA_CSC_wl.scala 747:45:@15393.6]
  wire [7:0] _T_2324; // @[NV_NVDLA_CSC_wl.scala 747:45:@15395.6]
  wire [7:0] _T_2325; // @[NV_NVDLA_CSC_wl.scala 747:45:@15397.6]
  wire [7:0] _T_2326; // @[NV_NVDLA_CSC_wl.scala 747:45:@15399.6]
  wire [7:0] _T_2327; // @[NV_NVDLA_CSC_wl.scala 747:45:@15401.6]
  wire [7:0] _T_2328; // @[NV_NVDLA_CSC_wl.scala 747:45:@15403.6]
  wire [7:0] _T_2329; // @[NV_NVDLA_CSC_wl.scala 747:45:@15405.6]
  wire [7:0] _T_2330; // @[NV_NVDLA_CSC_wl.scala 747:45:@15407.6]
  wire [7:0] _T_2331; // @[NV_NVDLA_CSC_wl.scala 747:45:@15409.6]
  wire [7:0] _T_2332; // @[NV_NVDLA_CSC_wl.scala 747:45:@15411.6]
  wire [7:0] _T_2333; // @[NV_NVDLA_CSC_wl.scala 747:45:@15413.6]
  wire [7:0] _T_2334; // @[NV_NVDLA_CSC_wl.scala 747:45:@15415.6]
  wire [7:0] _T_2335; // @[NV_NVDLA_CSC_wl.scala 747:45:@15417.6]
  wire [7:0] _T_2336; // @[NV_NVDLA_CSC_wl.scala 747:45:@15419.6]
  wire [7:0] _T_2337; // @[NV_NVDLA_CSC_wl.scala 747:45:@15421.6]
  wire [7:0] _T_2338; // @[NV_NVDLA_CSC_wl.scala 747:45:@15423.6]
  wire [7:0] _T_2339; // @[NV_NVDLA_CSC_wl.scala 747:45:@15425.6]
  wire [7:0] _T_2340; // @[NV_NVDLA_CSC_wl.scala 747:45:@15427.6]
  wire [7:0] _T_2341; // @[NV_NVDLA_CSC_wl.scala 747:45:@15429.6]
  wire [7:0] _T_2342; // @[NV_NVDLA_CSC_wl.scala 747:45:@15431.6]
  wire [7:0] _T_2343; // @[NV_NVDLA_CSC_wl.scala 747:45:@15433.6]
  wire [7:0] _T_2344; // @[NV_NVDLA_CSC_wl.scala 747:45:@15435.6]
  wire [7:0] _T_2345; // @[NV_NVDLA_CSC_wl.scala 747:45:@15437.6]
  wire [7:0] _T_2346; // @[NV_NVDLA_CSC_wl.scala 747:45:@15439.6]
  wire [7:0] _T_2347; // @[NV_NVDLA_CSC_wl.scala 747:45:@15441.6]
  wire [7:0] _T_2348; // @[NV_NVDLA_CSC_wl.scala 747:45:@15443.6]
  wire [7:0] _T_2349; // @[NV_NVDLA_CSC_wl.scala 747:45:@15445.6]
  wire [7:0] _T_2350; // @[NV_NVDLA_CSC_wl.scala 747:45:@15447.6]
  wire [7:0] _T_2351; // @[NV_NVDLA_CSC_wl.scala 747:45:@15449.6]
  wire [7:0] _T_2352; // @[NV_NVDLA_CSC_wl.scala 747:45:@15451.6]
  wire [7:0] _T_2353; // @[NV_NVDLA_CSC_wl.scala 747:45:@15453.6]
  wire [7:0] _T_2354; // @[NV_NVDLA_CSC_wl.scala 747:45:@15455.6]
  wire [7:0] _T_2355; // @[NV_NVDLA_CSC_wl.scala 747:45:@15457.6]
  wire [7:0] _T_2356; // @[NV_NVDLA_CSC_wl.scala 747:45:@15459.6]
  wire [7:0] _GEN_79; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_80; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_81; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_82; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_83; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_84; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_85; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_86; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_87; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_88; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_89; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_90; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_91; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_92; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_93; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_94; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_95; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_96; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_97; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_98; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_99; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_100; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_101; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_102; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_103; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_104; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_106; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_107; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_108; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_109; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_110; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_111; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_112; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_113; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_114; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_115; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_116; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_117; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_118; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_119; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_120; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_121; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_122; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_123; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_124; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_125; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_126; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_127; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_128; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_129; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_130; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_131; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_132; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_133; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_134; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_135; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_136; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_137; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_138; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_139; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_140; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  reg  _T_2359; // @[NV_NVDLA_CSC_wl.scala 753:41:@15462.4]
  reg [31:0] _RAND_161;
  reg [31:0] _T_2362; // @[NV_NVDLA_CSC_wl.scala 754:32:@15463.4]
  reg [31:0] _RAND_162;
  wire [30:0] _T_2364; // @[NV_NVDLA_CSC_wl.scala 757:41:@15464.4]
  wire  _T_2365; // @[NV_NVDLA_CSC_wl.scala 757:77:@15465.4]
  wire [31:0] _T_2366; // @[Cat.scala 30:58:@15466.4]
  wire [31:0] _T_2367; // @[NV_NVDLA_CSC_wl.scala 756:27:@15467.4]
  wire  _GEN_143; // @[NV_NVDLA_CSC_wl.scala 759:27:@15468.4]
  wire [31:0] _GEN_144; // @[NV_NVDLA_CSC_wl.scala 759:27:@15468.4]
  reg  _T_2472; // @[NV_NVDLA_CSC_wl.scala 767:39:@15569.4]
  reg [31:0] _RAND_163;
  reg  _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_164;
  reg  _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_165;
  reg  _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_166;
  reg  _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_167;
  reg  _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_168;
  reg  _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_169;
  reg  _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_170;
  reg  _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_171;
  reg  _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_172;
  reg  _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_173;
  reg  _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_174;
  reg  _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_175;
  reg  _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_176;
  reg  _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_177;
  reg  _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_178;
  reg  _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_179;
  reg  _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_180;
  reg  _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_181;
  reg  _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_182;
  reg  _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_183;
  reg  _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_184;
  reg  _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_185;
  reg  _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_186;
  reg  _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_187;
  reg  _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_188;
  reg  _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_189;
  reg  _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_190;
  reg  _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_191;
  reg  _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_192;
  reg  _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_193;
  reg  _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_194;
  reg  _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_195;
  reg  _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_196;
  reg  _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_197;
  reg  _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_198;
  reg  _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_199;
  reg  _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_200;
  reg  _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_201;
  reg  _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_202;
  reg  _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_203;
  reg  _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_204;
  reg  _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_205;
  reg  _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_206;
  reg  _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_207;
  reg  _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_208;
  reg  _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_209;
  reg  _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_210;
  reg  _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_211;
  reg  _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_212;
  reg  _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_213;
  reg  _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_214;
  reg  _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_215;
  reg  _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_216;
  reg  _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_217;
  reg  _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_218;
  reg  _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_219;
  reg  _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_220;
  reg  _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_221;
  reg  _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_222;
  reg  _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_223;
  reg  _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_224;
  reg  _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_225;
  reg  _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_226;
  reg  _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 768:33:@15635.4]
  reg [31:0] _RAND_227;
  reg [9:0] _T_2938; // @[NV_NVDLA_CSC_wl.scala 769:36:@15636.4]
  reg [31:0] _RAND_228;
  wire  _T_2939; // @[NV_NVDLA_CSC_wl.scala 773:86:@15639.6]
  wire  _T_2940; // @[NV_NVDLA_CSC_wl.scala 773:86:@15640.6]
  wire  _T_2941; // @[NV_NVDLA_CSC_wl.scala 773:86:@15641.6]
  wire  _T_2942; // @[NV_NVDLA_CSC_wl.scala 773:86:@15642.6]
  wire  _T_2943; // @[NV_NVDLA_CSC_wl.scala 773:86:@15643.6]
  wire  _T_2944; // @[NV_NVDLA_CSC_wl.scala 773:86:@15644.6]
  wire  _T_2945; // @[NV_NVDLA_CSC_wl.scala 773:86:@15645.6]
  wire  _T_2946; // @[NV_NVDLA_CSC_wl.scala 773:86:@15646.6]
  wire  _T_2947; // @[NV_NVDLA_CSC_wl.scala 773:86:@15647.6]
  wire  _T_2948; // @[NV_NVDLA_CSC_wl.scala 773:86:@15648.6]
  wire  _T_2949; // @[NV_NVDLA_CSC_wl.scala 773:86:@15649.6]
  wire  _T_2950; // @[NV_NVDLA_CSC_wl.scala 773:86:@15650.6]
  wire  _T_2951; // @[NV_NVDLA_CSC_wl.scala 773:86:@15651.6]
  wire  _T_2952; // @[NV_NVDLA_CSC_wl.scala 773:86:@15652.6]
  wire  _T_2953; // @[NV_NVDLA_CSC_wl.scala 773:86:@15653.6]
  wire  _T_2954; // @[NV_NVDLA_CSC_wl.scala 773:86:@15654.6]
  wire  _T_2955; // @[NV_NVDLA_CSC_wl.scala 773:86:@15655.6]
  wire  _T_2956; // @[NV_NVDLA_CSC_wl.scala 773:86:@15656.6]
  wire  _T_2957; // @[NV_NVDLA_CSC_wl.scala 773:86:@15657.6]
  wire  _T_2958; // @[NV_NVDLA_CSC_wl.scala 773:86:@15658.6]
  wire  _T_2959; // @[NV_NVDLA_CSC_wl.scala 773:86:@15659.6]
  wire  _T_2960; // @[NV_NVDLA_CSC_wl.scala 773:86:@15660.6]
  wire  _T_2961; // @[NV_NVDLA_CSC_wl.scala 773:86:@15661.6]
  wire  _T_2962; // @[NV_NVDLA_CSC_wl.scala 773:86:@15662.6]
  wire  _T_2963; // @[NV_NVDLA_CSC_wl.scala 773:86:@15663.6]
  wire  _T_2964; // @[NV_NVDLA_CSC_wl.scala 773:86:@15664.6]
  wire  _T_2965; // @[NV_NVDLA_CSC_wl.scala 773:86:@15665.6]
  wire  _T_2966; // @[NV_NVDLA_CSC_wl.scala 773:86:@15666.6]
  wire  _T_2967; // @[NV_NVDLA_CSC_wl.scala 773:86:@15667.6]
  wire  _T_2968; // @[NV_NVDLA_CSC_wl.scala 773:86:@15668.6]
  wire  _T_2969; // @[NV_NVDLA_CSC_wl.scala 773:86:@15669.6]
  wire  _T_2970; // @[NV_NVDLA_CSC_wl.scala 773:86:@15670.6]
  wire  _T_2971; // @[NV_NVDLA_CSC_wl.scala 773:86:@15671.6]
  wire  _T_2972; // @[NV_NVDLA_CSC_wl.scala 773:86:@15672.6]
  wire  _T_2973; // @[NV_NVDLA_CSC_wl.scala 773:86:@15673.6]
  wire  _T_2974; // @[NV_NVDLA_CSC_wl.scala 773:86:@15674.6]
  wire  _T_2975; // @[NV_NVDLA_CSC_wl.scala 773:86:@15675.6]
  wire  _T_2976; // @[NV_NVDLA_CSC_wl.scala 773:86:@15676.6]
  wire  _T_2977; // @[NV_NVDLA_CSC_wl.scala 773:86:@15677.6]
  wire  _T_2978; // @[NV_NVDLA_CSC_wl.scala 773:86:@15678.6]
  wire  _T_2979; // @[NV_NVDLA_CSC_wl.scala 773:86:@15679.6]
  wire  _T_2980; // @[NV_NVDLA_CSC_wl.scala 773:86:@15680.6]
  wire  _T_2981; // @[NV_NVDLA_CSC_wl.scala 773:86:@15681.6]
  wire  _T_2982; // @[NV_NVDLA_CSC_wl.scala 773:86:@15682.6]
  wire  _T_2983; // @[NV_NVDLA_CSC_wl.scala 773:86:@15683.6]
  wire  _T_2984; // @[NV_NVDLA_CSC_wl.scala 773:86:@15684.6]
  wire  _T_2985; // @[NV_NVDLA_CSC_wl.scala 773:86:@15685.6]
  wire  _T_2986; // @[NV_NVDLA_CSC_wl.scala 773:86:@15686.6]
  wire  _T_2987; // @[NV_NVDLA_CSC_wl.scala 773:86:@15687.6]
  wire  _T_2988; // @[NV_NVDLA_CSC_wl.scala 773:86:@15688.6]
  wire  _T_2989; // @[NV_NVDLA_CSC_wl.scala 773:86:@15689.6]
  wire  _T_2990; // @[NV_NVDLA_CSC_wl.scala 773:86:@15690.6]
  wire  _T_2991; // @[NV_NVDLA_CSC_wl.scala 773:86:@15691.6]
  wire  _T_2992; // @[NV_NVDLA_CSC_wl.scala 773:86:@15692.6]
  wire  _T_2993; // @[NV_NVDLA_CSC_wl.scala 773:86:@15693.6]
  wire  _T_2994; // @[NV_NVDLA_CSC_wl.scala 773:86:@15694.6]
  wire  _T_2995; // @[NV_NVDLA_CSC_wl.scala 773:86:@15695.6]
  wire  _T_2996; // @[NV_NVDLA_CSC_wl.scala 773:86:@15696.6]
  wire  _T_2997; // @[NV_NVDLA_CSC_wl.scala 773:86:@15697.6]
  wire  _T_2998; // @[NV_NVDLA_CSC_wl.scala 773:86:@15698.6]
  wire  _T_2999; // @[NV_NVDLA_CSC_wl.scala 773:86:@15699.6]
  wire  _T_3000; // @[NV_NVDLA_CSC_wl.scala 773:86:@15700.6]
  wire  _T_3001; // @[NV_NVDLA_CSC_wl.scala 773:86:@15701.6]
  wire  _T_3002; // @[NV_NVDLA_CSC_wl.scala 773:86:@15702.6]
  wire  _GEN_145; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_146; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_147; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_148; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_149; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_150; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_151; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_152; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_153; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_154; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_155; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  wire [9:0] _T_3076; // @[Bitwise.scala 72:12:@15834.4]
  wire  _T_3077; // @[Bitwise.scala 72:15:@16002.4]
  wire [15:0] _T_3080; // @[Bitwise.scala 72:12:@16003.4]
  wire [7:0] _T_3087; // @[NV_NVDLA_CSC_wl.scala 794:92:@16010.4]
  wire [15:0] _T_3095; // @[NV_NVDLA_CSC_wl.scala 794:92:@16018.4]
  wire [7:0] _T_3102; // @[NV_NVDLA_CSC_wl.scala 794:92:@16025.4]
  wire [31:0] _T_3111; // @[NV_NVDLA_CSC_wl.scala 794:92:@16034.4]
  wire [15:0] _T_3112; // @[NV_NVDLA_CSC_wl.scala 794:99:@16035.4]
  wire [15:0] _T_3113; // @[NV_NVDLA_CSC_wl.scala 794:71:@16036.4]
  wire [15:0] _T_3149; // @[NV_NVDLA_CSC_wl.scala 795:99:@16070.4]
  wire [15:0] _T_3150; // @[NV_NVDLA_CSC_wl.scala 795:71:@16071.4]
  wire  _T_3152; // @[NV_NVDLA_CSC_wl.scala 796:49:@16072.4]
  wire  _T_3154; // @[NV_NVDLA_CSC_wl.scala 797:49:@16073.4]
  reg  _T_3157; // @[NV_NVDLA_CSC_wl.scala 799:39:@16074.4]
  reg [31:0] _RAND_229;
  reg  _T_3160; // @[NV_NVDLA_CSC_wl.scala 800:39:@16075.4]
  reg [31:0] _RAND_230;
  reg  _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_231;
  reg  _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_232;
  reg  _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_233;
  reg  _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_234;
  reg  _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_235;
  reg  _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_236;
  reg  _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_237;
  reg  _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_238;
  reg  _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_239;
  reg  _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_240;
  reg  _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_241;
  reg  _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_242;
  reg  _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_243;
  reg  _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_244;
  reg  _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_245;
  reg  _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_246;
  reg  _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_247;
  reg  _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_248;
  reg  _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_249;
  reg  _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_250;
  reg  _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_251;
  reg  _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_252;
  reg  _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_253;
  reg  _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_254;
  reg  _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_255;
  reg  _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_256;
  reg  _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_257;
  reg  _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_258;
  reg  _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_259;
  reg  _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_260;
  reg  _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_261;
  reg  _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_262;
  reg  _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_263;
  reg  _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_264;
  reg  _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_265;
  reg  _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_266;
  reg  _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_267;
  reg  _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_268;
  reg  _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_269;
  reg  _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_270;
  reg  _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_271;
  reg  _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_272;
  reg  _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_273;
  reg  _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_274;
  reg  _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_275;
  reg  _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_276;
  reg  _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_277;
  reg  _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_278;
  reg  _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_279;
  reg  _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_280;
  reg  _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_281;
  reg  _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_282;
  reg  _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_283;
  reg  _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_284;
  reg  _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_285;
  reg  _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_286;
  reg  _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_287;
  reg  _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_288;
  reg  _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_289;
  reg  _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_290;
  reg  _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_291;
  reg  _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_292;
  reg  _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_293;
  reg  _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 801:39:@16141.4]
  reg [31:0] _RAND_294;
  reg  _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_295;
  reg  _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_296;
  reg  _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_297;
  reg  _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_298;
  reg  _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_299;
  reg  _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_300;
  reg  _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_301;
  reg  _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_302;
  reg  _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_303;
  reg  _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_304;
  reg  _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_305;
  reg  _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_306;
  reg  _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_307;
  reg  _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_308;
  reg  _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_309;
  reg  _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_310;
  reg  _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_311;
  reg  _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_312;
  reg  _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_313;
  reg  _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_314;
  reg  _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_315;
  reg  _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_316;
  reg  _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_317;
  reg  _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_318;
  reg  _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_319;
  reg  _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_320;
  reg  _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_321;
  reg  _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_322;
  reg  _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_323;
  reg  _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_324;
  reg  _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_325;
  reg  _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_326;
  reg  _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_327;
  reg  _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_328;
  reg  _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_329;
  reg  _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_330;
  reg  _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_331;
  reg  _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_332;
  reg  _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_333;
  reg  _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_334;
  reg  _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_335;
  reg  _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_336;
  reg  _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_337;
  reg  _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_338;
  reg  _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_339;
  reg  _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_340;
  reg  _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_341;
  reg  _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_342;
  reg  _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_343;
  reg  _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_344;
  reg  _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_345;
  reg  _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_346;
  reg  _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_347;
  reg  _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_348;
  reg  _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_349;
  reg  _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_350;
  reg  _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_351;
  reg  _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_352;
  reg  _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_353;
  reg  _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_354;
  reg  _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_355;
  reg  _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_356;
  reg  _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_357;
  reg  _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 802:39:@16207.4]
  reg [31:0] _RAND_358;
  reg  _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_359;
  reg  _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_360;
  reg  _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_361;
  reg  _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_362;
  reg  _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_363;
  reg  _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_364;
  reg  _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_365;
  reg  _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_366;
  reg  _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_367;
  reg  _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_368;
  reg  _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_369;
  reg  _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_370;
  reg  _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_371;
  reg  _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_372;
  reg  _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_373;
  reg  _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 803:38:@16225.4]
  reg [31:0] _RAND_374;
  reg  _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_375;
  reg  _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_376;
  reg  _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_377;
  reg  _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_378;
  reg  _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_379;
  reg  _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_380;
  reg  _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_381;
  reg  _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_382;
  reg  _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_383;
  reg  _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_384;
  reg  _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_385;
  reg  _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_386;
  reg  _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_387;
  reg  _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_388;
  reg  _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_389;
  reg  _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 804:38:@16243.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4344_0; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4344_1; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4344_2; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4344_3; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4344_4; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4344_5; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4344_6; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4344_7; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4344_8; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4344_9; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4344_10; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4344_11; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4344_12; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4344_13; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4344_14; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4344_15; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4344_16; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4344_17; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4344_18; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4344_19; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4344_20; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_411;
  reg [7:0] _T_4344_21; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_412;
  reg [7:0] _T_4344_22; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_413;
  reg [7:0] _T_4344_23; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_414;
  reg [7:0] _T_4344_24; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_415;
  reg [7:0] _T_4344_25; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_416;
  reg [7:0] _T_4344_26; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_417;
  reg [7:0] _T_4344_27; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_418;
  reg [7:0] _T_4344_28; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_419;
  reg [7:0] _T_4344_29; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_420;
  reg [7:0] _T_4344_30; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_421;
  reg [7:0] _T_4344_31; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_422;
  reg [7:0] _T_4344_32; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_423;
  reg [7:0] _T_4344_33; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_424;
  reg [7:0] _T_4344_34; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_425;
  reg [7:0] _T_4344_35; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_426;
  reg [7:0] _T_4344_36; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_427;
  reg [7:0] _T_4344_37; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_428;
  reg [7:0] _T_4344_38; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_429;
  reg [7:0] _T_4344_39; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_430;
  reg [7:0] _T_4344_40; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_431;
  reg [7:0] _T_4344_41; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_432;
  reg [7:0] _T_4344_42; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_433;
  reg [7:0] _T_4344_43; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_434;
  reg [7:0] _T_4344_44; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_435;
  reg [7:0] _T_4344_45; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_436;
  reg [7:0] _T_4344_46; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_437;
  reg [7:0] _T_4344_47; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_438;
  reg [7:0] _T_4344_48; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_439;
  reg [7:0] _T_4344_49; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_440;
  reg [7:0] _T_4344_50; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_441;
  reg [7:0] _T_4344_51; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_442;
  reg [7:0] _T_4344_52; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_443;
  reg [7:0] _T_4344_53; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_444;
  reg [7:0] _T_4344_54; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_445;
  reg [7:0] _T_4344_55; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_446;
  reg [7:0] _T_4344_56; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_447;
  reg [7:0] _T_4344_57; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_448;
  reg [7:0] _T_4344_58; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_449;
  reg [7:0] _T_4344_59; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_450;
  reg [7:0] _T_4344_60; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_451;
  reg [7:0] _T_4344_61; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_452;
  reg [7:0] _T_4344_62; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_453;
  reg [7:0] _T_4344_63; // @[NV_NVDLA_CSC_wl.scala 805:35:@16244.4]
  reg [31:0] _RAND_454;
  reg [7:0] _T_4414_0; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_455;
  reg [7:0] _T_4414_1; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_456;
  reg [7:0] _T_4414_2; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_457;
  reg [7:0] _T_4414_3; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_458;
  reg [7:0] _T_4414_4; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_459;
  reg [7:0] _T_4414_5; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_460;
  reg [7:0] _T_4414_6; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_461;
  reg [7:0] _T_4414_7; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_462;
  reg [7:0] _T_4414_8; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_463;
  reg [7:0] _T_4414_9; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_464;
  reg [7:0] _T_4414_10; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_465;
  reg [7:0] _T_4414_11; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_466;
  reg [7:0] _T_4414_12; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_467;
  reg [7:0] _T_4414_13; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_468;
  reg [7:0] _T_4414_14; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_469;
  reg [7:0] _T_4414_15; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_470;
  reg [7:0] _T_4414_16; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_471;
  reg [7:0] _T_4414_17; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_472;
  reg [7:0] _T_4414_18; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_473;
  reg [7:0] _T_4414_19; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_474;
  reg [7:0] _T_4414_20; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_475;
  reg [7:0] _T_4414_21; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_476;
  reg [7:0] _T_4414_22; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_477;
  reg [7:0] _T_4414_23; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_478;
  reg [7:0] _T_4414_24; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_479;
  reg [7:0] _T_4414_25; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_480;
  reg [7:0] _T_4414_26; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_481;
  reg [7:0] _T_4414_27; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_482;
  reg [7:0] _T_4414_28; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_483;
  reg [7:0] _T_4414_29; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_484;
  reg [7:0] _T_4414_30; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_485;
  reg [7:0] _T_4414_31; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_486;
  reg [7:0] _T_4414_32; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_487;
  reg [7:0] _T_4414_33; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_488;
  reg [7:0] _T_4414_34; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_489;
  reg [7:0] _T_4414_35; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_490;
  reg [7:0] _T_4414_36; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_491;
  reg [7:0] _T_4414_37; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_492;
  reg [7:0] _T_4414_38; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_493;
  reg [7:0] _T_4414_39; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_494;
  reg [7:0] _T_4414_40; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_495;
  reg [7:0] _T_4414_41; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_496;
  reg [7:0] _T_4414_42; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_497;
  reg [7:0] _T_4414_43; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_498;
  reg [7:0] _T_4414_44; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_499;
  reg [7:0] _T_4414_45; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_500;
  reg [7:0] _T_4414_46; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_501;
  reg [7:0] _T_4414_47; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_502;
  reg [7:0] _T_4414_48; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_503;
  reg [7:0] _T_4414_49; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_504;
  reg [7:0] _T_4414_50; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_505;
  reg [7:0] _T_4414_51; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_506;
  reg [7:0] _T_4414_52; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_507;
  reg [7:0] _T_4414_53; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_508;
  reg [7:0] _T_4414_54; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_509;
  reg [7:0] _T_4414_55; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_510;
  reg [7:0] _T_4414_56; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_511;
  reg [7:0] _T_4414_57; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_512;
  reg [7:0] _T_4414_58; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_513;
  reg [7:0] _T_4414_59; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_514;
  reg [7:0] _T_4414_60; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_515;
  reg [7:0] _T_4414_61; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_516;
  reg [7:0] _T_4414_62; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_517;
  reg [7:0] _T_4414_63; // @[NV_NVDLA_CSC_wl.scala 806:35:@16245.4]
  reg [31:0] _RAND_518;
  wire  _T_4481; // @[NV_NVDLA_CSC_wl.scala 807:91:@16246.4]
  wire  _T_4482; // @[NV_NVDLA_CSC_wl.scala 807:97:@16247.4]
  wire  _T_4483; // @[NV_NVDLA_CSC_wl.scala 807:91:@16248.4]
  wire  _T_4484; // @[NV_NVDLA_CSC_wl.scala 807:97:@16249.4]
  wire  _T_4485; // @[NV_NVDLA_CSC_wl.scala 807:91:@16250.4]
  wire  _T_4486; // @[NV_NVDLA_CSC_wl.scala 807:97:@16251.4]
  wire  _T_4487; // @[NV_NVDLA_CSC_wl.scala 807:91:@16252.4]
  wire  _T_4488; // @[NV_NVDLA_CSC_wl.scala 807:97:@16253.4]
  wire  _T_4489; // @[NV_NVDLA_CSC_wl.scala 807:91:@16254.4]
  wire  _T_4490; // @[NV_NVDLA_CSC_wl.scala 807:97:@16255.4]
  wire  _T_4491; // @[NV_NVDLA_CSC_wl.scala 807:91:@16256.4]
  wire  _T_4492; // @[NV_NVDLA_CSC_wl.scala 807:97:@16257.4]
  wire  _T_4493; // @[NV_NVDLA_CSC_wl.scala 807:91:@16258.4]
  wire  _T_4494; // @[NV_NVDLA_CSC_wl.scala 807:97:@16259.4]
  wire  _T_4495; // @[NV_NVDLA_CSC_wl.scala 807:91:@16260.4]
  wire  _T_4496; // @[NV_NVDLA_CSC_wl.scala 807:97:@16261.4]
  wire  _T_4497; // @[NV_NVDLA_CSC_wl.scala 807:91:@16262.4]
  wire  _T_4498; // @[NV_NVDLA_CSC_wl.scala 807:97:@16263.4]
  wire  _T_4499; // @[NV_NVDLA_CSC_wl.scala 807:91:@16264.4]
  wire  _T_4500; // @[NV_NVDLA_CSC_wl.scala 807:97:@16265.4]
  wire  _T_4501; // @[NV_NVDLA_CSC_wl.scala 807:91:@16266.4]
  wire  _T_4502; // @[NV_NVDLA_CSC_wl.scala 807:97:@16267.4]
  wire  _T_4503; // @[NV_NVDLA_CSC_wl.scala 807:91:@16268.4]
  wire  _T_4504; // @[NV_NVDLA_CSC_wl.scala 807:97:@16269.4]
  wire  _T_4505; // @[NV_NVDLA_CSC_wl.scala 807:91:@16270.4]
  wire  _T_4506; // @[NV_NVDLA_CSC_wl.scala 807:97:@16271.4]
  wire  _T_4507; // @[NV_NVDLA_CSC_wl.scala 807:91:@16272.4]
  wire  _T_4508; // @[NV_NVDLA_CSC_wl.scala 807:97:@16273.4]
  wire  _T_4509; // @[NV_NVDLA_CSC_wl.scala 807:91:@16274.4]
  wire  _T_4510; // @[NV_NVDLA_CSC_wl.scala 807:97:@16275.4]
  wire  _T_4511; // @[NV_NVDLA_CSC_wl.scala 807:91:@16276.4]
  wire  _T_4512; // @[NV_NVDLA_CSC_wl.scala 807:97:@16277.4]
  wire  _T_4513; // @[NV_NVDLA_CSC_wl.scala 807:91:@16278.4]
  wire  _T_4514; // @[NV_NVDLA_CSC_wl.scala 807:97:@16279.4]
  wire  _T_4515; // @[NV_NVDLA_CSC_wl.scala 807:91:@16280.4]
  wire  _T_4516; // @[NV_NVDLA_CSC_wl.scala 807:97:@16281.4]
  wire  _T_4517; // @[NV_NVDLA_CSC_wl.scala 807:91:@16282.4]
  wire  _T_4518; // @[NV_NVDLA_CSC_wl.scala 807:97:@16283.4]
  wire  _T_4519; // @[NV_NVDLA_CSC_wl.scala 807:91:@16284.4]
  wire  _T_4520; // @[NV_NVDLA_CSC_wl.scala 807:97:@16285.4]
  wire  _T_4521; // @[NV_NVDLA_CSC_wl.scala 807:91:@16286.4]
  wire  _T_4522; // @[NV_NVDLA_CSC_wl.scala 807:97:@16287.4]
  wire  _T_4523; // @[NV_NVDLA_CSC_wl.scala 807:91:@16288.4]
  wire  _T_4524; // @[NV_NVDLA_CSC_wl.scala 807:97:@16289.4]
  wire  _T_4525; // @[NV_NVDLA_CSC_wl.scala 807:91:@16290.4]
  wire  _T_4526; // @[NV_NVDLA_CSC_wl.scala 807:97:@16291.4]
  wire  _T_4527; // @[NV_NVDLA_CSC_wl.scala 807:91:@16292.4]
  wire  _T_4528; // @[NV_NVDLA_CSC_wl.scala 807:97:@16293.4]
  wire  _T_4529; // @[NV_NVDLA_CSC_wl.scala 807:91:@16294.4]
  wire  _T_4530; // @[NV_NVDLA_CSC_wl.scala 807:97:@16295.4]
  wire  _T_4531; // @[NV_NVDLA_CSC_wl.scala 807:91:@16296.4]
  wire  _T_4532; // @[NV_NVDLA_CSC_wl.scala 807:97:@16297.4]
  wire  _T_4533; // @[NV_NVDLA_CSC_wl.scala 807:91:@16298.4]
  wire  _T_4534; // @[NV_NVDLA_CSC_wl.scala 807:97:@16299.4]
  wire  _T_4535; // @[NV_NVDLA_CSC_wl.scala 807:91:@16300.4]
  wire  _T_4536; // @[NV_NVDLA_CSC_wl.scala 807:97:@16301.4]
  wire  _T_4537; // @[NV_NVDLA_CSC_wl.scala 807:91:@16302.4]
  wire  _T_4538; // @[NV_NVDLA_CSC_wl.scala 807:97:@16303.4]
  wire  _T_4539; // @[NV_NVDLA_CSC_wl.scala 807:91:@16304.4]
  wire  _T_4540; // @[NV_NVDLA_CSC_wl.scala 807:97:@16305.4]
  wire  _T_4541; // @[NV_NVDLA_CSC_wl.scala 807:91:@16306.4]
  wire  _T_4542; // @[NV_NVDLA_CSC_wl.scala 807:97:@16307.4]
  wire  _T_4543; // @[NV_NVDLA_CSC_wl.scala 807:91:@16308.4]
  wire  _T_4544; // @[NV_NVDLA_CSC_wl.scala 807:97:@16309.4]
  wire  _T_4545; // @[NV_NVDLA_CSC_wl.scala 807:91:@16310.4]
  wire  _T_4546; // @[NV_NVDLA_CSC_wl.scala 807:97:@16311.4]
  wire  _T_4547; // @[NV_NVDLA_CSC_wl.scala 807:91:@16312.4]
  wire  _T_4548; // @[NV_NVDLA_CSC_wl.scala 807:97:@16313.4]
  wire  _T_4549; // @[NV_NVDLA_CSC_wl.scala 807:91:@16314.4]
  wire  _T_4550; // @[NV_NVDLA_CSC_wl.scala 807:97:@16315.4]
  wire  _T_4551; // @[NV_NVDLA_CSC_wl.scala 807:91:@16316.4]
  wire  _T_4552; // @[NV_NVDLA_CSC_wl.scala 807:97:@16317.4]
  wire  _T_4553; // @[NV_NVDLA_CSC_wl.scala 807:91:@16318.4]
  wire  _T_4554; // @[NV_NVDLA_CSC_wl.scala 807:97:@16319.4]
  wire  _T_4555; // @[NV_NVDLA_CSC_wl.scala 807:91:@16320.4]
  wire  _T_4556; // @[NV_NVDLA_CSC_wl.scala 807:97:@16321.4]
  wire  _T_4557; // @[NV_NVDLA_CSC_wl.scala 807:91:@16322.4]
  wire  _T_4558; // @[NV_NVDLA_CSC_wl.scala 807:97:@16323.4]
  wire  _T_4559; // @[NV_NVDLA_CSC_wl.scala 807:91:@16324.4]
  wire  _T_4560; // @[NV_NVDLA_CSC_wl.scala 807:97:@16325.4]
  wire  _T_4561; // @[NV_NVDLA_CSC_wl.scala 807:91:@16326.4]
  wire  _T_4562; // @[NV_NVDLA_CSC_wl.scala 807:97:@16327.4]
  wire  _T_4563; // @[NV_NVDLA_CSC_wl.scala 807:91:@16328.4]
  wire  _T_4564; // @[NV_NVDLA_CSC_wl.scala 807:97:@16329.4]
  wire  _T_4565; // @[NV_NVDLA_CSC_wl.scala 807:91:@16330.4]
  wire  _T_4566; // @[NV_NVDLA_CSC_wl.scala 807:97:@16331.4]
  wire  _T_4567; // @[NV_NVDLA_CSC_wl.scala 807:91:@16332.4]
  wire  _T_4568; // @[NV_NVDLA_CSC_wl.scala 807:97:@16333.4]
  wire  _T_4569; // @[NV_NVDLA_CSC_wl.scala 807:91:@16334.4]
  wire  _T_4570; // @[NV_NVDLA_CSC_wl.scala 807:97:@16335.4]
  wire  _T_4571; // @[NV_NVDLA_CSC_wl.scala 807:91:@16336.4]
  wire  _T_4572; // @[NV_NVDLA_CSC_wl.scala 807:97:@16337.4]
  wire  _T_4573; // @[NV_NVDLA_CSC_wl.scala 807:91:@16338.4]
  wire  _T_4574; // @[NV_NVDLA_CSC_wl.scala 807:97:@16339.4]
  wire  _T_4575; // @[NV_NVDLA_CSC_wl.scala 807:91:@16340.4]
  wire  _T_4576; // @[NV_NVDLA_CSC_wl.scala 807:97:@16341.4]
  wire  _T_4577; // @[NV_NVDLA_CSC_wl.scala 807:91:@16342.4]
  wire  _T_4578; // @[NV_NVDLA_CSC_wl.scala 807:97:@16343.4]
  wire  _T_4579; // @[NV_NVDLA_CSC_wl.scala 807:91:@16344.4]
  wire  _T_4580; // @[NV_NVDLA_CSC_wl.scala 807:97:@16345.4]
  wire  _T_4581; // @[NV_NVDLA_CSC_wl.scala 807:91:@16346.4]
  wire  _T_4582; // @[NV_NVDLA_CSC_wl.scala 807:97:@16347.4]
  wire  _T_4583; // @[NV_NVDLA_CSC_wl.scala 807:91:@16348.4]
  wire  _T_4584; // @[NV_NVDLA_CSC_wl.scala 807:97:@16349.4]
  wire  _T_4585; // @[NV_NVDLA_CSC_wl.scala 807:91:@16350.4]
  wire  _T_4586; // @[NV_NVDLA_CSC_wl.scala 807:97:@16351.4]
  wire  _T_4587; // @[NV_NVDLA_CSC_wl.scala 807:91:@16352.4]
  wire  _T_4588; // @[NV_NVDLA_CSC_wl.scala 807:97:@16353.4]
  wire  _T_4589; // @[NV_NVDLA_CSC_wl.scala 807:91:@16354.4]
  wire  _T_4590; // @[NV_NVDLA_CSC_wl.scala 807:97:@16355.4]
  wire  _T_4591; // @[NV_NVDLA_CSC_wl.scala 807:91:@16356.4]
  wire  _T_4592; // @[NV_NVDLA_CSC_wl.scala 807:97:@16357.4]
  wire  _T_4593; // @[NV_NVDLA_CSC_wl.scala 807:91:@16358.4]
  wire  _T_4594; // @[NV_NVDLA_CSC_wl.scala 807:97:@16359.4]
  wire  _T_4595; // @[NV_NVDLA_CSC_wl.scala 807:91:@16360.4]
  wire  _T_4596; // @[NV_NVDLA_CSC_wl.scala 807:97:@16361.4]
  wire  _T_4597; // @[NV_NVDLA_CSC_wl.scala 807:91:@16362.4]
  wire  _T_4598; // @[NV_NVDLA_CSC_wl.scala 807:97:@16363.4]
  wire  _T_4599; // @[NV_NVDLA_CSC_wl.scala 807:91:@16364.4]
  wire  _T_4600; // @[NV_NVDLA_CSC_wl.scala 807:97:@16365.4]
  wire  _T_4601; // @[NV_NVDLA_CSC_wl.scala 807:91:@16366.4]
  wire  _T_4602; // @[NV_NVDLA_CSC_wl.scala 807:97:@16367.4]
  wire  _T_4603; // @[NV_NVDLA_CSC_wl.scala 807:91:@16368.4]
  wire  _T_4604; // @[NV_NVDLA_CSC_wl.scala 807:97:@16369.4]
  wire  _T_4605; // @[NV_NVDLA_CSC_wl.scala 807:91:@16370.4]
  wire  _T_4606; // @[NV_NVDLA_CSC_wl.scala 807:97:@16371.4]
  wire  _T_4607; // @[NV_NVDLA_CSC_wl.scala 807:91:@16372.4]
  wire  _T_4608; // @[NV_NVDLA_CSC_wl.scala 807:97:@16373.4]
  wire  _T_4680; // @[NV_NVDLA_CSC_wl.scala 808:97:@16440.4]
  wire  _T_4682; // @[NV_NVDLA_CSC_wl.scala 808:97:@16442.4]
  wire  _T_4684; // @[NV_NVDLA_CSC_wl.scala 808:97:@16444.4]
  wire  _T_4686; // @[NV_NVDLA_CSC_wl.scala 808:97:@16446.4]
  wire  _T_4688; // @[NV_NVDLA_CSC_wl.scala 808:97:@16448.4]
  wire  _T_4690; // @[NV_NVDLA_CSC_wl.scala 808:97:@16450.4]
  wire  _T_4692; // @[NV_NVDLA_CSC_wl.scala 808:97:@16452.4]
  wire  _T_4694; // @[NV_NVDLA_CSC_wl.scala 808:97:@16454.4]
  wire  _T_4696; // @[NV_NVDLA_CSC_wl.scala 808:97:@16456.4]
  wire  _T_4698; // @[NV_NVDLA_CSC_wl.scala 808:97:@16458.4]
  wire  _T_4700; // @[NV_NVDLA_CSC_wl.scala 808:97:@16460.4]
  wire  _T_4702; // @[NV_NVDLA_CSC_wl.scala 808:97:@16462.4]
  wire  _T_4704; // @[NV_NVDLA_CSC_wl.scala 808:97:@16464.4]
  wire  _T_4706; // @[NV_NVDLA_CSC_wl.scala 808:97:@16466.4]
  wire  _T_4708; // @[NV_NVDLA_CSC_wl.scala 808:97:@16468.4]
  wire  _T_4710; // @[NV_NVDLA_CSC_wl.scala 808:97:@16470.4]
  wire  _T_4712; // @[NV_NVDLA_CSC_wl.scala 808:97:@16472.4]
  wire  _T_4714; // @[NV_NVDLA_CSC_wl.scala 808:97:@16474.4]
  wire  _T_4716; // @[NV_NVDLA_CSC_wl.scala 808:97:@16476.4]
  wire  _T_4718; // @[NV_NVDLA_CSC_wl.scala 808:97:@16478.4]
  wire  _T_4720; // @[NV_NVDLA_CSC_wl.scala 808:97:@16480.4]
  wire  _T_4722; // @[NV_NVDLA_CSC_wl.scala 808:97:@16482.4]
  wire  _T_4724; // @[NV_NVDLA_CSC_wl.scala 808:97:@16484.4]
  wire  _T_4726; // @[NV_NVDLA_CSC_wl.scala 808:97:@16486.4]
  wire  _T_4728; // @[NV_NVDLA_CSC_wl.scala 808:97:@16488.4]
  wire  _T_4730; // @[NV_NVDLA_CSC_wl.scala 808:97:@16490.4]
  wire  _T_4732; // @[NV_NVDLA_CSC_wl.scala 808:97:@16492.4]
  wire  _T_4734; // @[NV_NVDLA_CSC_wl.scala 808:97:@16494.4]
  wire  _T_4736; // @[NV_NVDLA_CSC_wl.scala 808:97:@16496.4]
  wire  _T_4738; // @[NV_NVDLA_CSC_wl.scala 808:97:@16498.4]
  wire  _T_4740; // @[NV_NVDLA_CSC_wl.scala 808:97:@16500.4]
  wire  _T_4742; // @[NV_NVDLA_CSC_wl.scala 808:97:@16502.4]
  wire  _T_4744; // @[NV_NVDLA_CSC_wl.scala 808:97:@16504.4]
  wire  _T_4746; // @[NV_NVDLA_CSC_wl.scala 808:97:@16506.4]
  wire  _T_4748; // @[NV_NVDLA_CSC_wl.scala 808:97:@16508.4]
  wire  _T_4750; // @[NV_NVDLA_CSC_wl.scala 808:97:@16510.4]
  wire  _T_4752; // @[NV_NVDLA_CSC_wl.scala 808:97:@16512.4]
  wire  _T_4754; // @[NV_NVDLA_CSC_wl.scala 808:97:@16514.4]
  wire  _T_4756; // @[NV_NVDLA_CSC_wl.scala 808:97:@16516.4]
  wire  _T_4758; // @[NV_NVDLA_CSC_wl.scala 808:97:@16518.4]
  wire  _T_4760; // @[NV_NVDLA_CSC_wl.scala 808:97:@16520.4]
  wire  _T_4762; // @[NV_NVDLA_CSC_wl.scala 808:97:@16522.4]
  wire  _T_4764; // @[NV_NVDLA_CSC_wl.scala 808:97:@16524.4]
  wire  _T_4766; // @[NV_NVDLA_CSC_wl.scala 808:97:@16526.4]
  wire  _T_4768; // @[NV_NVDLA_CSC_wl.scala 808:97:@16528.4]
  wire  _T_4770; // @[NV_NVDLA_CSC_wl.scala 808:97:@16530.4]
  wire  _T_4772; // @[NV_NVDLA_CSC_wl.scala 808:97:@16532.4]
  wire  _T_4774; // @[NV_NVDLA_CSC_wl.scala 808:97:@16534.4]
  wire  _T_4776; // @[NV_NVDLA_CSC_wl.scala 808:97:@16536.4]
  wire  _T_4778; // @[NV_NVDLA_CSC_wl.scala 808:97:@16538.4]
  wire  _T_4780; // @[NV_NVDLA_CSC_wl.scala 808:97:@16540.4]
  wire  _T_4782; // @[NV_NVDLA_CSC_wl.scala 808:97:@16542.4]
  wire  _T_4784; // @[NV_NVDLA_CSC_wl.scala 808:97:@16544.4]
  wire  _T_4786; // @[NV_NVDLA_CSC_wl.scala 808:97:@16546.4]
  wire  _T_4788; // @[NV_NVDLA_CSC_wl.scala 808:97:@16548.4]
  wire  _T_4790; // @[NV_NVDLA_CSC_wl.scala 808:97:@16550.4]
  wire  _T_4792; // @[NV_NVDLA_CSC_wl.scala 808:97:@16552.4]
  wire  _T_4794; // @[NV_NVDLA_CSC_wl.scala 808:97:@16554.4]
  wire  _T_4796; // @[NV_NVDLA_CSC_wl.scala 808:97:@16556.4]
  wire  _T_4798; // @[NV_NVDLA_CSC_wl.scala 808:97:@16558.4]
  wire  _T_4800; // @[NV_NVDLA_CSC_wl.scala 808:97:@16560.4]
  wire  _T_4802; // @[NV_NVDLA_CSC_wl.scala 808:97:@16562.4]
  wire  _T_4804; // @[NV_NVDLA_CSC_wl.scala 808:97:@16564.4]
  wire  _T_4806; // @[NV_NVDLA_CSC_wl.scala 808:97:@16566.4]
  wire  _T_4877; // @[NV_NVDLA_CSC_wl.scala 812:29:@16634.4]
  wire  _T_4878; // @[NV_NVDLA_CSC_wl.scala 814:96:@16700.6]
  wire  _T_4879; // @[NV_NVDLA_CSC_wl.scala 814:96:@16701.6]
  wire  _T_4880; // @[NV_NVDLA_CSC_wl.scala 814:96:@16702.6]
  wire  _T_4881; // @[NV_NVDLA_CSC_wl.scala 814:96:@16703.6]
  wire  _T_4882; // @[NV_NVDLA_CSC_wl.scala 814:96:@16704.6]
  wire  _T_4883; // @[NV_NVDLA_CSC_wl.scala 814:96:@16705.6]
  wire  _T_4884; // @[NV_NVDLA_CSC_wl.scala 814:96:@16706.6]
  wire  _T_4885; // @[NV_NVDLA_CSC_wl.scala 814:96:@16707.6]
  wire  _T_4886; // @[NV_NVDLA_CSC_wl.scala 814:96:@16708.6]
  wire  _T_4887; // @[NV_NVDLA_CSC_wl.scala 814:96:@16709.6]
  wire  _T_4888; // @[NV_NVDLA_CSC_wl.scala 814:96:@16710.6]
  wire  _T_4889; // @[NV_NVDLA_CSC_wl.scala 814:96:@16711.6]
  wire  _T_4890; // @[NV_NVDLA_CSC_wl.scala 814:96:@16712.6]
  wire  _T_4891; // @[NV_NVDLA_CSC_wl.scala 814:96:@16713.6]
  wire  _T_4892; // @[NV_NVDLA_CSC_wl.scala 814:96:@16714.6]
  wire  _T_4893; // @[NV_NVDLA_CSC_wl.scala 814:96:@16715.6]
  wire  _GEN_209; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_220; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_221; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_222; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_223; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_224; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_230; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_231; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_232; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_233; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_234; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_235; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_236; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_237; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_238; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_239; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_240; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_241; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_242; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_243; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_244; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_245; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_246; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_247; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_248; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_249; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_250; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_251; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_252; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_253; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_254; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_255; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_256; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_257; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_258; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_259; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_260; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_261; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_262; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_263; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_264; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_265; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_266; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_267; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_268; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_269; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_270; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_271; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_272; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_273; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_274; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_275; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_276; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_277; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_278; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_279; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_280; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_281; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_282; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_283; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  wire  _T_4916; // @[NV_NVDLA_CSC_wl.scala 816:29:@16750.4]
  wire  _T_4917; // @[NV_NVDLA_CSC_wl.scala 818:96:@16816.6]
  wire  _T_4918; // @[NV_NVDLA_CSC_wl.scala 818:96:@16817.6]
  wire  _T_4919; // @[NV_NVDLA_CSC_wl.scala 818:96:@16818.6]
  wire  _T_4920; // @[NV_NVDLA_CSC_wl.scala 818:96:@16819.6]
  wire  _T_4921; // @[NV_NVDLA_CSC_wl.scala 818:96:@16820.6]
  wire  _T_4922; // @[NV_NVDLA_CSC_wl.scala 818:96:@16821.6]
  wire  _T_4923; // @[NV_NVDLA_CSC_wl.scala 818:96:@16822.6]
  wire  _T_4924; // @[NV_NVDLA_CSC_wl.scala 818:96:@16823.6]
  wire  _T_4925; // @[NV_NVDLA_CSC_wl.scala 818:96:@16824.6]
  wire  _T_4926; // @[NV_NVDLA_CSC_wl.scala 818:96:@16825.6]
  wire  _T_4927; // @[NV_NVDLA_CSC_wl.scala 818:96:@16826.6]
  wire  _T_4928; // @[NV_NVDLA_CSC_wl.scala 818:96:@16827.6]
  wire  _T_4929; // @[NV_NVDLA_CSC_wl.scala 818:96:@16828.6]
  wire  _T_4930; // @[NV_NVDLA_CSC_wl.scala 818:96:@16829.6]
  wire  _T_4931; // @[NV_NVDLA_CSC_wl.scala 818:96:@16830.6]
  wire  _T_4932; // @[NV_NVDLA_CSC_wl.scala 818:96:@16831.6]
  wire  _GEN_289; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_348; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_349; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_350; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_351; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_352; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_353; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_354; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_355; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_356; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_357; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_358; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_359; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_360; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_361; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_362; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_363; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_364; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_365; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_366; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_367; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  wire  _GEN_368; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  NV_NVDLA_CSC_WL_dec NV_NVDLA_CSC_WL_dec ( // @[NV_NVDLA_CSC_wl.scala 778:23:@15836.4]
    .reset(NV_NVDLA_CSC_WL_dec_reset),
    .io_nvdla_core_clk(NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk),
    .io_input_valid(NV_NVDLA_CSC_WL_dec_io_input_valid),
    .io_input_bits_mask_0(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0),
    .io_input_bits_mask_1(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1),
    .io_input_bits_mask_2(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2),
    .io_input_bits_mask_3(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3),
    .io_input_bits_mask_4(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4),
    .io_input_bits_mask_5(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5),
    .io_input_bits_mask_6(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6),
    .io_input_bits_mask_7(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7),
    .io_input_bits_mask_8(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8),
    .io_input_bits_mask_9(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9),
    .io_input_bits_mask_10(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10),
    .io_input_bits_mask_11(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11),
    .io_input_bits_mask_12(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12),
    .io_input_bits_mask_13(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13),
    .io_input_bits_mask_14(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14),
    .io_input_bits_mask_15(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15),
    .io_input_bits_mask_16(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16),
    .io_input_bits_mask_17(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17),
    .io_input_bits_mask_18(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18),
    .io_input_bits_mask_19(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19),
    .io_input_bits_mask_20(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20),
    .io_input_bits_mask_21(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21),
    .io_input_bits_mask_22(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22),
    .io_input_bits_mask_23(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23),
    .io_input_bits_mask_24(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24),
    .io_input_bits_mask_25(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25),
    .io_input_bits_mask_26(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26),
    .io_input_bits_mask_27(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27),
    .io_input_bits_mask_28(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28),
    .io_input_bits_mask_29(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29),
    .io_input_bits_mask_30(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30),
    .io_input_bits_mask_31(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31),
    .io_input_bits_mask_32(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32),
    .io_input_bits_mask_33(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33),
    .io_input_bits_mask_34(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34),
    .io_input_bits_mask_35(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35),
    .io_input_bits_mask_36(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36),
    .io_input_bits_mask_37(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37),
    .io_input_bits_mask_38(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38),
    .io_input_bits_mask_39(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39),
    .io_input_bits_mask_40(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40),
    .io_input_bits_mask_41(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41),
    .io_input_bits_mask_42(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42),
    .io_input_bits_mask_43(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43),
    .io_input_bits_mask_44(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44),
    .io_input_bits_mask_45(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45),
    .io_input_bits_mask_46(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46),
    .io_input_bits_mask_47(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47),
    .io_input_bits_mask_48(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48),
    .io_input_bits_mask_49(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49),
    .io_input_bits_mask_50(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50),
    .io_input_bits_mask_51(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51),
    .io_input_bits_mask_52(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52),
    .io_input_bits_mask_53(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53),
    .io_input_bits_mask_54(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54),
    .io_input_bits_mask_55(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55),
    .io_input_bits_mask_56(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56),
    .io_input_bits_mask_57(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57),
    .io_input_bits_mask_58(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58),
    .io_input_bits_mask_59(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59),
    .io_input_bits_mask_60(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60),
    .io_input_bits_mask_61(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61),
    .io_input_bits_mask_62(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62),
    .io_input_bits_mask_63(NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63),
    .io_input_bits_data_0(NV_NVDLA_CSC_WL_dec_io_input_bits_data_0),
    .io_input_bits_data_1(NV_NVDLA_CSC_WL_dec_io_input_bits_data_1),
    .io_input_bits_data_2(NV_NVDLA_CSC_WL_dec_io_input_bits_data_2),
    .io_input_bits_data_3(NV_NVDLA_CSC_WL_dec_io_input_bits_data_3),
    .io_input_bits_data_4(NV_NVDLA_CSC_WL_dec_io_input_bits_data_4),
    .io_input_bits_data_5(NV_NVDLA_CSC_WL_dec_io_input_bits_data_5),
    .io_input_bits_data_6(NV_NVDLA_CSC_WL_dec_io_input_bits_data_6),
    .io_input_bits_data_7(NV_NVDLA_CSC_WL_dec_io_input_bits_data_7),
    .io_input_bits_data_8(NV_NVDLA_CSC_WL_dec_io_input_bits_data_8),
    .io_input_bits_data_9(NV_NVDLA_CSC_WL_dec_io_input_bits_data_9),
    .io_input_bits_data_10(NV_NVDLA_CSC_WL_dec_io_input_bits_data_10),
    .io_input_bits_data_11(NV_NVDLA_CSC_WL_dec_io_input_bits_data_11),
    .io_input_bits_data_12(NV_NVDLA_CSC_WL_dec_io_input_bits_data_12),
    .io_input_bits_data_13(NV_NVDLA_CSC_WL_dec_io_input_bits_data_13),
    .io_input_bits_data_14(NV_NVDLA_CSC_WL_dec_io_input_bits_data_14),
    .io_input_bits_data_15(NV_NVDLA_CSC_WL_dec_io_input_bits_data_15),
    .io_input_bits_data_16(NV_NVDLA_CSC_WL_dec_io_input_bits_data_16),
    .io_input_bits_data_17(NV_NVDLA_CSC_WL_dec_io_input_bits_data_17),
    .io_input_bits_data_18(NV_NVDLA_CSC_WL_dec_io_input_bits_data_18),
    .io_input_bits_data_19(NV_NVDLA_CSC_WL_dec_io_input_bits_data_19),
    .io_input_bits_data_20(NV_NVDLA_CSC_WL_dec_io_input_bits_data_20),
    .io_input_bits_data_21(NV_NVDLA_CSC_WL_dec_io_input_bits_data_21),
    .io_input_bits_data_22(NV_NVDLA_CSC_WL_dec_io_input_bits_data_22),
    .io_input_bits_data_23(NV_NVDLA_CSC_WL_dec_io_input_bits_data_23),
    .io_input_bits_data_24(NV_NVDLA_CSC_WL_dec_io_input_bits_data_24),
    .io_input_bits_data_25(NV_NVDLA_CSC_WL_dec_io_input_bits_data_25),
    .io_input_bits_data_26(NV_NVDLA_CSC_WL_dec_io_input_bits_data_26),
    .io_input_bits_data_27(NV_NVDLA_CSC_WL_dec_io_input_bits_data_27),
    .io_input_bits_data_28(NV_NVDLA_CSC_WL_dec_io_input_bits_data_28),
    .io_input_bits_data_29(NV_NVDLA_CSC_WL_dec_io_input_bits_data_29),
    .io_input_bits_data_30(NV_NVDLA_CSC_WL_dec_io_input_bits_data_30),
    .io_input_bits_data_31(NV_NVDLA_CSC_WL_dec_io_input_bits_data_31),
    .io_input_bits_data_32(NV_NVDLA_CSC_WL_dec_io_input_bits_data_32),
    .io_input_bits_data_33(NV_NVDLA_CSC_WL_dec_io_input_bits_data_33),
    .io_input_bits_data_34(NV_NVDLA_CSC_WL_dec_io_input_bits_data_34),
    .io_input_bits_data_35(NV_NVDLA_CSC_WL_dec_io_input_bits_data_35),
    .io_input_bits_data_36(NV_NVDLA_CSC_WL_dec_io_input_bits_data_36),
    .io_input_bits_data_37(NV_NVDLA_CSC_WL_dec_io_input_bits_data_37),
    .io_input_bits_data_38(NV_NVDLA_CSC_WL_dec_io_input_bits_data_38),
    .io_input_bits_data_39(NV_NVDLA_CSC_WL_dec_io_input_bits_data_39),
    .io_input_bits_data_40(NV_NVDLA_CSC_WL_dec_io_input_bits_data_40),
    .io_input_bits_data_41(NV_NVDLA_CSC_WL_dec_io_input_bits_data_41),
    .io_input_bits_data_42(NV_NVDLA_CSC_WL_dec_io_input_bits_data_42),
    .io_input_bits_data_43(NV_NVDLA_CSC_WL_dec_io_input_bits_data_43),
    .io_input_bits_data_44(NV_NVDLA_CSC_WL_dec_io_input_bits_data_44),
    .io_input_bits_data_45(NV_NVDLA_CSC_WL_dec_io_input_bits_data_45),
    .io_input_bits_data_46(NV_NVDLA_CSC_WL_dec_io_input_bits_data_46),
    .io_input_bits_data_47(NV_NVDLA_CSC_WL_dec_io_input_bits_data_47),
    .io_input_bits_data_48(NV_NVDLA_CSC_WL_dec_io_input_bits_data_48),
    .io_input_bits_data_49(NV_NVDLA_CSC_WL_dec_io_input_bits_data_49),
    .io_input_bits_data_50(NV_NVDLA_CSC_WL_dec_io_input_bits_data_50),
    .io_input_bits_data_51(NV_NVDLA_CSC_WL_dec_io_input_bits_data_51),
    .io_input_bits_data_52(NV_NVDLA_CSC_WL_dec_io_input_bits_data_52),
    .io_input_bits_data_53(NV_NVDLA_CSC_WL_dec_io_input_bits_data_53),
    .io_input_bits_data_54(NV_NVDLA_CSC_WL_dec_io_input_bits_data_54),
    .io_input_bits_data_55(NV_NVDLA_CSC_WL_dec_io_input_bits_data_55),
    .io_input_bits_data_56(NV_NVDLA_CSC_WL_dec_io_input_bits_data_56),
    .io_input_bits_data_57(NV_NVDLA_CSC_WL_dec_io_input_bits_data_57),
    .io_input_bits_data_58(NV_NVDLA_CSC_WL_dec_io_input_bits_data_58),
    .io_input_bits_data_59(NV_NVDLA_CSC_WL_dec_io_input_bits_data_59),
    .io_input_bits_data_60(NV_NVDLA_CSC_WL_dec_io_input_bits_data_60),
    .io_input_bits_data_61(NV_NVDLA_CSC_WL_dec_io_input_bits_data_61),
    .io_input_bits_data_62(NV_NVDLA_CSC_WL_dec_io_input_bits_data_62),
    .io_input_bits_data_63(NV_NVDLA_CSC_WL_dec_io_input_bits_data_63),
    .io_input_bits_sel_0(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0),
    .io_input_bits_sel_1(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1),
    .io_input_bits_sel_2(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2),
    .io_input_bits_sel_3(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3),
    .io_input_bits_sel_4(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4),
    .io_input_bits_sel_5(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5),
    .io_input_bits_sel_6(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6),
    .io_input_bits_sel_7(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7),
    .io_input_bits_sel_8(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8),
    .io_input_bits_sel_9(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9),
    .io_input_bits_sel_10(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10),
    .io_input_bits_sel_11(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11),
    .io_input_bits_sel_12(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12),
    .io_input_bits_sel_13(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13),
    .io_input_bits_sel_14(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14),
    .io_input_bits_sel_15(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15),
    .io_input_bits_sel_16(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16),
    .io_input_bits_sel_17(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17),
    .io_input_bits_sel_18(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18),
    .io_input_bits_sel_19(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19),
    .io_input_bits_sel_20(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20),
    .io_input_bits_sel_21(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21),
    .io_input_bits_sel_22(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22),
    .io_input_bits_sel_23(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23),
    .io_input_bits_sel_24(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24),
    .io_input_bits_sel_25(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25),
    .io_input_bits_sel_26(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26),
    .io_input_bits_sel_27(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27),
    .io_input_bits_sel_28(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28),
    .io_input_bits_sel_29(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29),
    .io_input_bits_sel_30(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30),
    .io_input_bits_sel_31(NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31),
    .io_input_mask_en(NV_NVDLA_CSC_WL_dec_io_input_mask_en),
    .io_output_valid(NV_NVDLA_CSC_WL_dec_io_output_valid),
    .io_output_bits_mask_0(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0),
    .io_output_bits_mask_1(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1),
    .io_output_bits_mask_2(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2),
    .io_output_bits_mask_3(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3),
    .io_output_bits_mask_4(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4),
    .io_output_bits_mask_5(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5),
    .io_output_bits_mask_6(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6),
    .io_output_bits_mask_7(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7),
    .io_output_bits_mask_8(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8),
    .io_output_bits_mask_9(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9),
    .io_output_bits_mask_10(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10),
    .io_output_bits_mask_11(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11),
    .io_output_bits_mask_12(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12),
    .io_output_bits_mask_13(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13),
    .io_output_bits_mask_14(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14),
    .io_output_bits_mask_15(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15),
    .io_output_bits_mask_16(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16),
    .io_output_bits_mask_17(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17),
    .io_output_bits_mask_18(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18),
    .io_output_bits_mask_19(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19),
    .io_output_bits_mask_20(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20),
    .io_output_bits_mask_21(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21),
    .io_output_bits_mask_22(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22),
    .io_output_bits_mask_23(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23),
    .io_output_bits_mask_24(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24),
    .io_output_bits_mask_25(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25),
    .io_output_bits_mask_26(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26),
    .io_output_bits_mask_27(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27),
    .io_output_bits_mask_28(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28),
    .io_output_bits_mask_29(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29),
    .io_output_bits_mask_30(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30),
    .io_output_bits_mask_31(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31),
    .io_output_bits_mask_32(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32),
    .io_output_bits_mask_33(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33),
    .io_output_bits_mask_34(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34),
    .io_output_bits_mask_35(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35),
    .io_output_bits_mask_36(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36),
    .io_output_bits_mask_37(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37),
    .io_output_bits_mask_38(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38),
    .io_output_bits_mask_39(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39),
    .io_output_bits_mask_40(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40),
    .io_output_bits_mask_41(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41),
    .io_output_bits_mask_42(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42),
    .io_output_bits_mask_43(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43),
    .io_output_bits_mask_44(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44),
    .io_output_bits_mask_45(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45),
    .io_output_bits_mask_46(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46),
    .io_output_bits_mask_47(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47),
    .io_output_bits_mask_48(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48),
    .io_output_bits_mask_49(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49),
    .io_output_bits_mask_50(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50),
    .io_output_bits_mask_51(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51),
    .io_output_bits_mask_52(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52),
    .io_output_bits_mask_53(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53),
    .io_output_bits_mask_54(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54),
    .io_output_bits_mask_55(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55),
    .io_output_bits_mask_56(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56),
    .io_output_bits_mask_57(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57),
    .io_output_bits_mask_58(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58),
    .io_output_bits_mask_59(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59),
    .io_output_bits_mask_60(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60),
    .io_output_bits_mask_61(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61),
    .io_output_bits_mask_62(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62),
    .io_output_bits_mask_63(NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63),
    .io_output_bits_data_0(NV_NVDLA_CSC_WL_dec_io_output_bits_data_0),
    .io_output_bits_data_1(NV_NVDLA_CSC_WL_dec_io_output_bits_data_1),
    .io_output_bits_data_2(NV_NVDLA_CSC_WL_dec_io_output_bits_data_2),
    .io_output_bits_data_3(NV_NVDLA_CSC_WL_dec_io_output_bits_data_3),
    .io_output_bits_data_4(NV_NVDLA_CSC_WL_dec_io_output_bits_data_4),
    .io_output_bits_data_5(NV_NVDLA_CSC_WL_dec_io_output_bits_data_5),
    .io_output_bits_data_6(NV_NVDLA_CSC_WL_dec_io_output_bits_data_6),
    .io_output_bits_data_7(NV_NVDLA_CSC_WL_dec_io_output_bits_data_7),
    .io_output_bits_data_8(NV_NVDLA_CSC_WL_dec_io_output_bits_data_8),
    .io_output_bits_data_9(NV_NVDLA_CSC_WL_dec_io_output_bits_data_9),
    .io_output_bits_data_10(NV_NVDLA_CSC_WL_dec_io_output_bits_data_10),
    .io_output_bits_data_11(NV_NVDLA_CSC_WL_dec_io_output_bits_data_11),
    .io_output_bits_data_12(NV_NVDLA_CSC_WL_dec_io_output_bits_data_12),
    .io_output_bits_data_13(NV_NVDLA_CSC_WL_dec_io_output_bits_data_13),
    .io_output_bits_data_14(NV_NVDLA_CSC_WL_dec_io_output_bits_data_14),
    .io_output_bits_data_15(NV_NVDLA_CSC_WL_dec_io_output_bits_data_15),
    .io_output_bits_data_16(NV_NVDLA_CSC_WL_dec_io_output_bits_data_16),
    .io_output_bits_data_17(NV_NVDLA_CSC_WL_dec_io_output_bits_data_17),
    .io_output_bits_data_18(NV_NVDLA_CSC_WL_dec_io_output_bits_data_18),
    .io_output_bits_data_19(NV_NVDLA_CSC_WL_dec_io_output_bits_data_19),
    .io_output_bits_data_20(NV_NVDLA_CSC_WL_dec_io_output_bits_data_20),
    .io_output_bits_data_21(NV_NVDLA_CSC_WL_dec_io_output_bits_data_21),
    .io_output_bits_data_22(NV_NVDLA_CSC_WL_dec_io_output_bits_data_22),
    .io_output_bits_data_23(NV_NVDLA_CSC_WL_dec_io_output_bits_data_23),
    .io_output_bits_data_24(NV_NVDLA_CSC_WL_dec_io_output_bits_data_24),
    .io_output_bits_data_25(NV_NVDLA_CSC_WL_dec_io_output_bits_data_25),
    .io_output_bits_data_26(NV_NVDLA_CSC_WL_dec_io_output_bits_data_26),
    .io_output_bits_data_27(NV_NVDLA_CSC_WL_dec_io_output_bits_data_27),
    .io_output_bits_data_28(NV_NVDLA_CSC_WL_dec_io_output_bits_data_28),
    .io_output_bits_data_29(NV_NVDLA_CSC_WL_dec_io_output_bits_data_29),
    .io_output_bits_data_30(NV_NVDLA_CSC_WL_dec_io_output_bits_data_30),
    .io_output_bits_data_31(NV_NVDLA_CSC_WL_dec_io_output_bits_data_31),
    .io_output_bits_data_32(NV_NVDLA_CSC_WL_dec_io_output_bits_data_32),
    .io_output_bits_data_33(NV_NVDLA_CSC_WL_dec_io_output_bits_data_33),
    .io_output_bits_data_34(NV_NVDLA_CSC_WL_dec_io_output_bits_data_34),
    .io_output_bits_data_35(NV_NVDLA_CSC_WL_dec_io_output_bits_data_35),
    .io_output_bits_data_36(NV_NVDLA_CSC_WL_dec_io_output_bits_data_36),
    .io_output_bits_data_37(NV_NVDLA_CSC_WL_dec_io_output_bits_data_37),
    .io_output_bits_data_38(NV_NVDLA_CSC_WL_dec_io_output_bits_data_38),
    .io_output_bits_data_39(NV_NVDLA_CSC_WL_dec_io_output_bits_data_39),
    .io_output_bits_data_40(NV_NVDLA_CSC_WL_dec_io_output_bits_data_40),
    .io_output_bits_data_41(NV_NVDLA_CSC_WL_dec_io_output_bits_data_41),
    .io_output_bits_data_42(NV_NVDLA_CSC_WL_dec_io_output_bits_data_42),
    .io_output_bits_data_43(NV_NVDLA_CSC_WL_dec_io_output_bits_data_43),
    .io_output_bits_data_44(NV_NVDLA_CSC_WL_dec_io_output_bits_data_44),
    .io_output_bits_data_45(NV_NVDLA_CSC_WL_dec_io_output_bits_data_45),
    .io_output_bits_data_46(NV_NVDLA_CSC_WL_dec_io_output_bits_data_46),
    .io_output_bits_data_47(NV_NVDLA_CSC_WL_dec_io_output_bits_data_47),
    .io_output_bits_data_48(NV_NVDLA_CSC_WL_dec_io_output_bits_data_48),
    .io_output_bits_data_49(NV_NVDLA_CSC_WL_dec_io_output_bits_data_49),
    .io_output_bits_data_50(NV_NVDLA_CSC_WL_dec_io_output_bits_data_50),
    .io_output_bits_data_51(NV_NVDLA_CSC_WL_dec_io_output_bits_data_51),
    .io_output_bits_data_52(NV_NVDLA_CSC_WL_dec_io_output_bits_data_52),
    .io_output_bits_data_53(NV_NVDLA_CSC_WL_dec_io_output_bits_data_53),
    .io_output_bits_data_54(NV_NVDLA_CSC_WL_dec_io_output_bits_data_54),
    .io_output_bits_data_55(NV_NVDLA_CSC_WL_dec_io_output_bits_data_55),
    .io_output_bits_data_56(NV_NVDLA_CSC_WL_dec_io_output_bits_data_56),
    .io_output_bits_data_57(NV_NVDLA_CSC_WL_dec_io_output_bits_data_57),
    .io_output_bits_data_58(NV_NVDLA_CSC_WL_dec_io_output_bits_data_58),
    .io_output_bits_data_59(NV_NVDLA_CSC_WL_dec_io_output_bits_data_59),
    .io_output_bits_data_60(NV_NVDLA_CSC_WL_dec_io_output_bits_data_60),
    .io_output_bits_data_61(NV_NVDLA_CSC_WL_dec_io_output_bits_data_61),
    .io_output_bits_data_62(NV_NVDLA_CSC_WL_dec_io_output_bits_data_62),
    .io_output_bits_data_63(NV_NVDLA_CSC_WL_dec_io_output_bits_data_63),
    .io_output_bits_sel_0(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0),
    .io_output_bits_sel_1(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1),
    .io_output_bits_sel_2(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2),
    .io_output_bits_sel_3(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3),
    .io_output_bits_sel_4(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4),
    .io_output_bits_sel_5(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5),
    .io_output_bits_sel_6(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6),
    .io_output_bits_sel_7(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7),
    .io_output_bits_sel_8(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8),
    .io_output_bits_sel_9(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9),
    .io_output_bits_sel_10(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10),
    .io_output_bits_sel_11(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11),
    .io_output_bits_sel_12(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12),
    .io_output_bits_sel_13(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13),
    .io_output_bits_sel_14(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14),
    .io_output_bits_sel_15(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15),
    .io_output_bits_sel_16(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16),
    .io_output_bits_sel_17(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17),
    .io_output_bits_sel_18(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18),
    .io_output_bits_sel_19(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19),
    .io_output_bits_sel_20(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20),
    .io_output_bits_sel_21(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21),
    .io_output_bits_sel_22(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22),
    .io_output_bits_sel_23(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23),
    .io_output_bits_sel_24(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24),
    .io_output_bits_sel_25(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25),
    .io_output_bits_sel_26(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26),
    .io_output_bits_sel_27(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27),
    .io_output_bits_sel_28(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28),
    .io_output_bits_sel_29(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29),
    .io_output_bits_sel_30(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30),
    .io_output_bits_sel_31(NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31)
  );
  assign _T_700 = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_wl.scala 97:35:@14287.4]
  assign _T_704 = io_sc_state == 2'h2; // @[NV_NVDLA_CSC_wl.scala 99:38:@14289.4]
  assign _T_706 = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_wl.scala 100:35:@14290.4]
  assign _T_707 = ~ _T_698; // @[NV_NVDLA_CSC_wl.scala 101:37:@14291.4]
  assign _T_708 = _T_704 & _T_707; // @[NV_NVDLA_CSC_wl.scala 101:35:@14292.4]
  assign _T_743 = io_reg2dp_op_en & _T_700; // @[NV_NVDLA_CSC_wl.scala 115:36:@14304.4]
  assign _T_749 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 120:42:@14308.6]
  assign _T_750 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 120:42:@14309.6]
  assign _T_752 = io_reg2dp_weight_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 121:46:@14311.6]
  assign _T_753 = io_reg2dp_weight_bank + 5'h1; // @[NV_NVDLA_CSC_wl.scala 121:46:@14312.6]
  assign _T_755 = 9'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_wl.scala 122:42:@14314.6]
  assign _T_756 = _T_755[5:3]; // @[NV_NVDLA_CSC_wl.scala 122:67:@14315.6]
  assign _GEN_0 = _T_743 ? _T_750 : _T_715; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  assign _GEN_1 = _T_743 ? _T_753 : _T_722; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  assign _GEN_2 = _T_743 ? _T_756 : _T_739; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  assign _GEN_3 = _T_743 ? io_reg2dp_weight_format : _T_742; // @[NV_NVDLA_CSC_wl.scala 119:19:@14307.4]
  assign _T_757 = _T_706 & io_reg2dp_skip_weight_rls; // @[NV_NVDLA_CSC_wl.scala 125:21:@14319.4]
  assign _T_758 = io_reg2dp_weight_bytes[20:6]; // @[NV_NVDLA_CSC_wl.scala 126:54:@14321.6]
  assign _T_759 = io_reg2dp_wmb_bytes[14:6]; // @[NV_NVDLA_CSC_wl.scala 127:70:@14323.6]
  assign _T_761 = _T_742 ? _T_759 : 9'h0; // @[NV_NVDLA_CSC_wl.scala 127:32:@14324.6]
  assign _GEN_4 = _T_757 ? _T_758 : _T_729; // @[NV_NVDLA_CSC_wl.scala 125:49:@14320.4]
  assign _GEN_5 = _T_757 ? _T_761 : _T_736; // @[NV_NVDLA_CSC_wl.scala 125:49:@14320.4]
  assign _T_1759 = _T_1712[35]; // @[NV_NVDLA_CSC_wl.scala 693:34:@15202.4]
  assign _T_857 = _T_1692 & _T_1759; // @[NV_NVDLA_CSC_wl.scala 203:36:@14402.4]
  assign _T_858 = io_sg2wl_reuse_rls | _T_857; // @[NV_NVDLA_CSC_wl.scala 207:25:@14403.4]
  assign _T_1755 = _T_1712[31:17]; // @[NV_NVDLA_CSC_wl.scala 689:44:@15197.4]
  assign _T_859 = io_sg2wl_reuse_rls ? _T_729 : _T_1755; // @[NV_NVDLA_CSC_wl.scala 208:29:@14405.4]
  assign _T_1754 = _T_1712[16:8]; // @[NV_NVDLA_CSC_wl.scala 688:45:@15195.4]
  assign _T_860 = io_sg2wl_reuse_rls ? _T_736 : _T_1754; // @[NV_NVDLA_CSC_wl.scala 209:30:@14407.4]
  assign _T_799 = _T_798 + _T_859; // @[NV_NVDLA_CSC_wl.scala 155:39:@14349.4]
  assign _T_800 = _T_798 + _T_859; // @[NV_NVDLA_CSC_wl.scala 155:39:@14350.4]
  assign _T_802 = {_T_722,9'h0}; // @[Cat.scala 30:58:@14351.4]
  assign _GEN_497 = {{1'd0}, _T_802}; // @[NV_NVDLA_CSC_wl.scala 156:48:@14352.4]
  assign _T_803 = _T_800 - _GEN_497; // @[NV_NVDLA_CSC_wl.scala 156:48:@14352.4]
  assign _T_804 = $unsigned(_T_803); // @[NV_NVDLA_CSC_wl.scala 156:48:@14353.4]
  assign _T_805 = _T_804[14:0]; // @[NV_NVDLA_CSC_wl.scala 156:48:@14354.4]
  assign _T_808 = _T_800 >= _GEN_497; // @[NV_NVDLA_CSC_wl.scala 157:48:@14356.4]
  assign _T_810 = ~ _T_858; // @[NV_NVDLA_CSC_wl.scala 158:88:@14357.4]
  assign _T_811 = _T_808 ? _T_805 : _T_800; // @[NV_NVDLA_CSC_wl.scala 158:113:@14358.4]
  assign _T_812 = _T_810 ? _T_798 : _T_811; // @[NV_NVDLA_CSC_wl.scala 158:87:@14359.4]
  assign _T_813 = io_sc2cdma_wt_pending_req ? 15'h0 : _T_812; // @[NV_NVDLA_CSC_wl.scala 158:28:@14360.4]
  assign _T_847 = io_sc2cdma_wt_pending_req | _T_858; // @[NV_NVDLA_CSC_wl.scala 184:21:@14388.4]
  assign _GEN_8 = _T_847 ? _T_813 : _T_798; // @[NV_NVDLA_CSC_wl.scala 184:30:@14389.4]
  assign _GEN_12 = _T_858 ? _T_859 : _T_867; // @[Reg.scala 20:19:@14414.4]
  assign _GEN_13 = _T_858 ? _T_860 : _T_871; // @[Reg.scala 20:19:@14420.4]
  assign _T_879 = io_sg2wl_pd_bits[0]; // @[NV_NVDLA_CSC_wl.scala 224:26:@14427.4 NV_NVDLA_CSC_wl.scala 228:19:@14430.4]
  assign _GEN_14 = io_sg2wl_pd_valid ? {{17'd0}, _T_879} : _T_882; // @[NV_NVDLA_CSC_wl.scala 232:30:@14432.4]
  assign _T_883 = _T_882[6:0]; // @[NV_NVDLA_CSC_wl.scala 241:31:@14435.4]
  assign _T_884 = _T_882[12:7]; // @[NV_NVDLA_CSC_wl.scala 242:31:@14436.4]
  assign _T_885 = _T_882[14:13]; // @[NV_NVDLA_CSC_wl.scala 243:29:@14437.4]
  assign _T_886 = _T_882[15]; // @[NV_NVDLA_CSC_wl.scala 244:31:@14438.4]
  assign _T_887 = _T_882[16]; // @[NV_NVDLA_CSC_wl.scala 245:29:@14439.4]
  assign _T_888 = _T_882[17]; // @[NV_NVDLA_CSC_wl.scala 246:30:@14440.4]
  assign _T_898 = _T_893 + 5'h1; // @[NV_NVDLA_CSC_wl.scala 257:37:@14444.4]
  assign _T_899 = _T_893 + 5'h1; // @[NV_NVDLA_CSC_wl.scala 257:37:@14445.4]
  assign _T_904 = _T_884[4:0]; // @[NV_NVDLA_CSC_wl.scala 259:39:@14448.4]
  assign _T_905 = _T_899 == _T_904; // @[NV_NVDLA_CSC_wl.scala 260:38:@14449.4]
  assign _T_902 = _T_905 ? 5'h0 : _T_899; // @[NV_NVDLA_CSC_wl.scala 258:59:@14446.4]
  assign _T_903 = _T_743 ? 5'h0 : _T_902; // @[NV_NVDLA_CSC_wl.scala 258:27:@14447.4]
  assign _T_908 = _T_893 != 5'h0; // @[NV_NVDLA_CSC_wl.scala 262:64:@14451.4]
  assign _T_909 = ~ _T_908; // @[NV_NVDLA_CSC_wl.scala 262:51:@14452.4]
  assign _T_911 = _T_909 ? 1'h0 : _T_896; // @[NV_NVDLA_CSC_wl.scala 262:50:@14453.4]
  assign _T_912 = _T_877 ? 1'h1 : _T_911; // @[NV_NVDLA_CSC_wl.scala 262:29:@14454.4]
  assign _T_913 = _T_743 | _T_912; // @[NV_NVDLA_CSC_wl.scala 263:38:@14455.4]
  assign _GEN_15 = _T_913 ? _T_903 : _T_893; // @[NV_NVDLA_CSC_wl.scala 265:28:@14456.4]
  assign _T_966 = _T_912 & _T_742; // @[NV_NVDLA_CSC_wl.scala 289:37:@14493.4]
  assign _T_964 = 2'h0 == _T_885; // @[Mux.scala 46:19:@14490.4]
  assign _T_942 = {1'h0,_T_883}; // @[Cat.scala 30:58:@14476.4]
  assign _T_962 = 2'h1 == _T_885; // @[Mux.scala 46:19:@14488.4]
  assign _T_951 = _T_942[6:0]; // @[NV_NVDLA_CSC_wl.scala 285:101:@14480.4]
  assign _T_954 = {1'h0,_T_951,1'h0}; // @[Cat.scala 30:58:@14482.4]
  assign _T_960 = 2'h2 == _T_885; // @[Mux.scala 46:19:@14486.4]
  assign _T_958 = {_T_951,1'h0}; // @[Cat.scala 30:58:@14484.4]
  assign _T_959 = _T_958 + _T_942; // @[NV_NVDLA_CSC_wl.scala 286:109:@14485.4]
  assign _T_944 = _T_942[5:0]; // @[NV_NVDLA_CSC_wl.scala 282:92:@14477.4]
  assign _T_947 = {1'h0,_T_944,2'h0}; // @[Cat.scala 30:58:@14479.4]
  assign _T_961 = _T_960 ? _T_959 : _T_947; // @[Mux.scala 46:16:@14487.4]
  assign _T_963 = _T_962 ? _T_954 : _T_961; // @[Mux.scala 46:16:@14489.4]
  assign _T_965 = _T_964 ? {{1'd0}, _T_942} : _T_963; // @[Mux.scala 46:16:@14491.4]
  assign _T_917 = _T_965[7:0]; // @[NV_NVDLA_CSC_wl.scala 271:31:@14460.4 NV_NVDLA_CSC_wl.scala 282:21:@14492.4]
  assign _T_968 = {3'h0,_T_917}; // @[Cat.scala 30:58:@14494.4]
  assign _T_969 = _T_920 < _T_968; // @[NV_NVDLA_CSC_wl.scala 289:75:@14495.4]
  assign _T_970 = _T_966 & _T_969; // @[NV_NVDLA_CSC_wl.scala 289:56:@14496.4]
  assign _T_924 = ~ _T_970; // @[NV_NVDLA_CSC_wl.scala 275:35:@14463.4]
  assign _T_927 = _T_924 ? 11'h0 : 11'h200; // @[NV_NVDLA_CSC_wl.scala 275:34:@14464.4]
  assign _T_929 = _T_912 ? _T_917 : 8'h0; // @[NV_NVDLA_CSC_wl.scala 276:34:@14465.4]
  assign _T_930 = _T_920 + _T_927; // @[NV_NVDLA_CSC_wl.scala 277:47:@14466.4]
  assign _T_931 = _T_920 + _T_927; // @[NV_NVDLA_CSC_wl.scala 277:47:@14467.4]
  assign _GEN_501 = {{3'd0}, _T_929}; // @[NV_NVDLA_CSC_wl.scala 277:69:@14468.4]
  assign _T_932 = _T_931 - _GEN_501; // @[NV_NVDLA_CSC_wl.scala 277:69:@14468.4]
  assign _T_933 = $unsigned(_T_932); // @[NV_NVDLA_CSC_wl.scala 277:69:@14469.4]
  assign _T_934 = _T_933[10:0]; // @[NV_NVDLA_CSC_wl.scala 277:69:@14470.4]
  assign _T_936 = ~ _T_887; // @[NV_NVDLA_CSC_wl.scala 278:82:@14471.4]
  assign _T_937 = _T_905 & _T_936; // @[NV_NVDLA_CSC_wl.scala 278:80:@14472.4]
  assign _T_938 = _T_937 & _T_886; // @[NV_NVDLA_CSC_wl.scala 278:96:@14473.4]
  assign _T_939 = _T_938 ? _T_923 : _T_934; // @[NV_NVDLA_CSC_wl.scala 278:65:@14474.4]
  assign _T_940 = _T_743 ? 11'h0 : _T_939; // @[NV_NVDLA_CSC_wl.scala 278:32:@14475.4]
  assign _T_972 = _T_743 | _T_966; // @[NV_NVDLA_CSC_wl.scala 290:43:@14499.4]
  assign _T_974 = _T_966 & _T_905; // @[NV_NVDLA_CSC_wl.scala 291:85:@14501.4]
  assign _T_975 = _T_974 & _T_887; // @[NV_NVDLA_CSC_wl.scala 291:101:@14502.4]
  assign _T_976 = _T_743 | _T_975; // @[NV_NVDLA_CSC_wl.scala 291:48:@14503.4]
  assign _GEN_16 = _T_972 ? _T_940 : _T_920; // @[NV_NVDLA_CSC_wl.scala 293:33:@14504.4]
  assign _GEN_17 = _T_976 ? _T_940 : _T_923; // @[NV_NVDLA_CSC_wl.scala 296:38:@14507.4]
  assign _T_1007 = _T_887 & _T_905; // @[NV_NVDLA_CSC_wl.scala 321:58:@14537.4]
  assign _T_1008 = _T_743 | _T_1007; // @[NV_NVDLA_CSC_wl.scala 321:42:@14538.4]
  assign _T_1010 = _T_886 & _T_905; // @[NV_NVDLA_CSC_wl.scala 322:48:@14539.4]
  assign _T_1012 = _T_1010 ? 1'h1 : _T_1003; // @[NV_NVDLA_CSC_wl.scala 322:32:@14540.4]
  assign _T_1013 = _T_1008 ? 1'h0 : _T_1012; // @[NV_NVDLA_CSC_wl.scala 321:32:@14541.4]
  assign _T_1015 = _T_1006 + 9'h1; // @[NV_NVDLA_CSC_wl.scala 323:39:@14542.4]
  assign _T_1016 = _T_1006 + 9'h1; // @[NV_NVDLA_CSC_wl.scala 323:39:@14543.4]
  assign _T_1018 = _T_905 & _T_887; // @[NV_NVDLA_CSC_wl.scala 325:43:@14544.4]
  assign _T_1020 = _T_1018 ? 9'h0 : _T_1016; // @[NV_NVDLA_CSC_wl.scala 325:28:@14545.4]
  assign _T_1021 = _T_743 ? 9'h0 : _T_1020; // @[NV_NVDLA_CSC_wl.scala 324:28:@14546.4]
  assign _T_1022 = _T_742 & _T_912; // @[NV_NVDLA_CSC_wl.scala 326:58:@14547.4]
  assign _T_1023 = _T_1022 & _T_905; // @[NV_NVDLA_CSC_wl.scala 326:75:@14548.4]
  assign _T_1024 = _T_1023 & _T_887; // @[NV_NVDLA_CSC_wl.scala 326:91:@14549.4]
  assign _T_1025 = _T_743 | _T_1024; // @[NV_NVDLA_CSC_wl.scala 326:39:@14550.4]
  assign _T_1026 = _T_742 & _T_970; // @[NV_NVDLA_CSC_wl.scala 326:126:@14551.4]
  assign _T_1027 = ~ _T_1003; // @[NV_NVDLA_CSC_wl.scala 326:144:@14552.4]
  assign _T_1028 = _T_1026 & _T_1027; // @[NV_NVDLA_CSC_wl.scala 326:142:@14553.4]
  assign _T_1029 = _T_1025 | _T_1028; // @[NV_NVDLA_CSC_wl.scala 326:107:@14554.4]
  assign _T_1031 = _T_1003 | _T_924; // @[NV_NVDLA_CSC_wl.scala 327:47:@14556.4]
  assign _T_1032 = _T_1031 ? _T_1006 : _T_1016; // @[NV_NVDLA_CSC_wl.scala 327:30:@14557.4]
  assign _GEN_20 = _T_1029 ? _T_1021 : _T_1006; // @[NV_NVDLA_CSC_wl.scala 330:29:@14559.4]
  assign _GEN_22 = _T_912 ? _T_883 : _T_1041; // @[NV_NVDLA_CSC_wl.scala 351:25:@14577.4]
  assign _GEN_23 = _T_912 ? _T_917 : _T_1044; // @[NV_NVDLA_CSC_wl.scala 351:25:@14577.4]
  assign _T_1063 = _T_912 & _T_888; // @[NV_NVDLA_CSC_wl.scala 355:25:@14581.4]
  assign _T_1064 = _T_1063 & _T_905; // @[NV_NVDLA_CSC_wl.scala 355:41:@14582.4]
  assign _GEN_24 = _T_1064 ? _T_1032 : _T_1047; // @[NV_NVDLA_CSC_wl.scala 355:57:@14583.4]
  assign _T_1067 = _T_888 & _T_905; // @[NV_NVDLA_CSC_wl.scala 362:41:@14592.6]
  assign _GEN_25 = _T_912 ? _T_905 : _T_1050; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  assign _GEN_26 = _T_912 ? _T_1010 : _T_1053; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  assign _GEN_27 = _T_912 ? _T_1007 : _T_1056; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  assign _GEN_28 = _T_912 ? _T_1067 : _T_1059; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  assign _GEN_29 = _T_912 ? _T_885 : _T_1062; // @[NV_NVDLA_CSC_wl.scala 358:25:@14586.4]
  assign _T_1076 = {_T_1062,1'h0,_T_1059,_T_1056,_T_1053,_T_1050,_T_1047,_T_1044,_T_1041}; // @[Cat.scala 30:58:@14603.4]
  assign _GEN_30 = _T_896 ? _T_1076 : _T_1101; // @[NV_NVDLA_CSC_wl.scala 394:37:@14621.4]
  assign _GEN_31 = _T_1081 ? _T_1101 : _T_1104; // @[NV_NVDLA_CSC_wl.scala 394:37:@14625.4]
  assign _GEN_32 = _T_1084 ? _T_1104 : _T_1107; // @[NV_NVDLA_CSC_wl.scala 394:37:@14629.4]
  assign _GEN_33 = _T_1087 ? _T_1107 : _T_1110; // @[NV_NVDLA_CSC_wl.scala 394:37:@14633.4]
  assign _GEN_34 = _T_1090 ? _T_1110 : _T_1113; // @[NV_NVDLA_CSC_wl.scala 394:37:@14637.4]
  assign _GEN_35 = _T_1093 ? _T_1113 : _T_1116; // @[NV_NVDLA_CSC_wl.scala 394:37:@14641.4]
  assign _T_1117 = _T_1116[6:0]; // @[NV_NVDLA_CSC_wl.scala 404:46:@14644.4]
  assign _T_1118 = _T_1116[14:7]; // @[NV_NVDLA_CSC_wl.scala 405:42:@14645.4]
  assign _T_1119 = _T_1116[23:15]; // @[NV_NVDLA_CSC_wl.scala 406:46:@14646.4]
  assign _T_1120 = _T_1116[24]; // @[NV_NVDLA_CSC_wl.scala 407:45:@14647.4]
  assign _T_1121 = _T_1116[25]; // @[NV_NVDLA_CSC_wl.scala 408:46:@14648.4]
  assign _T_1122 = _T_1116[26]; // @[NV_NVDLA_CSC_wl.scala 409:44:@14649.4]
  assign _T_1123 = _T_1116[27]; // @[NV_NVDLA_CSC_wl.scala 410:38:@14650.4]
  assign _T_1124 = _T_1116[30:29]; // @[NV_NVDLA_CSC_wl.scala 411:44:@14651.4]
  assign _T_1137 = ~ _T_1122; // @[NV_NVDLA_CSC_wl.scala 421:91:@14656.4]
  assign _T_1138 = _T_1121 & _T_1137; // @[NV_NVDLA_CSC_wl.scala 421:89:@14657.4]
  assign _T_1145 = _T_1096 & _T_1122; // @[NV_NVDLA_CSC_wl.scala 422:72:@14664.4]
  assign _T_1146 = _T_1145 & _T_742; // @[NV_NVDLA_CSC_wl.scala 422:92:@14665.4]
  assign _T_1147 = _T_743 | _T_1146; // @[NV_NVDLA_CSC_wl.scala 422:51:@14666.4]
  assign _T_1148 = _T_1096 & _T_742; // @[NV_NVDLA_CSC_wl.scala 424:40:@14667.4]
  assign _T_1149 = _T_743 | _T_1148; // @[NV_NVDLA_CSC_wl.scala 424:19:@14668.4]
  assign _T_1170 = _T_1163[63:0]; // @[NV_NVDLA_CSC_wl.scala 437:63:@14684.4]
  assign _T_1171 = {{127'd0}, _T_1170}; // @[NV_NVDLA_CSC_wl.scala 437:45:@14685.4]
  assign _T_1172 = ~ _T_742; // @[NV_NVDLA_CSC_wl.scala 437:108:@14686.4]
  assign _T_1176 = _T_1172 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12:@14688.4]
  assign _GEN_503 = {{127'd0}, _T_1176}; // @[NV_NVDLA_CSC_wl.scala 437:85:@14689.4]
  assign _T_1177 = _T_1171 | _GEN_503; // @[NV_NVDLA_CSC_wl.scala 437:85:@14689.4]
  assign _T_1183 = 319'hffffffffffffffff << _T_1118; // @[NV_NVDLA_CSC_wl.scala 438:56:@14691.4]
  assign _T_1184 = ~ _T_1183; // @[NV_NVDLA_CSC_wl.scala 438:25:@14692.4]
  assign _T_1185 = _T_1177[63:0]; // @[NV_NVDLA_CSC_wl.scala 439:41:@14693.4]
  assign _GEN_504 = {{255'd0}, _T_1185}; // @[NV_NVDLA_CSC_wl.scala 439:63:@14694.4]
  assign _T_1186 = _GEN_504 & _T_1184; // @[NV_NVDLA_CSC_wl.scala 439:63:@14694.4]
  assign _GEN_38 = _T_1096 ? _T_1186 : _T_1156; // @[NV_NVDLA_CSC_wl.scala 441:28:@14695.4]
  assign _T_1199 = _T_1163 >> _T_1118; // @[NV_NVDLA_CSC_wl.scala 450:49:@14705.4]
  assign _T_1208 = _T_1138 ? _T_1193 : _T_1199; // @[NV_NVDLA_CSC_wl.scala 453:84:@14710.4]
  assign _T_1209 = _T_743 ? 512'h0 : _T_1208; // @[NV_NVDLA_CSC_wl.scala 453:33:@14711.4]
  assign _T_1215 = _T_1117[4:0]; // @[NV_NVDLA_CSC_wl.scala 456:52:@14717.4]
  assign _T_1217 = {_T_1215,1'h0}; // @[Cat.scala 30:58:@14718.4]
  assign _GEN_506 = {{1'd0}, _T_1215}; // @[NV_NVDLA_CSC_wl.scala 456:69:@14720.4]
  assign _T_1219 = _T_1217 + _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@14720.4]
  assign _T_1220 = _T_1217 + _GEN_506; // @[NV_NVDLA_CSC_wl.scala 456:69:@14721.4]
  assign _GEN_39 = _T_1149 ? _T_1209 : _T_1163; // @[NV_NVDLA_CSC_wl.scala 458:34:@14722.4]
  assign _GEN_40 = _T_1147 ? _T_1209 : _T_1193; // @[NV_NVDLA_CSC_wl.scala 461:39:@14725.4]
  assign _GEN_41 = _T_1096 ? _T_1117 : _T_1226; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_42 = _T_1096 ? _T_1120 : _T_1229; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_43 = _T_1096 ? _T_1121 : _T_1232; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_44 = _T_1096 ? _T_1122 : _T_1235; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_45 = _T_1096 ? _T_1123 : _T_1238; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_46 = _T_1096 ? _T_1119 : _T_1241; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_47 = _T_1096 ? _T_1124 : _T_1244; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _GEN_48 = _T_1096 ? {{1'd0}, _T_1220} : _T_1247; // @[NV_NVDLA_CSC_wl.scala 477:28:@14738.4]
  assign _T_1318 = _T_1156[0]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14749.4]
  assign _T_1319 = _T_1156[1]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14751.4]
  assign _T_1320 = _T_1156[2]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14753.4]
  assign _T_1321 = _T_1156[3]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14755.4]
  assign _T_1322 = _T_1156[4]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14757.4]
  assign _T_1323 = _T_1156[5]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14759.4]
  assign _T_1324 = _T_1156[6]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14761.4]
  assign _T_1325 = _T_1156[7]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14763.4]
  assign _T_1326 = _T_1156[8]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14765.4]
  assign _T_1327 = _T_1156[9]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14767.4]
  assign _T_1328 = _T_1156[10]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14769.4]
  assign _T_1329 = _T_1156[11]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14771.4]
  assign _T_1330 = _T_1156[12]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14773.4]
  assign _T_1331 = _T_1156[13]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14775.4]
  assign _T_1332 = _T_1156[14]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14777.4]
  assign _T_1333 = _T_1156[15]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14779.4]
  assign _T_1334 = _T_1156[16]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14781.4]
  assign _T_1335 = _T_1156[17]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14783.4]
  assign _T_1336 = _T_1156[18]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14785.4]
  assign _T_1337 = _T_1156[19]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14787.4]
  assign _T_1338 = _T_1156[20]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14789.4]
  assign _T_1339 = _T_1156[21]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14791.4]
  assign _T_1340 = _T_1156[22]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14793.4]
  assign _T_1341 = _T_1156[23]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14795.4]
  assign _T_1342 = _T_1156[24]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14797.4]
  assign _T_1343 = _T_1156[25]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14799.4]
  assign _T_1344 = _T_1156[26]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14801.4]
  assign _T_1345 = _T_1156[27]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14803.4]
  assign _T_1346 = _T_1156[28]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14805.4]
  assign _T_1347 = _T_1156[29]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14807.4]
  assign _T_1348 = _T_1156[30]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14809.4]
  assign _T_1349 = _T_1156[31]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14811.4]
  assign _T_1350 = _T_1156[32]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14813.4]
  assign _T_1351 = _T_1156[33]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14815.4]
  assign _T_1352 = _T_1156[34]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14817.4]
  assign _T_1353 = _T_1156[35]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14819.4]
  assign _T_1354 = _T_1156[36]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14821.4]
  assign _T_1355 = _T_1156[37]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14823.4]
  assign _T_1356 = _T_1156[38]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14825.4]
  assign _T_1357 = _T_1156[39]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14827.4]
  assign _T_1358 = _T_1156[40]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14829.4]
  assign _T_1359 = _T_1156[41]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14831.4]
  assign _T_1360 = _T_1156[42]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14833.4]
  assign _T_1361 = _T_1156[43]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14835.4]
  assign _T_1362 = _T_1156[44]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14837.4]
  assign _T_1363 = _T_1156[45]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14839.4]
  assign _T_1364 = _T_1156[46]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14841.4]
  assign _T_1365 = _T_1156[47]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14843.4]
  assign _T_1366 = _T_1156[48]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14845.4]
  assign _T_1367 = _T_1156[49]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14847.4]
  assign _T_1368 = _T_1156[50]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14849.4]
  assign _T_1369 = _T_1156[51]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14851.4]
  assign _T_1370 = _T_1156[52]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14853.4]
  assign _T_1371 = _T_1156[53]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14855.4]
  assign _T_1372 = _T_1156[54]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14857.4]
  assign _T_1373 = _T_1156[55]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14859.4]
  assign _T_1374 = _T_1156[56]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14861.4]
  assign _T_1375 = _T_1156[57]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14863.4]
  assign _T_1376 = _T_1156[58]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14865.4]
  assign _T_1377 = _T_1156[59]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14867.4]
  assign _T_1378 = _T_1156[60]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14869.4]
  assign _T_1379 = _T_1156[61]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14871.4]
  assign _T_1380 = _T_1156[62]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14873.4]
  assign _T_1381 = _T_1156[63]; // @[NV_NVDLA_CSC_wl.scala 497:40:@14875.4]
  assign _T_1382 = _T_1318 + _T_1319; // @[NV_NVDLA_CSC_wl.scala 499:46:@14877.4]
  assign _GEN_507 = {{1'd0}, _T_1320}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14878.4]
  assign _T_1383 = _T_1382 + _GEN_507; // @[NV_NVDLA_CSC_wl.scala 499:46:@14878.4]
  assign _GEN_508 = {{2'd0}, _T_1321}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14879.4]
  assign _T_1384 = _T_1383 + _GEN_508; // @[NV_NVDLA_CSC_wl.scala 499:46:@14879.4]
  assign _GEN_509 = {{3'd0}, _T_1322}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14880.4]
  assign _T_1385 = _T_1384 + _GEN_509; // @[NV_NVDLA_CSC_wl.scala 499:46:@14880.4]
  assign _GEN_510 = {{4'd0}, _T_1323}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14881.4]
  assign _T_1386 = _T_1385 + _GEN_510; // @[NV_NVDLA_CSC_wl.scala 499:46:@14881.4]
  assign _GEN_511 = {{5'd0}, _T_1324}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14882.4]
  assign _T_1387 = _T_1386 + _GEN_511; // @[NV_NVDLA_CSC_wl.scala 499:46:@14882.4]
  assign _GEN_512 = {{6'd0}, _T_1325}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14883.4]
  assign _T_1388 = _T_1387 + _GEN_512; // @[NV_NVDLA_CSC_wl.scala 499:46:@14883.4]
  assign _GEN_513 = {{7'd0}, _T_1326}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14884.4]
  assign _T_1389 = _T_1388 + _GEN_513; // @[NV_NVDLA_CSC_wl.scala 499:46:@14884.4]
  assign _GEN_514 = {{8'd0}, _T_1327}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14885.4]
  assign _T_1390 = _T_1389 + _GEN_514; // @[NV_NVDLA_CSC_wl.scala 499:46:@14885.4]
  assign _GEN_515 = {{9'd0}, _T_1328}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14886.4]
  assign _T_1391 = _T_1390 + _GEN_515; // @[NV_NVDLA_CSC_wl.scala 499:46:@14886.4]
  assign _GEN_516 = {{10'd0}, _T_1329}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14887.4]
  assign _T_1392 = _T_1391 + _GEN_516; // @[NV_NVDLA_CSC_wl.scala 499:46:@14887.4]
  assign _GEN_517 = {{11'd0}, _T_1330}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14888.4]
  assign _T_1393 = _T_1392 + _GEN_517; // @[NV_NVDLA_CSC_wl.scala 499:46:@14888.4]
  assign _GEN_518 = {{12'd0}, _T_1331}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14889.4]
  assign _T_1394 = _T_1393 + _GEN_518; // @[NV_NVDLA_CSC_wl.scala 499:46:@14889.4]
  assign _GEN_519 = {{13'd0}, _T_1332}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14890.4]
  assign _T_1395 = _T_1394 + _GEN_519; // @[NV_NVDLA_CSC_wl.scala 499:46:@14890.4]
  assign _GEN_520 = {{14'd0}, _T_1333}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14891.4]
  assign _T_1396 = _T_1395 + _GEN_520; // @[NV_NVDLA_CSC_wl.scala 499:46:@14891.4]
  assign _GEN_521 = {{15'd0}, _T_1334}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14892.4]
  assign _T_1397 = _T_1396 + _GEN_521; // @[NV_NVDLA_CSC_wl.scala 499:46:@14892.4]
  assign _GEN_522 = {{16'd0}, _T_1335}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14893.4]
  assign _T_1398 = _T_1397 + _GEN_522; // @[NV_NVDLA_CSC_wl.scala 499:46:@14893.4]
  assign _GEN_523 = {{17'd0}, _T_1336}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14894.4]
  assign _T_1399 = _T_1398 + _GEN_523; // @[NV_NVDLA_CSC_wl.scala 499:46:@14894.4]
  assign _GEN_524 = {{18'd0}, _T_1337}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14895.4]
  assign _T_1400 = _T_1399 + _GEN_524; // @[NV_NVDLA_CSC_wl.scala 499:46:@14895.4]
  assign _GEN_525 = {{19'd0}, _T_1338}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14896.4]
  assign _T_1401 = _T_1400 + _GEN_525; // @[NV_NVDLA_CSC_wl.scala 499:46:@14896.4]
  assign _GEN_526 = {{20'd0}, _T_1339}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14897.4]
  assign _T_1402 = _T_1401 + _GEN_526; // @[NV_NVDLA_CSC_wl.scala 499:46:@14897.4]
  assign _GEN_527 = {{21'd0}, _T_1340}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14898.4]
  assign _T_1403 = _T_1402 + _GEN_527; // @[NV_NVDLA_CSC_wl.scala 499:46:@14898.4]
  assign _GEN_528 = {{22'd0}, _T_1341}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14899.4]
  assign _T_1404 = _T_1403 + _GEN_528; // @[NV_NVDLA_CSC_wl.scala 499:46:@14899.4]
  assign _GEN_529 = {{23'd0}, _T_1342}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14900.4]
  assign _T_1405 = _T_1404 + _GEN_529; // @[NV_NVDLA_CSC_wl.scala 499:46:@14900.4]
  assign _GEN_530 = {{24'd0}, _T_1343}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14901.4]
  assign _T_1406 = _T_1405 + _GEN_530; // @[NV_NVDLA_CSC_wl.scala 499:46:@14901.4]
  assign _GEN_531 = {{25'd0}, _T_1344}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14902.4]
  assign _T_1407 = _T_1406 + _GEN_531; // @[NV_NVDLA_CSC_wl.scala 499:46:@14902.4]
  assign _GEN_532 = {{26'd0}, _T_1345}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14903.4]
  assign _T_1408 = _T_1407 + _GEN_532; // @[NV_NVDLA_CSC_wl.scala 499:46:@14903.4]
  assign _GEN_533 = {{27'd0}, _T_1346}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14904.4]
  assign _T_1409 = _T_1408 + _GEN_533; // @[NV_NVDLA_CSC_wl.scala 499:46:@14904.4]
  assign _GEN_534 = {{28'd0}, _T_1347}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14905.4]
  assign _T_1410 = _T_1409 + _GEN_534; // @[NV_NVDLA_CSC_wl.scala 499:46:@14905.4]
  assign _GEN_535 = {{29'd0}, _T_1348}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14906.4]
  assign _T_1411 = _T_1410 + _GEN_535; // @[NV_NVDLA_CSC_wl.scala 499:46:@14906.4]
  assign _GEN_536 = {{30'd0}, _T_1349}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14907.4]
  assign _T_1412 = _T_1411 + _GEN_536; // @[NV_NVDLA_CSC_wl.scala 499:46:@14907.4]
  assign _GEN_537 = {{31'd0}, _T_1350}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14908.4]
  assign _T_1413 = _T_1412 + _GEN_537; // @[NV_NVDLA_CSC_wl.scala 499:46:@14908.4]
  assign _GEN_538 = {{32'd0}, _T_1351}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14909.4]
  assign _T_1414 = _T_1413 + _GEN_538; // @[NV_NVDLA_CSC_wl.scala 499:46:@14909.4]
  assign _GEN_539 = {{33'd0}, _T_1352}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14910.4]
  assign _T_1415 = _T_1414 + _GEN_539; // @[NV_NVDLA_CSC_wl.scala 499:46:@14910.4]
  assign _GEN_540 = {{34'd0}, _T_1353}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14911.4]
  assign _T_1416 = _T_1415 + _GEN_540; // @[NV_NVDLA_CSC_wl.scala 499:46:@14911.4]
  assign _GEN_541 = {{35'd0}, _T_1354}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14912.4]
  assign _T_1417 = _T_1416 + _GEN_541; // @[NV_NVDLA_CSC_wl.scala 499:46:@14912.4]
  assign _GEN_542 = {{36'd0}, _T_1355}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14913.4]
  assign _T_1418 = _T_1417 + _GEN_542; // @[NV_NVDLA_CSC_wl.scala 499:46:@14913.4]
  assign _GEN_543 = {{37'd0}, _T_1356}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14914.4]
  assign _T_1419 = _T_1418 + _GEN_543; // @[NV_NVDLA_CSC_wl.scala 499:46:@14914.4]
  assign _GEN_544 = {{38'd0}, _T_1357}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14915.4]
  assign _T_1420 = _T_1419 + _GEN_544; // @[NV_NVDLA_CSC_wl.scala 499:46:@14915.4]
  assign _GEN_545 = {{39'd0}, _T_1358}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14916.4]
  assign _T_1421 = _T_1420 + _GEN_545; // @[NV_NVDLA_CSC_wl.scala 499:46:@14916.4]
  assign _GEN_546 = {{40'd0}, _T_1359}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14917.4]
  assign _T_1422 = _T_1421 + _GEN_546; // @[NV_NVDLA_CSC_wl.scala 499:46:@14917.4]
  assign _GEN_547 = {{41'd0}, _T_1360}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14918.4]
  assign _T_1423 = _T_1422 + _GEN_547; // @[NV_NVDLA_CSC_wl.scala 499:46:@14918.4]
  assign _GEN_548 = {{42'd0}, _T_1361}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14919.4]
  assign _T_1424 = _T_1423 + _GEN_548; // @[NV_NVDLA_CSC_wl.scala 499:46:@14919.4]
  assign _GEN_549 = {{43'd0}, _T_1362}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14920.4]
  assign _T_1425 = _T_1424 + _GEN_549; // @[NV_NVDLA_CSC_wl.scala 499:46:@14920.4]
  assign _GEN_550 = {{44'd0}, _T_1363}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14921.4]
  assign _T_1426 = _T_1425 + _GEN_550; // @[NV_NVDLA_CSC_wl.scala 499:46:@14921.4]
  assign _GEN_551 = {{45'd0}, _T_1364}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14922.4]
  assign _T_1427 = _T_1426 + _GEN_551; // @[NV_NVDLA_CSC_wl.scala 499:46:@14922.4]
  assign _GEN_552 = {{46'd0}, _T_1365}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14923.4]
  assign _T_1428 = _T_1427 + _GEN_552; // @[NV_NVDLA_CSC_wl.scala 499:46:@14923.4]
  assign _GEN_553 = {{47'd0}, _T_1366}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14924.4]
  assign _T_1429 = _T_1428 + _GEN_553; // @[NV_NVDLA_CSC_wl.scala 499:46:@14924.4]
  assign _GEN_554 = {{48'd0}, _T_1367}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14925.4]
  assign _T_1430 = _T_1429 + _GEN_554; // @[NV_NVDLA_CSC_wl.scala 499:46:@14925.4]
  assign _GEN_555 = {{49'd0}, _T_1368}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14926.4]
  assign _T_1431 = _T_1430 + _GEN_555; // @[NV_NVDLA_CSC_wl.scala 499:46:@14926.4]
  assign _GEN_556 = {{50'd0}, _T_1369}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14927.4]
  assign _T_1432 = _T_1431 + _GEN_556; // @[NV_NVDLA_CSC_wl.scala 499:46:@14927.4]
  assign _GEN_557 = {{51'd0}, _T_1370}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14928.4]
  assign _T_1433 = _T_1432 + _GEN_557; // @[NV_NVDLA_CSC_wl.scala 499:46:@14928.4]
  assign _GEN_558 = {{52'd0}, _T_1371}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14929.4]
  assign _T_1434 = _T_1433 + _GEN_558; // @[NV_NVDLA_CSC_wl.scala 499:46:@14929.4]
  assign _GEN_559 = {{53'd0}, _T_1372}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14930.4]
  assign _T_1435 = _T_1434 + _GEN_559; // @[NV_NVDLA_CSC_wl.scala 499:46:@14930.4]
  assign _GEN_560 = {{54'd0}, _T_1373}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14931.4]
  assign _T_1436 = _T_1435 + _GEN_560; // @[NV_NVDLA_CSC_wl.scala 499:46:@14931.4]
  assign _GEN_561 = {{55'd0}, _T_1374}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14932.4]
  assign _T_1437 = _T_1436 + _GEN_561; // @[NV_NVDLA_CSC_wl.scala 499:46:@14932.4]
  assign _GEN_562 = {{56'd0}, _T_1375}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14933.4]
  assign _T_1438 = _T_1437 + _GEN_562; // @[NV_NVDLA_CSC_wl.scala 499:46:@14933.4]
  assign _GEN_563 = {{57'd0}, _T_1376}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14934.4]
  assign _T_1439 = _T_1438 + _GEN_563; // @[NV_NVDLA_CSC_wl.scala 499:46:@14934.4]
  assign _GEN_564 = {{58'd0}, _T_1377}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14935.4]
  assign _T_1440 = _T_1439 + _GEN_564; // @[NV_NVDLA_CSC_wl.scala 499:46:@14935.4]
  assign _GEN_565 = {{59'd0}, _T_1378}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14936.4]
  assign _T_1441 = _T_1440 + _GEN_565; // @[NV_NVDLA_CSC_wl.scala 499:46:@14936.4]
  assign _GEN_566 = {{60'd0}, _T_1379}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14937.4]
  assign _T_1442 = _T_1441 + _GEN_566; // @[NV_NVDLA_CSC_wl.scala 499:46:@14937.4]
  assign _GEN_567 = {{61'd0}, _T_1380}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14938.4]
  assign _T_1443 = _T_1442 + _GEN_567; // @[NV_NVDLA_CSC_wl.scala 499:46:@14938.4]
  assign _GEN_568 = {{62'd0}, _T_1381}; // @[NV_NVDLA_CSC_wl.scala 499:46:@14939.4]
  assign _T_1444 = _T_1443 + _GEN_568; // @[NV_NVDLA_CSC_wl.scala 499:46:@14939.4]
  assign _T_1453 = 191'hffffffffffffffff << _T_1226; // @[NV_NVDLA_CSC_wl.scala 505:57:@14942.4]
  assign _T_1454 = ~ _T_1453; // @[NV_NVDLA_CSC_wl.scala 505:26:@14943.4]
  assign _T_1456 = _T_1244 >= 2'h1; // @[NV_NVDLA_CSC_wl.scala 508:45:@14944.4]
  assign _T_1467 = _T_1456 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 508:27:@14947.4]
  assign _T_1469 = _T_1244 >= 2'h2; // @[NV_NVDLA_CSC_wl.scala 509:45:@14948.4]
  assign _T_1480 = _T_1469 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 509:27:@14951.4]
  assign _T_1482 = _T_1244 >= 2'h3; // @[NV_NVDLA_CSC_wl.scala 510:45:@14952.4]
  assign _T_1493 = _T_1482 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_wl.scala 510:27:@14955.4]
  assign _T_1494 = _T_1226[5:0]; // @[NV_NVDLA_CSC_wl.scala 514:50:@14956.4]
  assign _T_1496 = {_T_1494,1'h0}; // @[Cat.scala 30:58:@14957.4]
  assign _T_1497 = _T_1156[63:0]; // @[NV_NVDLA_CSC_wl.scala 515:39:@14958.4]
  assign _GEN_569 = {{127'd0}, _T_1497}; // @[NV_NVDLA_CSC_wl.scala 515:61:@14959.4]
  assign _T_1498 = _GEN_569 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 515:61:@14959.4]
  assign _T_1500 = _T_1497 >> _T_1226; // @[NV_NVDLA_CSC_wl.scala 516:62:@14961.4]
  assign _GEN_570 = {{127'd0}, _T_1500}; // @[NV_NVDLA_CSC_wl.scala 516:83:@14962.4]
  assign _T_1501 = _GEN_570 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 516:83:@14962.4]
  assign _GEN_571 = {{127'd0}, _T_1467}; // @[NV_NVDLA_CSC_wl.scala 516:100:@14963.4]
  assign _T_1502 = _T_1501 & _GEN_571; // @[NV_NVDLA_CSC_wl.scala 516:100:@14963.4]
  assign _T_1504 = _T_1497 >> _T_1496; // @[NV_NVDLA_CSC_wl.scala 517:62:@14965.4]
  assign _GEN_572 = {{127'd0}, _T_1504}; // @[NV_NVDLA_CSC_wl.scala 517:83:@14966.4]
  assign _T_1505 = _GEN_572 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 517:83:@14966.4]
  assign _GEN_573 = {{127'd0}, _T_1480}; // @[NV_NVDLA_CSC_wl.scala 517:100:@14967.4]
  assign _T_1506 = _T_1505 & _GEN_573; // @[NV_NVDLA_CSC_wl.scala 517:100:@14967.4]
  assign _T_1508 = _T_1497 >> _T_1247; // @[NV_NVDLA_CSC_wl.scala 518:62:@14969.4]
  assign _GEN_574 = {{127'd0}, _T_1508}; // @[NV_NVDLA_CSC_wl.scala 518:83:@14970.4]
  assign _T_1509 = _GEN_574 & _T_1454; // @[NV_NVDLA_CSC_wl.scala 518:83:@14970.4]
  assign _GEN_575 = {{127'd0}, _T_1493}; // @[NV_NVDLA_CSC_wl.scala 518:100:@14971.4]
  assign _T_1510 = _T_1509 & _GEN_575; // @[NV_NVDLA_CSC_wl.scala 518:100:@14971.4]
  assign _T_1517 = _T_739 == 3'h1; // @[NV_NVDLA_CSC_wl.scala 523:41:@14973.4]
  assign _T_1519 = _T_739 == 3'h2; // @[NV_NVDLA_CSC_wl.scala 524:41:@14974.4]
  assign _T_1520 = _T_1502[31:0]; // @[NV_NVDLA_CSC_wl.scala 524:82:@14975.4]
  assign _T_1521 = _T_1498[31:0]; // @[NV_NVDLA_CSC_wl.scala 524:122:@14976.4]
  assign _T_1522 = {_T_1520,_T_1521}; // @[Cat.scala 30:58:@14977.4]
  assign _T_1523 = _T_1510[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:44:@14978.4]
  assign _T_1524 = _T_1506[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:84:@14979.4]
  assign _T_1525 = _T_1502[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:124:@14980.4]
  assign _T_1526 = _T_1498[15:0]; // @[NV_NVDLA_CSC_wl.scala 525:164:@14981.4]
  assign _T_1529 = {_T_1523,_T_1524,_T_1525,_T_1526}; // @[Cat.scala 30:58:@14984.4]
  assign _T_1530 = _T_1519 ? _T_1522 : _T_1529; // @[NV_NVDLA_CSC_wl.scala 524:28:@14985.4]
  assign _T_1531 = _T_1517 ? _T_1498 : {{127'd0}, _T_1530}; // @[NV_NVDLA_CSC_wl.scala 523:28:@14986.4]
  assign _T_1532 = _T_743 ? 191'h0 : _T_1531; // @[NV_NVDLA_CSC_wl.scala 522:28:@14987.4]
  assign _GEN_576 = {{127'd0}, _T_1447}; // @[NV_NVDLA_CSC_wl.scala 528:61:@14988.4]
  assign _T_1533 = _T_1532 != _GEN_576; // @[NV_NVDLA_CSC_wl.scala 528:61:@14988.4]
  assign _T_1534 = _T_1223 & _T_1533; // @[NV_NVDLA_CSC_wl.scala 528:44:@14989.4]
  assign _GEN_577 = {{56'd0}, _T_1537}; // @[NV_NVDLA_CSC_wl.scala 534:57:@14992.4]
  assign _T_1541 = _GEN_577 < _T_1444; // @[NV_NVDLA_CSC_wl.scala 534:57:@14992.4]
  assign _T_1542 = _T_1223 & _T_1541; // @[NV_NVDLA_CSC_wl.scala 534:42:@14993.4]
  assign _T_1543 = ~ _T_1542; // @[NV_NVDLA_CSC_wl.scala 536:31:@14994.4]
  assign _T_1546 = _T_1543 ? 8'h0 : 8'h40; // @[NV_NVDLA_CSC_wl.scala 536:30:@14995.4]
  assign _T_1547 = _T_1537 + _T_1546; // @[NV_NVDLA_CSC_wl.scala 538:39:@14996.4]
  assign _T_1548 = _T_1537 + _T_1546; // @[NV_NVDLA_CSC_wl.scala 538:39:@14997.4]
  assign _GEN_578 = {{56'd0}, _T_1548}; // @[NV_NVDLA_CSC_wl.scala 538:57:@14998.4]
  assign _T_1549 = _GEN_578 - _T_1444; // @[NV_NVDLA_CSC_wl.scala 538:57:@14998.4]
  assign _T_1550 = $unsigned(_T_1549); // @[NV_NVDLA_CSC_wl.scala 538:57:@14999.4]
  assign _T_1551 = _T_1550[63:0]; // @[NV_NVDLA_CSC_wl.scala 538:57:@15000.4]
  assign _T_1553 = ~ _T_1235; // @[NV_NVDLA_CSC_wl.scala 540:29:@15001.4]
  assign _T_1554 = _T_1553 & _T_1232; // @[NV_NVDLA_CSC_wl.scala 540:47:@15002.4]
  assign _T_1555 = _T_1554 ? {{56'd0}, _T_1540} : _T_1551; // @[NV_NVDLA_CSC_wl.scala 540:28:@15003.4]
  assign _T_1556 = _T_743 ? 64'h0 : _T_1555; // @[NV_NVDLA_CSC_wl.scala 539:28:@15004.4]
  assign _T_1557 = _T_1223 & _T_1229; // @[NV_NVDLA_CSC_wl.scala 543:61:@15005.4]
  assign _T_1558 = _T_1557 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 543:81:@15006.4]
  assign _T_1559 = _T_743 | _T_1558; // @[NV_NVDLA_CSC_wl.scala 543:40:@15007.4]
  assign _T_1560 = _T_743 | _T_1223; // @[NV_NVDLA_CSC_wl.scala 545:19:@15008.4]
  assign _GEN_49 = _T_1560 ? _T_1556 : {{56'd0}, _T_1537}; // @[NV_NVDLA_CSC_wl.scala 545:39:@15009.4]
  assign _GEN_50 = _T_1559 ? _T_1556 : {{56'd0}, _T_1540}; // @[NV_NVDLA_CSC_wl.scala 548:30:@15012.4]
  assign _T_1568 = _T_1563 + 13'h1; // @[NV_NVDLA_CSC_wl.scala 556:39:@15017.4]
  assign _T_1569 = _T_1563 + 13'h1; // @[NV_NVDLA_CSC_wl.scala 556:39:@15018.4]
  assign _GEN_579 = {{1'd0}, _T_1569}; // @[NV_NVDLA_CSC_wl.scala 557:48:@15021.4]
  assign _T_1576 = _GEN_579 == _T_802; // @[NV_NVDLA_CSC_wl.scala 557:48:@15021.4]
  assign _T_1582 = _T_1576 ? 13'h0 : _T_1569; // @[NV_NVDLA_CSC_wl.scala 558:35:@15023.4]
  assign _T_1583 = _T_813[12:0]; // @[NV_NVDLA_CSC_wl.scala 560:53:@15024.4]
  assign _T_1586 = _T_1542 ? _T_1582 : _T_1563; // @[NV_NVDLA_CSC_wl.scala 562:28:@15027.4]
  assign _T_1587 = _T_1554 ? _T_1566 : _T_1586; // @[NV_NVDLA_CSC_wl.scala 561:28:@15028.4]
  assign _T_1588 = _T_708 ? _T_1583 : _T_1587; // @[NV_NVDLA_CSC_wl.scala 560:28:@15029.4]
  assign _T_1589 = _T_708 | _T_1542; // @[NV_NVDLA_CSC_wl.scala 566:40:@15030.4]
  assign _T_1590 = _T_1223 & _T_1232; // @[NV_NVDLA_CSC_wl.scala 566:76:@15031.4]
  assign _T_1591 = _T_1589 | _T_1590; // @[NV_NVDLA_CSC_wl.scala 566:55:@15032.4]
  assign _T_1592 = _T_1223 & _T_1223; // @[NV_NVDLA_CSC_wl.scala 567:66:@15033.4]
  assign _T_1593 = _T_1592 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 567:86:@15034.4]
  assign _T_1594 = _T_708 | _T_1593; // @[NV_NVDLA_CSC_wl.scala 567:45:@15035.4]
  assign _T_1600 = {_T_715,9'h0}; // @[Cat.scala 30:58:@15037.4]
  assign _GEN_580 = {{1'd0}, _T_1563}; // @[NV_NVDLA_CSC_wl.scala 568:39:@15038.4]
  assign _T_1601 = _GEN_580 + _T_1600; // @[NV_NVDLA_CSC_wl.scala 568:39:@15038.4]
  assign _T_1602 = _GEN_580 + _T_1600; // @[NV_NVDLA_CSC_wl.scala 568:39:@15039.4]
  assign _GEN_51 = _T_1591 ? _T_1588 : _T_1563; // @[NV_NVDLA_CSC_wl.scala 570:29:@15040.4]
  assign _GEN_52 = _T_1594 ? _T_1588 : _T_1566; // @[NV_NVDLA_CSC_wl.scala 573:34:@15043.4]
  assign _T_1609 = _T_743 | _T_1235; // @[NV_NVDLA_CSC_wl.scala 581:42:@15048.4]
  assign _T_1612 = _T_1232 ? 1'h1 : _T_1605; // @[NV_NVDLA_CSC_wl.scala 581:76:@15049.4]
  assign _T_1613 = _T_1609 ? 1'h0 : _T_1612; // @[NV_NVDLA_CSC_wl.scala 581:31:@15050.4]
  assign _T_1615 = _T_1608 + 15'h1; // @[NV_NVDLA_CSC_wl.scala 582:37:@15051.4]
  assign _T_1616 = _T_1608 + 15'h1; // @[NV_NVDLA_CSC_wl.scala 582:37:@15052.4]
  assign _T_1619 = _T_1235 ? 15'h0 : _T_1616; // @[NV_NVDLA_CSC_wl.scala 583:84:@15053.4]
  assign _T_1620 = _T_743 ? 15'h0 : _T_1619; // @[NV_NVDLA_CSC_wl.scala 583:27:@15054.4]
  assign _T_1621 = _T_1223 & _T_1235; // @[NV_NVDLA_CSC_wl.scala 584:59:@15055.4]
  assign _T_1622 = _T_743 | _T_1621; // @[NV_NVDLA_CSC_wl.scala 584:38:@15056.4]
  assign _T_1623 = ~ _T_1605; // @[NV_NVDLA_CSC_wl.scala 584:82:@15057.4]
  assign _T_1624 = _T_1623 & _T_1542; // @[NV_NVDLA_CSC_wl.scala 584:98:@15058.4]
  assign _T_1625 = _T_1622 | _T_1624; // @[NV_NVDLA_CSC_wl.scala 584:79:@15059.4]
  assign _T_1627 = _T_1605 | _T_1543; // @[NV_NVDLA_CSC_wl.scala 585:45:@15061.4]
  assign _T_1628 = _T_1627 ? _T_1608 : _T_1616; // @[NV_NVDLA_CSC_wl.scala 585:29:@15062.4]
  assign _GEN_53 = _T_1625 ? _T_1620 : _T_1608; // @[NV_NVDLA_CSC_wl.scala 588:28:@15064.4]
  assign _GEN_54 = _T_1542 ? _T_1602 : {{1'd0}, _T_1634}; // @[NV_NVDLA_CSC_wl.scala 609:23:@15079.4]
  assign _GEN_55 = _T_1223 ? _T_1229 : _T_1640; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  assign _GEN_56 = _T_1223 ? _T_1232 : _T_1643; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  assign _GEN_57 = _T_1223 ? _T_1235 : _T_1646; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  assign _GEN_58 = _T_1223 ? _T_1238 : _T_1649; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  assign _GEN_59 = _T_1223 ? _T_1444 : {{56'd0}, _T_1652}; // @[NV_NVDLA_CSC_wl.scala 613:28:@15083.4]
  assign _GEN_60 = _T_1560 ? _T_1532 : {{127'd0}, _T_1447}; // @[NV_NVDLA_CSC_wl.scala 621:39:@15091.4]
  assign _GEN_61 = _T_1223 ? _T_1241 : _T_1658; // @[NV_NVDLA_CSC_wl.scala 625:28:@15095.4]
  assign _T_1663 = _T_1223 & _T_1238; // @[NV_NVDLA_CSC_wl.scala 628:28:@15098.4]
  assign _GEN_62 = _T_1663 ? _T_1628 : _T_1661; // @[NV_NVDLA_CSC_wl.scala 628:41:@15099.4]
  assign _T_1672 = {_T_1649,_T_1646,_T_1643,_T_1640,_T_1661,_T_1658,_T_1652}; // @[Cat.scala 30:58:@15112.4]
  assign _GEN_63 = _T_1637 ? _T_1672 : _T_1697; // @[NV_NVDLA_CSC_wl.scala 669:36:@15146.4]
  assign _GEN_64 = _T_1655 ? _T_1447 : _T_1737; // @[NV_NVDLA_CSC_wl.scala 673:34:@15150.4]
  assign _GEN_65 = _T_1677 ? _T_1697 : _T_1700; // @[NV_NVDLA_CSC_wl.scala 669:36:@15154.4]
  assign _GEN_66 = _T_1717 ? _T_1737 : _T_1740; // @[NV_NVDLA_CSC_wl.scala 673:34:@15158.4]
  assign _GEN_67 = _T_1680 ? _T_1700 : _T_1703; // @[NV_NVDLA_CSC_wl.scala 669:36:@15162.4]
  assign _GEN_68 = _T_1720 ? _T_1740 : _T_1743; // @[NV_NVDLA_CSC_wl.scala 673:34:@15166.4]
  assign _GEN_69 = _T_1683 ? _T_1703 : _T_1706; // @[NV_NVDLA_CSC_wl.scala 669:36:@15170.4]
  assign _GEN_70 = _T_1723 ? _T_1743 : _T_1746; // @[NV_NVDLA_CSC_wl.scala 673:34:@15174.4]
  assign _GEN_71 = _T_1686 ? _T_1706 : _T_1709; // @[NV_NVDLA_CSC_wl.scala 669:36:@15178.4]
  assign _GEN_72 = _T_1726 ? _T_1746 : _T_1749; // @[NV_NVDLA_CSC_wl.scala 673:34:@15182.4]
  assign _GEN_73 = _T_1689 ? _T_1709 : _T_1712; // @[NV_NVDLA_CSC_wl.scala 669:36:@15186.4]
  assign _GEN_74 = _T_1729 ? _T_1749 : _T_1752; // @[NV_NVDLA_CSC_wl.scala 673:34:@15190.4]
  assign _T_1753 = _T_1712[7:0]; // @[NV_NVDLA_CSC_wl.scala 687:38:@15194.4]
  assign _T_1756 = _T_1712[32]; // @[NV_NVDLA_CSC_wl.scala 690:44:@15199.4]
  assign _T_1757 = _T_1712[33]; // @[NV_NVDLA_CSC_wl.scala 691:45:@15200.4]
  assign _T_1758 = _T_1712[34]; // @[NV_NVDLA_CSC_wl.scala 692:43:@15201.4]
  assign _T_1768 = io_sc2buf_wt_rd_data_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_wl.scala 702:37:@15206.4]
  assign _T_1770 = ~ _T_1758; // @[NV_NVDLA_CSC_wl.scala 704:55:@15207.4]
  assign _T_1771 = _T_1757 & _T_1770; // @[NV_NVDLA_CSC_wl.scala 704:53:@15208.4]
  assign _T_1773 = {2'h0,_T_1765}; // @[Cat.scala 30:58:@15209.4]
  assign _GEN_581 = {{1'd0}, _T_1762}; // @[NV_NVDLA_CSC_wl.scala 704:141:@15210.4]
  assign _T_1774 = _GEN_581 + _T_1768; // @[NV_NVDLA_CSC_wl.scala 704:141:@15210.4]
  assign _T_1775 = _GEN_581 + _T_1768; // @[NV_NVDLA_CSC_wl.scala 704:141:@15211.4]
  assign _T_1776 = _T_1775 - _T_1753; // @[NV_NVDLA_CSC_wl.scala 704:166:@15212.4]
  assign _T_1777 = $unsigned(_T_1776); // @[NV_NVDLA_CSC_wl.scala 704:166:@15213.4]
  assign _T_1778 = _T_1777[7:0]; // @[NV_NVDLA_CSC_wl.scala 704:166:@15214.4]
  assign _T_1779 = _T_1771 ? _T_1773 : {{1'd0}, _T_1778}; // @[NV_NVDLA_CSC_wl.scala 704:33:@15215.4]
  assign _T_1780 = _T_743 ? 9'h0 : _T_1779; // @[NV_NVDLA_CSC_wl.scala 703:35:@15216.4]
  assign _T_1781 = _T_1780[6:0]; // @[NV_NVDLA_CSC_wl.scala 704:182:@15217.4]
  assign _T_1782 = _T_743 | _T_1692; // @[NV_NVDLA_CSC_wl.scala 705:42:@15218.4]
  assign _T_1783 = _T_1692 & _T_1758; // @[NV_NVDLA_CSC_wl.scala 706:67:@15219.4]
  assign _T_1784 = _T_743 | _T_1783; // @[NV_NVDLA_CSC_wl.scala 706:47:@15220.4]
  assign _GEN_75 = _T_1782 ? _T_1781 : _T_1762; // @[NV_NVDLA_CSC_wl.scala 708:32:@15221.4]
  assign _GEN_76 = _T_1784 ? _T_1781 : _T_1765; // @[NV_NVDLA_CSC_wl.scala 711:37:@15224.4]
  assign _T_1790 = _T_1753 - _GEN_581; // @[NV_NVDLA_CSC_wl.scala 719:40:@15230.4]
  assign _T_1791 = $unsigned(_T_1790); // @[NV_NVDLA_CSC_wl.scala 719:40:@15231.4]
  assign _T_1792 = _T_1791[7:0]; // @[NV_NVDLA_CSC_wl.scala 719:40:@15232.4]
  assign _T_1795 = {_T_1792,3'h0}; // @[Cat.scala 30:58:@15234.4]
  assign _T_1796 = io_sc2buf_wt_rd_data_bits >> _T_1795; // @[NV_NVDLA_CSC_wl.scala 720:82:@15235.4]
  assign _T_1798 = _T_1762 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 721:58:@15236.4]
  assign _T_1799 = ~ _T_1798; // @[NV_NVDLA_CSC_wl.scala 721:38:@15237.4]
  assign _T_1801 = _T_1799 ? 512'h0 : _T_1786; // @[NV_NVDLA_CSC_wl.scala 721:36:@15238.4]
  assign _T_1803 = {_T_1753,3'h0}; // @[Cat.scala 30:58:@15239.4]
  assign _T_1804 = _T_1786 >> _T_1803; // @[NV_NVDLA_CSC_wl.scala 722:45:@15240.4]
  assign _T_1809 = _T_1765 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 725:98:@15243.4]
  assign _T_1810 = _T_1771 & _T_1809; // @[NV_NVDLA_CSC_wl.scala 725:71:@15244.4]
  assign _T_1811 = io_sc2buf_wt_rd_data_valid ? _T_1796 : _T_1804; // @[NV_NVDLA_CSC_wl.scala 726:31:@15245.4]
  assign _T_1812 = _T_1810 ? _T_1788 : _T_1811; // @[NV_NVDLA_CSC_wl.scala 725:31:@15246.4]
  assign _T_1813 = _T_743 ? 512'h0 : _T_1812; // @[NV_NVDLA_CSC_wl.scala 724:31:@15247.4]
  assign _T_1815 = _T_1781 != 7'h0; // @[NV_NVDLA_CSC_wl.scala 729:86:@15248.4]
  assign _T_1816 = _T_1692 & _T_1815; // @[NV_NVDLA_CSC_wl.scala 729:62:@15249.4]
  assign _T_1817 = _T_743 | _T_1816; // @[NV_NVDLA_CSC_wl.scala 729:42:@15250.4]
  assign _T_1821 = _T_1783 & _T_1815; // @[NV_NVDLA_CSC_wl.scala 730:86:@15253.4]
  assign _T_1822 = _T_743 | _T_1821; // @[NV_NVDLA_CSC_wl.scala 730:47:@15254.4]
  assign _T_1825 = {_T_1762,3'h0}; // @[Cat.scala 30:58:@15256.4]
  assign _GEN_583 = {{1023'd0}, io_sc2buf_wt_rd_data_bits}; // @[NV_NVDLA_CSC_wl.scala 731:55:@15257.4]
  assign _T_1826 = _GEN_583 << _T_1825; // @[NV_NVDLA_CSC_wl.scala 731:55:@15257.4]
  assign _T_1828 = io_sc2buf_wt_rd_data_valid ? _T_1826 : 1535'h0; // @[NV_NVDLA_CSC_wl.scala 732:32:@15258.4]
  assign _GEN_584 = {{1023'd0}, _T_1801}; // @[NV_NVDLA_CSC_wl.scala 744:42:@15331.4]
  assign _T_2292 = _T_1828 | _GEN_584; // @[NV_NVDLA_CSC_wl.scala 744:42:@15331.4]
  assign _T_2293 = _T_2292[7:0]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15333.6]
  assign _T_2294 = _T_2292[15:8]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15335.6]
  assign _T_2295 = _T_2292[23:16]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15337.6]
  assign _T_2296 = _T_2292[31:24]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15339.6]
  assign _T_2297 = _T_2292[39:32]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15341.6]
  assign _T_2298 = _T_2292[47:40]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15343.6]
  assign _T_2299 = _T_2292[55:48]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15345.6]
  assign _T_2300 = _T_2292[63:56]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15347.6]
  assign _T_2301 = _T_2292[71:64]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15349.6]
  assign _T_2302 = _T_2292[79:72]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15351.6]
  assign _T_2303 = _T_2292[87:80]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15353.6]
  assign _T_2304 = _T_2292[95:88]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15355.6]
  assign _T_2305 = _T_2292[103:96]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15357.6]
  assign _T_2306 = _T_2292[111:104]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15359.6]
  assign _T_2307 = _T_2292[119:112]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15361.6]
  assign _T_2308 = _T_2292[127:120]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15363.6]
  assign _T_2309 = _T_2292[135:128]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15365.6]
  assign _T_2310 = _T_2292[143:136]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15367.6]
  assign _T_2311 = _T_2292[151:144]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15369.6]
  assign _T_2312 = _T_2292[159:152]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15371.6]
  assign _T_2313 = _T_2292[167:160]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15373.6]
  assign _T_2314 = _T_2292[175:168]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15375.6]
  assign _T_2315 = _T_2292[183:176]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15377.6]
  assign _T_2316 = _T_2292[191:184]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15379.6]
  assign _T_2317 = _T_2292[199:192]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15381.6]
  assign _T_2318 = _T_2292[207:200]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15383.6]
  assign _T_2319 = _T_2292[215:208]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15385.6]
  assign _T_2320 = _T_2292[223:216]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15387.6]
  assign _T_2321 = _T_2292[231:224]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15389.6]
  assign _T_2322 = _T_2292[239:232]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15391.6]
  assign _T_2323 = _T_2292[247:240]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15393.6]
  assign _T_2324 = _T_2292[255:248]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15395.6]
  assign _T_2325 = _T_2292[263:256]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15397.6]
  assign _T_2326 = _T_2292[271:264]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15399.6]
  assign _T_2327 = _T_2292[279:272]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15401.6]
  assign _T_2328 = _T_2292[287:280]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15403.6]
  assign _T_2329 = _T_2292[295:288]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15405.6]
  assign _T_2330 = _T_2292[303:296]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15407.6]
  assign _T_2331 = _T_2292[311:304]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15409.6]
  assign _T_2332 = _T_2292[319:312]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15411.6]
  assign _T_2333 = _T_2292[327:320]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15413.6]
  assign _T_2334 = _T_2292[335:328]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15415.6]
  assign _T_2335 = _T_2292[343:336]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15417.6]
  assign _T_2336 = _T_2292[351:344]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15419.6]
  assign _T_2337 = _T_2292[359:352]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15421.6]
  assign _T_2338 = _T_2292[367:360]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15423.6]
  assign _T_2339 = _T_2292[375:368]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15425.6]
  assign _T_2340 = _T_2292[383:376]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15427.6]
  assign _T_2341 = _T_2292[391:384]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15429.6]
  assign _T_2342 = _T_2292[399:392]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15431.6]
  assign _T_2343 = _T_2292[407:400]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15433.6]
  assign _T_2344 = _T_2292[415:408]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15435.6]
  assign _T_2345 = _T_2292[423:416]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15437.6]
  assign _T_2346 = _T_2292[431:424]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15439.6]
  assign _T_2347 = _T_2292[439:432]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15441.6]
  assign _T_2348 = _T_2292[447:440]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15443.6]
  assign _T_2349 = _T_2292[455:448]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15445.6]
  assign _T_2350 = _T_2292[463:456]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15447.6]
  assign _T_2351 = _T_2292[471:464]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15449.6]
  assign _T_2352 = _T_2292[479:472]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15451.6]
  assign _T_2353 = _T_2292[487:480]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15453.6]
  assign _T_2354 = _T_2292[495:488]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15455.6]
  assign _T_2355 = _T_2292[503:496]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15457.6]
  assign _T_2356 = _T_2292[511:504]; // @[NV_NVDLA_CSC_wl.scala 747:45:@15459.6]
  assign _GEN_79 = _T_1692 ? _T_2293 : _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_80 = _T_1692 ? _T_2294 : _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_81 = _T_1692 ? _T_2295 : _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_82 = _T_1692 ? _T_2296 : _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_83 = _T_1692 ? _T_2297 : _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_84 = _T_1692 ? _T_2298 : _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_85 = _T_1692 ? _T_2299 : _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_86 = _T_1692 ? _T_2300 : _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_87 = _T_1692 ? _T_2301 : _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_88 = _T_1692 ? _T_2302 : _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_89 = _T_1692 ? _T_2303 : _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_90 = _T_1692 ? _T_2304 : _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_91 = _T_1692 ? _T_2305 : _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_92 = _T_1692 ? _T_2306 : _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_93 = _T_1692 ? _T_2307 : _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_94 = _T_1692 ? _T_2308 : _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_95 = _T_1692 ? _T_2309 : _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_96 = _T_1692 ? _T_2310 : _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_97 = _T_1692 ? _T_2311 : _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_98 = _T_1692 ? _T_2312 : _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_99 = _T_1692 ? _T_2313 : _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_100 = _T_1692 ? _T_2314 : _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_101 = _T_1692 ? _T_2315 : _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_102 = _T_1692 ? _T_2316 : _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_103 = _T_1692 ? _T_2317 : _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_104 = _T_1692 ? _T_2318 : _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_105 = _T_1692 ? _T_2319 : _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_106 = _T_1692 ? _T_2320 : _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_107 = _T_1692 ? _T_2321 : _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_108 = _T_1692 ? _T_2322 : _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_109 = _T_1692 ? _T_2323 : _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_110 = _T_1692 ? _T_2324 : _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_111 = _T_1692 ? _T_2325 : _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_112 = _T_1692 ? _T_2326 : _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_113 = _T_1692 ? _T_2327 : _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_114 = _T_1692 ? _T_2328 : _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_115 = _T_1692 ? _T_2329 : _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_116 = _T_1692 ? _T_2330 : _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_117 = _T_1692 ? _T_2331 : _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_118 = _T_1692 ? _T_2332 : _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_119 = _T_1692 ? _T_2333 : _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_120 = _T_1692 ? _T_2334 : _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_121 = _T_1692 ? _T_2335 : _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_122 = _T_1692 ? _T_2336 : _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_123 = _T_1692 ? _T_2337 : _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_124 = _T_1692 ? _T_2338 : _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_125 = _T_1692 ? _T_2339 : _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_126 = _T_1692 ? _T_2340 : _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_127 = _T_1692 ? _T_2341 : _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_128 = _T_1692 ? _T_2342 : _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_129 = _T_1692 ? _T_2343 : _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_130 = _T_1692 ? _T_2344 : _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_131 = _T_1692 ? _T_2345 : _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_132 = _T_1692 ? _T_2346 : _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_133 = _T_1692 ? _T_2347 : _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_134 = _T_1692 ? _T_2348 : _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_135 = _T_1692 ? _T_2349 : _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_136 = _T_1692 ? _T_2350 : _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_137 = _T_1692 ? _T_2351 : _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_138 = _T_1692 ? _T_2352 : _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_139 = _T_1692 ? _T_2353 : _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_140 = _T_1692 ? _T_2354 : _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_141 = _T_1692 ? _T_2355 : _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _GEN_142 = _T_1692 ? _T_2356 : _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 745:27:@15332.4]
  assign _T_2364 = _T_2362[30:0]; // @[NV_NVDLA_CSC_wl.scala 757:41:@15464.4]
  assign _T_2365 = _T_2362[31]; // @[NV_NVDLA_CSC_wl.scala 757:77:@15465.4]
  assign _T_2366 = {_T_2364,_T_2365}; // @[Cat.scala 30:58:@15466.4]
  assign _T_2367 = _T_2359 ? 32'h1 : _T_2366; // @[NV_NVDLA_CSC_wl.scala 756:27:@15467.4]
  assign _GEN_143 = _T_1692 ? _T_1756 : _T_2359; // @[NV_NVDLA_CSC_wl.scala 759:27:@15468.4]
  assign _GEN_144 = _T_1692 ? _T_2367 : _T_2362; // @[NV_NVDLA_CSC_wl.scala 759:27:@15468.4]
  assign _T_2939 = _T_1752[0]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15639.6]
  assign _T_2940 = _T_1752[1]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15640.6]
  assign _T_2941 = _T_1752[2]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15641.6]
  assign _T_2942 = _T_1752[3]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15642.6]
  assign _T_2943 = _T_1752[4]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15643.6]
  assign _T_2944 = _T_1752[5]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15644.6]
  assign _T_2945 = _T_1752[6]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15645.6]
  assign _T_2946 = _T_1752[7]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15646.6]
  assign _T_2947 = _T_1752[8]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15647.6]
  assign _T_2948 = _T_1752[9]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15648.6]
  assign _T_2949 = _T_1752[10]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15649.6]
  assign _T_2950 = _T_1752[11]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15650.6]
  assign _T_2951 = _T_1752[12]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15651.6]
  assign _T_2952 = _T_1752[13]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15652.6]
  assign _T_2953 = _T_1752[14]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15653.6]
  assign _T_2954 = _T_1752[15]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15654.6]
  assign _T_2955 = _T_1752[16]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15655.6]
  assign _T_2956 = _T_1752[17]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15656.6]
  assign _T_2957 = _T_1752[18]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15657.6]
  assign _T_2958 = _T_1752[19]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15658.6]
  assign _T_2959 = _T_1752[20]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15659.6]
  assign _T_2960 = _T_1752[21]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15660.6]
  assign _T_2961 = _T_1752[22]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15661.6]
  assign _T_2962 = _T_1752[23]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15662.6]
  assign _T_2963 = _T_1752[24]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15663.6]
  assign _T_2964 = _T_1752[25]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15664.6]
  assign _T_2965 = _T_1752[26]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15665.6]
  assign _T_2966 = _T_1752[27]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15666.6]
  assign _T_2967 = _T_1752[28]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15667.6]
  assign _T_2968 = _T_1752[29]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15668.6]
  assign _T_2969 = _T_1752[30]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15669.6]
  assign _T_2970 = _T_1752[31]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15670.6]
  assign _T_2971 = _T_1752[32]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15671.6]
  assign _T_2972 = _T_1752[33]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15672.6]
  assign _T_2973 = _T_1752[34]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15673.6]
  assign _T_2974 = _T_1752[35]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15674.6]
  assign _T_2975 = _T_1752[36]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15675.6]
  assign _T_2976 = _T_1752[37]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15676.6]
  assign _T_2977 = _T_1752[38]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15677.6]
  assign _T_2978 = _T_1752[39]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15678.6]
  assign _T_2979 = _T_1752[40]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15679.6]
  assign _T_2980 = _T_1752[41]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15680.6]
  assign _T_2981 = _T_1752[42]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15681.6]
  assign _T_2982 = _T_1752[43]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15682.6]
  assign _T_2983 = _T_1752[44]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15683.6]
  assign _T_2984 = _T_1752[45]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15684.6]
  assign _T_2985 = _T_1752[46]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15685.6]
  assign _T_2986 = _T_1752[47]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15686.6]
  assign _T_2987 = _T_1752[48]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15687.6]
  assign _T_2988 = _T_1752[49]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15688.6]
  assign _T_2989 = _T_1752[50]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15689.6]
  assign _T_2990 = _T_1752[51]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15690.6]
  assign _T_2991 = _T_1752[52]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15691.6]
  assign _T_2992 = _T_1752[53]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15692.6]
  assign _T_2993 = _T_1752[54]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15693.6]
  assign _T_2994 = _T_1752[55]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15694.6]
  assign _T_2995 = _T_1752[56]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15695.6]
  assign _T_2996 = _T_1752[57]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15696.6]
  assign _T_2997 = _T_1752[58]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15697.6]
  assign _T_2998 = _T_1752[59]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15698.6]
  assign _T_2999 = _T_1752[60]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15699.6]
  assign _T_3000 = _T_1752[61]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15700.6]
  assign _T_3001 = _T_1752[62]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15701.6]
  assign _T_3002 = _T_1752[63]; // @[NV_NVDLA_CSC_wl.scala 773:86:@15702.6]
  assign _GEN_145 = _T_1732 ? _T_2939 : _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_146 = _T_1732 ? _T_2940 : _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_147 = _T_1732 ? _T_2941 : _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_148 = _T_1732 ? _T_2942 : _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_149 = _T_1732 ? _T_2943 : _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_150 = _T_1732 ? _T_2944 : _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_151 = _T_1732 ? _T_2945 : _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_152 = _T_1732 ? _T_2946 : _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_153 = _T_1732 ? _T_2947 : _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_154 = _T_1732 ? _T_2948 : _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_155 = _T_1732 ? _T_2949 : _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_156 = _T_1732 ? _T_2950 : _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_157 = _T_1732 ? _T_2951 : _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_158 = _T_1732 ? _T_2952 : _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_159 = _T_1732 ? _T_2953 : _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_160 = _T_1732 ? _T_2954 : _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_161 = _T_1732 ? _T_2955 : _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_162 = _T_1732 ? _T_2956 : _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_163 = _T_1732 ? _T_2957 : _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_164 = _T_1732 ? _T_2958 : _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_165 = _T_1732 ? _T_2959 : _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_166 = _T_1732 ? _T_2960 : _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_167 = _T_1732 ? _T_2961 : _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_168 = _T_1732 ? _T_2962 : _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_169 = _T_1732 ? _T_2963 : _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_170 = _T_1732 ? _T_2964 : _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_171 = _T_1732 ? _T_2965 : _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_172 = _T_1732 ? _T_2966 : _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_173 = _T_1732 ? _T_2967 : _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_174 = _T_1732 ? _T_2968 : _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_175 = _T_1732 ? _T_2969 : _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_176 = _T_1732 ? _T_2970 : _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_177 = _T_1732 ? _T_2971 : _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_178 = _T_1732 ? _T_2972 : _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_179 = _T_1732 ? _T_2973 : _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_180 = _T_1732 ? _T_2974 : _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_181 = _T_1732 ? _T_2975 : _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_182 = _T_1732 ? _T_2976 : _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_183 = _T_1732 ? _T_2977 : _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_184 = _T_1732 ? _T_2978 : _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_185 = _T_1732 ? _T_2979 : _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_186 = _T_1732 ? _T_2980 : _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_187 = _T_1732 ? _T_2981 : _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_188 = _T_1732 ? _T_2982 : _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_189 = _T_1732 ? _T_2983 : _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_190 = _T_1732 ? _T_2984 : _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_191 = _T_1732 ? _T_2985 : _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_192 = _T_1732 ? _T_2986 : _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_193 = _T_1732 ? _T_2987 : _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_194 = _T_1732 ? _T_2988 : _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_195 = _T_1732 ? _T_2989 : _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_196 = _T_1732 ? _T_2990 : _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_197 = _T_1732 ? _T_2991 : _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_198 = _T_1732 ? _T_2992 : _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_199 = _T_1732 ? _T_2993 : _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_200 = _T_1732 ? _T_2994 : _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_201 = _T_1732 ? _T_2995 : _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_202 = _T_1732 ? _T_2996 : _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_203 = _T_1732 ? _T_2997 : _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_204 = _T_1732 ? _T_2998 : _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_205 = _T_1732 ? _T_2999 : _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_206 = _T_1732 ? _T_3000 : _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_207 = _T_1732 ? _T_3001 : _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _GEN_208 = _T_1732 ? _T_3002 : _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 772:25:@15638.4]
  assign _T_3076 = _T_1732 ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12:@15834.4]
  assign _T_3077 = NV_NVDLA_CSC_WL_dec_io_output_valid; // @[Bitwise.scala 72:15:@16002.4]
  assign _T_3080 = _T_3077 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@16003.4]
  assign _T_3087 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_7,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_6,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_5,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_4,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_3,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_2,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_1,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_0}; // @[NV_NVDLA_CSC_wl.scala 794:92:@16010.4]
  assign _T_3095 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_15,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_14,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_13,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_12,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_11,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_10,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_9,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_8,_T_3087}; // @[NV_NVDLA_CSC_wl.scala 794:92:@16018.4]
  assign _T_3102 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_23,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_22,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_21,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_20,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_19,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_18,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_17,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_16}; // @[NV_NVDLA_CSC_wl.scala 794:92:@16025.4]
  assign _T_3111 = {NV_NVDLA_CSC_WL_dec_io_output_bits_sel_31,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_30,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_29,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_28,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_27,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_26,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_25,NV_NVDLA_CSC_WL_dec_io_output_bits_sel_24,_T_3102,_T_3095}; // @[NV_NVDLA_CSC_wl.scala 794:92:@16034.4]
  assign _T_3112 = _T_3111[15:0]; // @[NV_NVDLA_CSC_wl.scala 794:99:@16035.4]
  assign _T_3113 = _T_3080 & _T_3112; // @[NV_NVDLA_CSC_wl.scala 794:71:@16036.4]
  assign _T_3149 = _T_3111[31:16]; // @[NV_NVDLA_CSC_wl.scala 795:99:@16070.4]
  assign _T_3150 = _T_3080 & _T_3149; // @[NV_NVDLA_CSC_wl.scala 795:71:@16071.4]
  assign _T_3152 = _T_3113 != 16'h0; // @[NV_NVDLA_CSC_wl.scala 796:49:@16072.4]
  assign _T_3154 = _T_3150 != 16'h0; // @[NV_NVDLA_CSC_wl.scala 797:49:@16073.4]
  assign _T_4481 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_0; // @[NV_NVDLA_CSC_wl.scala 807:91:@16246.4]
  assign _T_4482 = _T_4481 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16247.4]
  assign _T_4483 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_1; // @[NV_NVDLA_CSC_wl.scala 807:91:@16248.4]
  assign _T_4484 = _T_4483 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16249.4]
  assign _T_4485 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_2; // @[NV_NVDLA_CSC_wl.scala 807:91:@16250.4]
  assign _T_4486 = _T_4485 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16251.4]
  assign _T_4487 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_3; // @[NV_NVDLA_CSC_wl.scala 807:91:@16252.4]
  assign _T_4488 = _T_4487 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16253.4]
  assign _T_4489 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_4; // @[NV_NVDLA_CSC_wl.scala 807:91:@16254.4]
  assign _T_4490 = _T_4489 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16255.4]
  assign _T_4491 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_5; // @[NV_NVDLA_CSC_wl.scala 807:91:@16256.4]
  assign _T_4492 = _T_4491 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16257.4]
  assign _T_4493 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_6; // @[NV_NVDLA_CSC_wl.scala 807:91:@16258.4]
  assign _T_4494 = _T_4493 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16259.4]
  assign _T_4495 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_7; // @[NV_NVDLA_CSC_wl.scala 807:91:@16260.4]
  assign _T_4496 = _T_4495 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16261.4]
  assign _T_4497 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_8; // @[NV_NVDLA_CSC_wl.scala 807:91:@16262.4]
  assign _T_4498 = _T_4497 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16263.4]
  assign _T_4499 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_9; // @[NV_NVDLA_CSC_wl.scala 807:91:@16264.4]
  assign _T_4500 = _T_4499 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16265.4]
  assign _T_4501 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_10; // @[NV_NVDLA_CSC_wl.scala 807:91:@16266.4]
  assign _T_4502 = _T_4501 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16267.4]
  assign _T_4503 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_11; // @[NV_NVDLA_CSC_wl.scala 807:91:@16268.4]
  assign _T_4504 = _T_4503 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16269.4]
  assign _T_4505 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_12; // @[NV_NVDLA_CSC_wl.scala 807:91:@16270.4]
  assign _T_4506 = _T_4505 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16271.4]
  assign _T_4507 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_13; // @[NV_NVDLA_CSC_wl.scala 807:91:@16272.4]
  assign _T_4508 = _T_4507 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16273.4]
  assign _T_4509 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_14; // @[NV_NVDLA_CSC_wl.scala 807:91:@16274.4]
  assign _T_4510 = _T_4509 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16275.4]
  assign _T_4511 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_15; // @[NV_NVDLA_CSC_wl.scala 807:91:@16276.4]
  assign _T_4512 = _T_4511 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16277.4]
  assign _T_4513 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_16; // @[NV_NVDLA_CSC_wl.scala 807:91:@16278.4]
  assign _T_4514 = _T_4513 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16279.4]
  assign _T_4515 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_17; // @[NV_NVDLA_CSC_wl.scala 807:91:@16280.4]
  assign _T_4516 = _T_4515 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16281.4]
  assign _T_4517 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_18; // @[NV_NVDLA_CSC_wl.scala 807:91:@16282.4]
  assign _T_4518 = _T_4517 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16283.4]
  assign _T_4519 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_19; // @[NV_NVDLA_CSC_wl.scala 807:91:@16284.4]
  assign _T_4520 = _T_4519 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16285.4]
  assign _T_4521 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_20; // @[NV_NVDLA_CSC_wl.scala 807:91:@16286.4]
  assign _T_4522 = _T_4521 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16287.4]
  assign _T_4523 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_21; // @[NV_NVDLA_CSC_wl.scala 807:91:@16288.4]
  assign _T_4524 = _T_4523 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16289.4]
  assign _T_4525 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_22; // @[NV_NVDLA_CSC_wl.scala 807:91:@16290.4]
  assign _T_4526 = _T_4525 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16291.4]
  assign _T_4527 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_23; // @[NV_NVDLA_CSC_wl.scala 807:91:@16292.4]
  assign _T_4528 = _T_4527 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16293.4]
  assign _T_4529 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_24; // @[NV_NVDLA_CSC_wl.scala 807:91:@16294.4]
  assign _T_4530 = _T_4529 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16295.4]
  assign _T_4531 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_25; // @[NV_NVDLA_CSC_wl.scala 807:91:@16296.4]
  assign _T_4532 = _T_4531 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16297.4]
  assign _T_4533 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_26; // @[NV_NVDLA_CSC_wl.scala 807:91:@16298.4]
  assign _T_4534 = _T_4533 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16299.4]
  assign _T_4535 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_27; // @[NV_NVDLA_CSC_wl.scala 807:91:@16300.4]
  assign _T_4536 = _T_4535 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16301.4]
  assign _T_4537 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_28; // @[NV_NVDLA_CSC_wl.scala 807:91:@16302.4]
  assign _T_4538 = _T_4537 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16303.4]
  assign _T_4539 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_29; // @[NV_NVDLA_CSC_wl.scala 807:91:@16304.4]
  assign _T_4540 = _T_4539 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16305.4]
  assign _T_4541 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_30; // @[NV_NVDLA_CSC_wl.scala 807:91:@16306.4]
  assign _T_4542 = _T_4541 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16307.4]
  assign _T_4543 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_31; // @[NV_NVDLA_CSC_wl.scala 807:91:@16308.4]
  assign _T_4544 = _T_4543 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16309.4]
  assign _T_4545 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_32; // @[NV_NVDLA_CSC_wl.scala 807:91:@16310.4]
  assign _T_4546 = _T_4545 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16311.4]
  assign _T_4547 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_33; // @[NV_NVDLA_CSC_wl.scala 807:91:@16312.4]
  assign _T_4548 = _T_4547 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16313.4]
  assign _T_4549 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_34; // @[NV_NVDLA_CSC_wl.scala 807:91:@16314.4]
  assign _T_4550 = _T_4549 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16315.4]
  assign _T_4551 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_35; // @[NV_NVDLA_CSC_wl.scala 807:91:@16316.4]
  assign _T_4552 = _T_4551 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16317.4]
  assign _T_4553 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_36; // @[NV_NVDLA_CSC_wl.scala 807:91:@16318.4]
  assign _T_4554 = _T_4553 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16319.4]
  assign _T_4555 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_37; // @[NV_NVDLA_CSC_wl.scala 807:91:@16320.4]
  assign _T_4556 = _T_4555 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16321.4]
  assign _T_4557 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_38; // @[NV_NVDLA_CSC_wl.scala 807:91:@16322.4]
  assign _T_4558 = _T_4557 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16323.4]
  assign _T_4559 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_39; // @[NV_NVDLA_CSC_wl.scala 807:91:@16324.4]
  assign _T_4560 = _T_4559 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16325.4]
  assign _T_4561 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_40; // @[NV_NVDLA_CSC_wl.scala 807:91:@16326.4]
  assign _T_4562 = _T_4561 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16327.4]
  assign _T_4563 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_41; // @[NV_NVDLA_CSC_wl.scala 807:91:@16328.4]
  assign _T_4564 = _T_4563 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16329.4]
  assign _T_4565 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_42; // @[NV_NVDLA_CSC_wl.scala 807:91:@16330.4]
  assign _T_4566 = _T_4565 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16331.4]
  assign _T_4567 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_43; // @[NV_NVDLA_CSC_wl.scala 807:91:@16332.4]
  assign _T_4568 = _T_4567 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16333.4]
  assign _T_4569 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_44; // @[NV_NVDLA_CSC_wl.scala 807:91:@16334.4]
  assign _T_4570 = _T_4569 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16335.4]
  assign _T_4571 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_45; // @[NV_NVDLA_CSC_wl.scala 807:91:@16336.4]
  assign _T_4572 = _T_4571 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16337.4]
  assign _T_4573 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_46; // @[NV_NVDLA_CSC_wl.scala 807:91:@16338.4]
  assign _T_4574 = _T_4573 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16339.4]
  assign _T_4575 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_47; // @[NV_NVDLA_CSC_wl.scala 807:91:@16340.4]
  assign _T_4576 = _T_4575 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16341.4]
  assign _T_4577 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_48; // @[NV_NVDLA_CSC_wl.scala 807:91:@16342.4]
  assign _T_4578 = _T_4577 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16343.4]
  assign _T_4579 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_49; // @[NV_NVDLA_CSC_wl.scala 807:91:@16344.4]
  assign _T_4580 = _T_4579 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16345.4]
  assign _T_4581 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_50; // @[NV_NVDLA_CSC_wl.scala 807:91:@16346.4]
  assign _T_4582 = _T_4581 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16347.4]
  assign _T_4583 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_51; // @[NV_NVDLA_CSC_wl.scala 807:91:@16348.4]
  assign _T_4584 = _T_4583 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16349.4]
  assign _T_4585 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_52; // @[NV_NVDLA_CSC_wl.scala 807:91:@16350.4]
  assign _T_4586 = _T_4585 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16351.4]
  assign _T_4587 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_53; // @[NV_NVDLA_CSC_wl.scala 807:91:@16352.4]
  assign _T_4588 = _T_4587 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16353.4]
  assign _T_4589 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_54; // @[NV_NVDLA_CSC_wl.scala 807:91:@16354.4]
  assign _T_4590 = _T_4589 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16355.4]
  assign _T_4591 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_55; // @[NV_NVDLA_CSC_wl.scala 807:91:@16356.4]
  assign _T_4592 = _T_4591 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16357.4]
  assign _T_4593 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_56; // @[NV_NVDLA_CSC_wl.scala 807:91:@16358.4]
  assign _T_4594 = _T_4593 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16359.4]
  assign _T_4595 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_57; // @[NV_NVDLA_CSC_wl.scala 807:91:@16360.4]
  assign _T_4596 = _T_4595 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16361.4]
  assign _T_4597 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_58; // @[NV_NVDLA_CSC_wl.scala 807:91:@16362.4]
  assign _T_4598 = _T_4597 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16363.4]
  assign _T_4599 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_59; // @[NV_NVDLA_CSC_wl.scala 807:91:@16364.4]
  assign _T_4600 = _T_4599 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16365.4]
  assign _T_4601 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_60; // @[NV_NVDLA_CSC_wl.scala 807:91:@16366.4]
  assign _T_4602 = _T_4601 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16367.4]
  assign _T_4603 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_61; // @[NV_NVDLA_CSC_wl.scala 807:91:@16368.4]
  assign _T_4604 = _T_4603 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16369.4]
  assign _T_4605 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_62; // @[NV_NVDLA_CSC_wl.scala 807:91:@16370.4]
  assign _T_4606 = _T_4605 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16371.4]
  assign _T_4607 = NV_NVDLA_CSC_WL_dec_io_output_bits_mask_63; // @[NV_NVDLA_CSC_wl.scala 807:91:@16372.4]
  assign _T_4608 = _T_4607 & _T_3152; // @[NV_NVDLA_CSC_wl.scala 807:97:@16373.4]
  assign _T_4680 = _T_4481 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16440.4]
  assign _T_4682 = _T_4483 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16442.4]
  assign _T_4684 = _T_4485 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16444.4]
  assign _T_4686 = _T_4487 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16446.4]
  assign _T_4688 = _T_4489 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16448.4]
  assign _T_4690 = _T_4491 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16450.4]
  assign _T_4692 = _T_4493 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16452.4]
  assign _T_4694 = _T_4495 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16454.4]
  assign _T_4696 = _T_4497 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16456.4]
  assign _T_4698 = _T_4499 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16458.4]
  assign _T_4700 = _T_4501 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16460.4]
  assign _T_4702 = _T_4503 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16462.4]
  assign _T_4704 = _T_4505 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16464.4]
  assign _T_4706 = _T_4507 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16466.4]
  assign _T_4708 = _T_4509 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16468.4]
  assign _T_4710 = _T_4511 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16470.4]
  assign _T_4712 = _T_4513 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16472.4]
  assign _T_4714 = _T_4515 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16474.4]
  assign _T_4716 = _T_4517 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16476.4]
  assign _T_4718 = _T_4519 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16478.4]
  assign _T_4720 = _T_4521 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16480.4]
  assign _T_4722 = _T_4523 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16482.4]
  assign _T_4724 = _T_4525 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16484.4]
  assign _T_4726 = _T_4527 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16486.4]
  assign _T_4728 = _T_4529 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16488.4]
  assign _T_4730 = _T_4531 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16490.4]
  assign _T_4732 = _T_4533 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16492.4]
  assign _T_4734 = _T_4535 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16494.4]
  assign _T_4736 = _T_4537 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16496.4]
  assign _T_4738 = _T_4539 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16498.4]
  assign _T_4740 = _T_4541 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16500.4]
  assign _T_4742 = _T_4543 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16502.4]
  assign _T_4744 = _T_4545 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16504.4]
  assign _T_4746 = _T_4547 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16506.4]
  assign _T_4748 = _T_4549 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16508.4]
  assign _T_4750 = _T_4551 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16510.4]
  assign _T_4752 = _T_4553 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16512.4]
  assign _T_4754 = _T_4555 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16514.4]
  assign _T_4756 = _T_4557 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16516.4]
  assign _T_4758 = _T_4559 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16518.4]
  assign _T_4760 = _T_4561 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16520.4]
  assign _T_4762 = _T_4563 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16522.4]
  assign _T_4764 = _T_4565 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16524.4]
  assign _T_4766 = _T_4567 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16526.4]
  assign _T_4768 = _T_4569 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16528.4]
  assign _T_4770 = _T_4571 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16530.4]
  assign _T_4772 = _T_4573 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16532.4]
  assign _T_4774 = _T_4575 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16534.4]
  assign _T_4776 = _T_4577 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16536.4]
  assign _T_4778 = _T_4579 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16538.4]
  assign _T_4780 = _T_4581 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16540.4]
  assign _T_4782 = _T_4583 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16542.4]
  assign _T_4784 = _T_4585 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16544.4]
  assign _T_4786 = _T_4587 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16546.4]
  assign _T_4788 = _T_4589 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16548.4]
  assign _T_4790 = _T_4591 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16550.4]
  assign _T_4792 = _T_4593 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16552.4]
  assign _T_4794 = _T_4595 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16554.4]
  assign _T_4796 = _T_4597 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16556.4]
  assign _T_4798 = _T_4599 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16558.4]
  assign _T_4800 = _T_4601 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16560.4]
  assign _T_4802 = _T_4603 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16562.4]
  assign _T_4804 = _T_4605 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16564.4]
  assign _T_4806 = _T_4607 & _T_3154; // @[NV_NVDLA_CSC_wl.scala 808:97:@16566.4]
  assign _T_4877 = _T_3152 | _T_3157; // @[NV_NVDLA_CSC_wl.scala 812:29:@16634.4]
  assign _T_4878 = _T_3113[0]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16700.6]
  assign _T_4879 = _T_3113[1]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16701.6]
  assign _T_4880 = _T_3113[2]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16702.6]
  assign _T_4881 = _T_3113[3]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16703.6]
  assign _T_4882 = _T_3113[4]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16704.6]
  assign _T_4883 = _T_3113[5]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16705.6]
  assign _T_4884 = _T_3113[6]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16706.6]
  assign _T_4885 = _T_3113[7]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16707.6]
  assign _T_4886 = _T_3113[8]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16708.6]
  assign _T_4887 = _T_3113[9]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16709.6]
  assign _T_4888 = _T_3113[10]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16710.6]
  assign _T_4889 = _T_3113[11]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16711.6]
  assign _T_4890 = _T_3113[12]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16712.6]
  assign _T_4891 = _T_3113[13]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16713.6]
  assign _T_4892 = _T_3113[14]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16714.6]
  assign _T_4893 = _T_3113[15]; // @[NV_NVDLA_CSC_wl.scala 814:96:@16715.6]
  assign _GEN_209 = _T_4877 ? _T_4482 : _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_210 = _T_4877 ? _T_4484 : _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_211 = _T_4877 ? _T_4486 : _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_212 = _T_4877 ? _T_4488 : _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_213 = _T_4877 ? _T_4490 : _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_214 = _T_4877 ? _T_4492 : _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_215 = _T_4877 ? _T_4494 : _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_216 = _T_4877 ? _T_4496 : _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_217 = _T_4877 ? _T_4498 : _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_218 = _T_4877 ? _T_4500 : _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_219 = _T_4877 ? _T_4502 : _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_220 = _T_4877 ? _T_4504 : _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_221 = _T_4877 ? _T_4506 : _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_222 = _T_4877 ? _T_4508 : _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_223 = _T_4877 ? _T_4510 : _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_224 = _T_4877 ? _T_4512 : _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_225 = _T_4877 ? _T_4514 : _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_226 = _T_4877 ? _T_4516 : _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_227 = _T_4877 ? _T_4518 : _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_228 = _T_4877 ? _T_4520 : _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_229 = _T_4877 ? _T_4522 : _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_230 = _T_4877 ? _T_4524 : _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_231 = _T_4877 ? _T_4526 : _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_232 = _T_4877 ? _T_4528 : _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_233 = _T_4877 ? _T_4530 : _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_234 = _T_4877 ? _T_4532 : _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_235 = _T_4877 ? _T_4534 : _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_236 = _T_4877 ? _T_4536 : _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_237 = _T_4877 ? _T_4538 : _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_238 = _T_4877 ? _T_4540 : _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_239 = _T_4877 ? _T_4542 : _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_240 = _T_4877 ? _T_4544 : _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_241 = _T_4877 ? _T_4546 : _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_242 = _T_4877 ? _T_4548 : _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_243 = _T_4877 ? _T_4550 : _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_244 = _T_4877 ? _T_4552 : _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_245 = _T_4877 ? _T_4554 : _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_246 = _T_4877 ? _T_4556 : _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_247 = _T_4877 ? _T_4558 : _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_248 = _T_4877 ? _T_4560 : _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_249 = _T_4877 ? _T_4562 : _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_250 = _T_4877 ? _T_4564 : _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_251 = _T_4877 ? _T_4566 : _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_252 = _T_4877 ? _T_4568 : _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_253 = _T_4877 ? _T_4570 : _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_254 = _T_4877 ? _T_4572 : _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_255 = _T_4877 ? _T_4574 : _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_256 = _T_4877 ? _T_4576 : _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_257 = _T_4877 ? _T_4578 : _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_258 = _T_4877 ? _T_4580 : _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_259 = _T_4877 ? _T_4582 : _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_260 = _T_4877 ? _T_4584 : _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_261 = _T_4877 ? _T_4586 : _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_262 = _T_4877 ? _T_4588 : _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_263 = _T_4877 ? _T_4590 : _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_264 = _T_4877 ? _T_4592 : _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_265 = _T_4877 ? _T_4594 : _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_266 = _T_4877 ? _T_4596 : _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_267 = _T_4877 ? _T_4598 : _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_268 = _T_4877 ? _T_4600 : _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_269 = _T_4877 ? _T_4602 : _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_270 = _T_4877 ? _T_4604 : _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_271 = _T_4877 ? _T_4606 : _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_272 = _T_4877 ? _T_4608 : _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_273 = _T_4877 ? _T_4878 : _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_274 = _T_4877 ? _T_4879 : _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_275 = _T_4877 ? _T_4880 : _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_276 = _T_4877 ? _T_4881 : _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_277 = _T_4877 ? _T_4882 : _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_278 = _T_4877 ? _T_4883 : _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_279 = _T_4877 ? _T_4884 : _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_280 = _T_4877 ? _T_4885 : _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_281 = _T_4877 ? _T_4886 : _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_282 = _T_4877 ? _T_4887 : _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_283 = _T_4877 ? _T_4888 : _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_284 = _T_4877 ? _T_4889 : _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_285 = _T_4877 ? _T_4890 : _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_286 = _T_4877 ? _T_4891 : _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_287 = _T_4877 ? _T_4892 : _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _GEN_288 = _T_4877 ? _T_4893 : _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 812:52:@16635.4]
  assign _T_4916 = _T_3154 | _T_3160; // @[NV_NVDLA_CSC_wl.scala 816:29:@16750.4]
  assign _T_4917 = _T_3150[0]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16816.6]
  assign _T_4918 = _T_3150[1]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16817.6]
  assign _T_4919 = _T_3150[2]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16818.6]
  assign _T_4920 = _T_3150[3]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16819.6]
  assign _T_4921 = _T_3150[4]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16820.6]
  assign _T_4922 = _T_3150[5]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16821.6]
  assign _T_4923 = _T_3150[6]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16822.6]
  assign _T_4924 = _T_3150[7]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16823.6]
  assign _T_4925 = _T_3150[8]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16824.6]
  assign _T_4926 = _T_3150[9]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16825.6]
  assign _T_4927 = _T_3150[10]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16826.6]
  assign _T_4928 = _T_3150[11]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16827.6]
  assign _T_4929 = _T_3150[12]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16828.6]
  assign _T_4930 = _T_3150[13]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16829.6]
  assign _T_4931 = _T_3150[14]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16830.6]
  assign _T_4932 = _T_3150[15]; // @[NV_NVDLA_CSC_wl.scala 818:96:@16831.6]
  assign _GEN_289 = _T_4916 ? _T_4680 : _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_290 = _T_4916 ? _T_4682 : _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_291 = _T_4916 ? _T_4684 : _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_292 = _T_4916 ? _T_4686 : _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_293 = _T_4916 ? _T_4688 : _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_294 = _T_4916 ? _T_4690 : _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_295 = _T_4916 ? _T_4692 : _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_296 = _T_4916 ? _T_4694 : _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_297 = _T_4916 ? _T_4696 : _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_298 = _T_4916 ? _T_4698 : _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_299 = _T_4916 ? _T_4700 : _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_300 = _T_4916 ? _T_4702 : _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_301 = _T_4916 ? _T_4704 : _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_302 = _T_4916 ? _T_4706 : _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_303 = _T_4916 ? _T_4708 : _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_304 = _T_4916 ? _T_4710 : _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_305 = _T_4916 ? _T_4712 : _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_306 = _T_4916 ? _T_4714 : _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_307 = _T_4916 ? _T_4716 : _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_308 = _T_4916 ? _T_4718 : _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_309 = _T_4916 ? _T_4720 : _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_310 = _T_4916 ? _T_4722 : _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_311 = _T_4916 ? _T_4724 : _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_312 = _T_4916 ? _T_4726 : _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_313 = _T_4916 ? _T_4728 : _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_314 = _T_4916 ? _T_4730 : _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_315 = _T_4916 ? _T_4732 : _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_316 = _T_4916 ? _T_4734 : _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_317 = _T_4916 ? _T_4736 : _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_318 = _T_4916 ? _T_4738 : _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_319 = _T_4916 ? _T_4740 : _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_320 = _T_4916 ? _T_4742 : _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_321 = _T_4916 ? _T_4744 : _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_322 = _T_4916 ? _T_4746 : _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_323 = _T_4916 ? _T_4748 : _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_324 = _T_4916 ? _T_4750 : _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_325 = _T_4916 ? _T_4752 : _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_326 = _T_4916 ? _T_4754 : _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_327 = _T_4916 ? _T_4756 : _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_328 = _T_4916 ? _T_4758 : _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_329 = _T_4916 ? _T_4760 : _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_330 = _T_4916 ? _T_4762 : _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_331 = _T_4916 ? _T_4764 : _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_332 = _T_4916 ? _T_4766 : _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_333 = _T_4916 ? _T_4768 : _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_334 = _T_4916 ? _T_4770 : _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_335 = _T_4916 ? _T_4772 : _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_336 = _T_4916 ? _T_4774 : _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_337 = _T_4916 ? _T_4776 : _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_338 = _T_4916 ? _T_4778 : _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_339 = _T_4916 ? _T_4780 : _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_340 = _T_4916 ? _T_4782 : _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_341 = _T_4916 ? _T_4784 : _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_342 = _T_4916 ? _T_4786 : _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_343 = _T_4916 ? _T_4788 : _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_344 = _T_4916 ? _T_4790 : _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_345 = _T_4916 ? _T_4792 : _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_346 = _T_4916 ? _T_4794 : _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_347 = _T_4916 ? _T_4796 : _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_348 = _T_4916 ? _T_4798 : _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_349 = _T_4916 ? _T_4800 : _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_350 = _T_4916 ? _T_4802 : _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_351 = _T_4916 ? _T_4804 : _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_352 = _T_4916 ? _T_4806 : _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_353 = _T_4916 ? _T_4917 : _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_354 = _T_4916 ? _T_4918 : _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_355 = _T_4916 ? _T_4919 : _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_356 = _T_4916 ? _T_4920 : _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_357 = _T_4916 ? _T_4921 : _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_358 = _T_4916 ? _T_4922 : _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_359 = _T_4916 ? _T_4923 : _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_360 = _T_4916 ? _T_4924 : _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_361 = _T_4916 ? _T_4925 : _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_362 = _T_4916 ? _T_4926 : _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_363 = _T_4916 ? _T_4927 : _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_364 = _T_4916 ? _T_4928 : _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_365 = _T_4916 ? _T_4929 : _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_366 = _T_4916 ? _T_4930 : _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_367 = _T_4916 ? _T_4931 : _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign _GEN_368 = _T_4916 ? _T_4932 : _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 816:52:@16751.4]
  assign io_sc2cdma_wt_updt_valid = _T_863; // @[NV_NVDLA_CSC_wl.scala 212:30:@14411.4]
  assign io_sc2cdma_wt_updt_bits_entries = _T_867; // @[NV_NVDLA_CSC_wl.scala 213:37:@14417.4]
  assign io_sc2cdma_wt_updt_bits_kernels = 14'h0; // @[NV_NVDLA_CSC_wl.scala 217:37:@14424.4]
  assign io_sc2cdma_wmb_entries = _T_871; // @[NV_NVDLA_CSC_wl.scala 214:28:@14423.4]
  assign io_sc2buf_wt_rd_addr_valid = _T_1631; // @[NV_NVDLA_CSC_wl.scala 631:32:@15102.4]
  assign io_sc2buf_wt_rd_addr_bits = _T_1634; // @[NV_NVDLA_CSC_wl.scala 632:31:@15103.4]
  assign io_sc2mac_wt_a_valid = _T_3157; // @[NV_NVDLA_CSC_wl.scala 829:26:@17250.4]
  assign io_sc2mac_wt_a_bits_sel_0 = _T_4161_0; // @[NV_NVDLA_CSC_wl.scala 833:29:@17380.4]
  assign io_sc2mac_wt_a_bits_sel_1 = _T_4161_1; // @[NV_NVDLA_CSC_wl.scala 833:29:@17381.4]
  assign io_sc2mac_wt_a_bits_sel_2 = _T_4161_2; // @[NV_NVDLA_CSC_wl.scala 833:29:@17382.4]
  assign io_sc2mac_wt_a_bits_sel_3 = _T_4161_3; // @[NV_NVDLA_CSC_wl.scala 833:29:@17383.4]
  assign io_sc2mac_wt_a_bits_sel_4 = _T_4161_4; // @[NV_NVDLA_CSC_wl.scala 833:29:@17384.4]
  assign io_sc2mac_wt_a_bits_sel_5 = _T_4161_5; // @[NV_NVDLA_CSC_wl.scala 833:29:@17385.4]
  assign io_sc2mac_wt_a_bits_sel_6 = _T_4161_6; // @[NV_NVDLA_CSC_wl.scala 833:29:@17386.4]
  assign io_sc2mac_wt_a_bits_sel_7 = _T_4161_7; // @[NV_NVDLA_CSC_wl.scala 833:29:@17387.4]
  assign io_sc2mac_wt_a_bits_sel_8 = _T_4161_8; // @[NV_NVDLA_CSC_wl.scala 833:29:@17388.4]
  assign io_sc2mac_wt_a_bits_sel_9 = _T_4161_9; // @[NV_NVDLA_CSC_wl.scala 833:29:@17389.4]
  assign io_sc2mac_wt_a_bits_sel_10 = _T_4161_10; // @[NV_NVDLA_CSC_wl.scala 833:29:@17390.4]
  assign io_sc2mac_wt_a_bits_sel_11 = _T_4161_11; // @[NV_NVDLA_CSC_wl.scala 833:29:@17391.4]
  assign io_sc2mac_wt_a_bits_sel_12 = _T_4161_12; // @[NV_NVDLA_CSC_wl.scala 833:29:@17392.4]
  assign io_sc2mac_wt_a_bits_sel_13 = _T_4161_13; // @[NV_NVDLA_CSC_wl.scala 833:29:@17393.4]
  assign io_sc2mac_wt_a_bits_sel_14 = _T_4161_14; // @[NV_NVDLA_CSC_wl.scala 833:29:@17394.4]
  assign io_sc2mac_wt_a_bits_sel_15 = _T_4161_15; // @[NV_NVDLA_CSC_wl.scala 833:29:@17395.4]
  assign io_sc2mac_wt_a_bits_mask_0 = _T_3427_0; // @[NV_NVDLA_CSC_wl.scala 831:30:@17252.4]
  assign io_sc2mac_wt_a_bits_mask_1 = _T_3427_1; // @[NV_NVDLA_CSC_wl.scala 831:30:@17253.4]
  assign io_sc2mac_wt_a_bits_mask_2 = _T_3427_2; // @[NV_NVDLA_CSC_wl.scala 831:30:@17254.4]
  assign io_sc2mac_wt_a_bits_mask_3 = _T_3427_3; // @[NV_NVDLA_CSC_wl.scala 831:30:@17255.4]
  assign io_sc2mac_wt_a_bits_mask_4 = _T_3427_4; // @[NV_NVDLA_CSC_wl.scala 831:30:@17256.4]
  assign io_sc2mac_wt_a_bits_mask_5 = _T_3427_5; // @[NV_NVDLA_CSC_wl.scala 831:30:@17257.4]
  assign io_sc2mac_wt_a_bits_mask_6 = _T_3427_6; // @[NV_NVDLA_CSC_wl.scala 831:30:@17258.4]
  assign io_sc2mac_wt_a_bits_mask_7 = _T_3427_7; // @[NV_NVDLA_CSC_wl.scala 831:30:@17259.4]
  assign io_sc2mac_wt_a_bits_mask_8 = _T_3427_8; // @[NV_NVDLA_CSC_wl.scala 831:30:@17260.4]
  assign io_sc2mac_wt_a_bits_mask_9 = _T_3427_9; // @[NV_NVDLA_CSC_wl.scala 831:30:@17261.4]
  assign io_sc2mac_wt_a_bits_mask_10 = _T_3427_10; // @[NV_NVDLA_CSC_wl.scala 831:30:@17262.4]
  assign io_sc2mac_wt_a_bits_mask_11 = _T_3427_11; // @[NV_NVDLA_CSC_wl.scala 831:30:@17263.4]
  assign io_sc2mac_wt_a_bits_mask_12 = _T_3427_12; // @[NV_NVDLA_CSC_wl.scala 831:30:@17264.4]
  assign io_sc2mac_wt_a_bits_mask_13 = _T_3427_13; // @[NV_NVDLA_CSC_wl.scala 831:30:@17265.4]
  assign io_sc2mac_wt_a_bits_mask_14 = _T_3427_14; // @[NV_NVDLA_CSC_wl.scala 831:30:@17266.4]
  assign io_sc2mac_wt_a_bits_mask_15 = _T_3427_15; // @[NV_NVDLA_CSC_wl.scala 831:30:@17267.4]
  assign io_sc2mac_wt_a_bits_mask_16 = _T_3427_16; // @[NV_NVDLA_CSC_wl.scala 831:30:@17268.4]
  assign io_sc2mac_wt_a_bits_mask_17 = _T_3427_17; // @[NV_NVDLA_CSC_wl.scala 831:30:@17269.4]
  assign io_sc2mac_wt_a_bits_mask_18 = _T_3427_18; // @[NV_NVDLA_CSC_wl.scala 831:30:@17270.4]
  assign io_sc2mac_wt_a_bits_mask_19 = _T_3427_19; // @[NV_NVDLA_CSC_wl.scala 831:30:@17271.4]
  assign io_sc2mac_wt_a_bits_mask_20 = _T_3427_20; // @[NV_NVDLA_CSC_wl.scala 831:30:@17272.4]
  assign io_sc2mac_wt_a_bits_mask_21 = _T_3427_21; // @[NV_NVDLA_CSC_wl.scala 831:30:@17273.4]
  assign io_sc2mac_wt_a_bits_mask_22 = _T_3427_22; // @[NV_NVDLA_CSC_wl.scala 831:30:@17274.4]
  assign io_sc2mac_wt_a_bits_mask_23 = _T_3427_23; // @[NV_NVDLA_CSC_wl.scala 831:30:@17275.4]
  assign io_sc2mac_wt_a_bits_mask_24 = _T_3427_24; // @[NV_NVDLA_CSC_wl.scala 831:30:@17276.4]
  assign io_sc2mac_wt_a_bits_mask_25 = _T_3427_25; // @[NV_NVDLA_CSC_wl.scala 831:30:@17277.4]
  assign io_sc2mac_wt_a_bits_mask_26 = _T_3427_26; // @[NV_NVDLA_CSC_wl.scala 831:30:@17278.4]
  assign io_sc2mac_wt_a_bits_mask_27 = _T_3427_27; // @[NV_NVDLA_CSC_wl.scala 831:30:@17279.4]
  assign io_sc2mac_wt_a_bits_mask_28 = _T_3427_28; // @[NV_NVDLA_CSC_wl.scala 831:30:@17280.4]
  assign io_sc2mac_wt_a_bits_mask_29 = _T_3427_29; // @[NV_NVDLA_CSC_wl.scala 831:30:@17281.4]
  assign io_sc2mac_wt_a_bits_mask_30 = _T_3427_30; // @[NV_NVDLA_CSC_wl.scala 831:30:@17282.4]
  assign io_sc2mac_wt_a_bits_mask_31 = _T_3427_31; // @[NV_NVDLA_CSC_wl.scala 831:30:@17283.4]
  assign io_sc2mac_wt_a_bits_mask_32 = _T_3427_32; // @[NV_NVDLA_CSC_wl.scala 831:30:@17284.4]
  assign io_sc2mac_wt_a_bits_mask_33 = _T_3427_33; // @[NV_NVDLA_CSC_wl.scala 831:30:@17285.4]
  assign io_sc2mac_wt_a_bits_mask_34 = _T_3427_34; // @[NV_NVDLA_CSC_wl.scala 831:30:@17286.4]
  assign io_sc2mac_wt_a_bits_mask_35 = _T_3427_35; // @[NV_NVDLA_CSC_wl.scala 831:30:@17287.4]
  assign io_sc2mac_wt_a_bits_mask_36 = _T_3427_36; // @[NV_NVDLA_CSC_wl.scala 831:30:@17288.4]
  assign io_sc2mac_wt_a_bits_mask_37 = _T_3427_37; // @[NV_NVDLA_CSC_wl.scala 831:30:@17289.4]
  assign io_sc2mac_wt_a_bits_mask_38 = _T_3427_38; // @[NV_NVDLA_CSC_wl.scala 831:30:@17290.4]
  assign io_sc2mac_wt_a_bits_mask_39 = _T_3427_39; // @[NV_NVDLA_CSC_wl.scala 831:30:@17291.4]
  assign io_sc2mac_wt_a_bits_mask_40 = _T_3427_40; // @[NV_NVDLA_CSC_wl.scala 831:30:@17292.4]
  assign io_sc2mac_wt_a_bits_mask_41 = _T_3427_41; // @[NV_NVDLA_CSC_wl.scala 831:30:@17293.4]
  assign io_sc2mac_wt_a_bits_mask_42 = _T_3427_42; // @[NV_NVDLA_CSC_wl.scala 831:30:@17294.4]
  assign io_sc2mac_wt_a_bits_mask_43 = _T_3427_43; // @[NV_NVDLA_CSC_wl.scala 831:30:@17295.4]
  assign io_sc2mac_wt_a_bits_mask_44 = _T_3427_44; // @[NV_NVDLA_CSC_wl.scala 831:30:@17296.4]
  assign io_sc2mac_wt_a_bits_mask_45 = _T_3427_45; // @[NV_NVDLA_CSC_wl.scala 831:30:@17297.4]
  assign io_sc2mac_wt_a_bits_mask_46 = _T_3427_46; // @[NV_NVDLA_CSC_wl.scala 831:30:@17298.4]
  assign io_sc2mac_wt_a_bits_mask_47 = _T_3427_47; // @[NV_NVDLA_CSC_wl.scala 831:30:@17299.4]
  assign io_sc2mac_wt_a_bits_mask_48 = _T_3427_48; // @[NV_NVDLA_CSC_wl.scala 831:30:@17300.4]
  assign io_sc2mac_wt_a_bits_mask_49 = _T_3427_49; // @[NV_NVDLA_CSC_wl.scala 831:30:@17301.4]
  assign io_sc2mac_wt_a_bits_mask_50 = _T_3427_50; // @[NV_NVDLA_CSC_wl.scala 831:30:@17302.4]
  assign io_sc2mac_wt_a_bits_mask_51 = _T_3427_51; // @[NV_NVDLA_CSC_wl.scala 831:30:@17303.4]
  assign io_sc2mac_wt_a_bits_mask_52 = _T_3427_52; // @[NV_NVDLA_CSC_wl.scala 831:30:@17304.4]
  assign io_sc2mac_wt_a_bits_mask_53 = _T_3427_53; // @[NV_NVDLA_CSC_wl.scala 831:30:@17305.4]
  assign io_sc2mac_wt_a_bits_mask_54 = _T_3427_54; // @[NV_NVDLA_CSC_wl.scala 831:30:@17306.4]
  assign io_sc2mac_wt_a_bits_mask_55 = _T_3427_55; // @[NV_NVDLA_CSC_wl.scala 831:30:@17307.4]
  assign io_sc2mac_wt_a_bits_mask_56 = _T_3427_56; // @[NV_NVDLA_CSC_wl.scala 831:30:@17308.4]
  assign io_sc2mac_wt_a_bits_mask_57 = _T_3427_57; // @[NV_NVDLA_CSC_wl.scala 831:30:@17309.4]
  assign io_sc2mac_wt_a_bits_mask_58 = _T_3427_58; // @[NV_NVDLA_CSC_wl.scala 831:30:@17310.4]
  assign io_sc2mac_wt_a_bits_mask_59 = _T_3427_59; // @[NV_NVDLA_CSC_wl.scala 831:30:@17311.4]
  assign io_sc2mac_wt_a_bits_mask_60 = _T_3427_60; // @[NV_NVDLA_CSC_wl.scala 831:30:@17312.4]
  assign io_sc2mac_wt_a_bits_mask_61 = _T_3427_61; // @[NV_NVDLA_CSC_wl.scala 831:30:@17313.4]
  assign io_sc2mac_wt_a_bits_mask_62 = _T_3427_62; // @[NV_NVDLA_CSC_wl.scala 831:30:@17314.4]
  assign io_sc2mac_wt_a_bits_mask_63 = _T_3427_63; // @[NV_NVDLA_CSC_wl.scala 831:30:@17315.4]
  assign io_sc2mac_wt_a_bits_data_0 = _T_4344_0; // @[NV_NVDLA_CSC_wl.scala 835:30:@17412.4]
  assign io_sc2mac_wt_a_bits_data_1 = _T_4344_1; // @[NV_NVDLA_CSC_wl.scala 835:30:@17413.4]
  assign io_sc2mac_wt_a_bits_data_2 = _T_4344_2; // @[NV_NVDLA_CSC_wl.scala 835:30:@17414.4]
  assign io_sc2mac_wt_a_bits_data_3 = _T_4344_3; // @[NV_NVDLA_CSC_wl.scala 835:30:@17415.4]
  assign io_sc2mac_wt_a_bits_data_4 = _T_4344_4; // @[NV_NVDLA_CSC_wl.scala 835:30:@17416.4]
  assign io_sc2mac_wt_a_bits_data_5 = _T_4344_5; // @[NV_NVDLA_CSC_wl.scala 835:30:@17417.4]
  assign io_sc2mac_wt_a_bits_data_6 = _T_4344_6; // @[NV_NVDLA_CSC_wl.scala 835:30:@17418.4]
  assign io_sc2mac_wt_a_bits_data_7 = _T_4344_7; // @[NV_NVDLA_CSC_wl.scala 835:30:@17419.4]
  assign io_sc2mac_wt_a_bits_data_8 = _T_4344_8; // @[NV_NVDLA_CSC_wl.scala 835:30:@17420.4]
  assign io_sc2mac_wt_a_bits_data_9 = _T_4344_9; // @[NV_NVDLA_CSC_wl.scala 835:30:@17421.4]
  assign io_sc2mac_wt_a_bits_data_10 = _T_4344_10; // @[NV_NVDLA_CSC_wl.scala 835:30:@17422.4]
  assign io_sc2mac_wt_a_bits_data_11 = _T_4344_11; // @[NV_NVDLA_CSC_wl.scala 835:30:@17423.4]
  assign io_sc2mac_wt_a_bits_data_12 = _T_4344_12; // @[NV_NVDLA_CSC_wl.scala 835:30:@17424.4]
  assign io_sc2mac_wt_a_bits_data_13 = _T_4344_13; // @[NV_NVDLA_CSC_wl.scala 835:30:@17425.4]
  assign io_sc2mac_wt_a_bits_data_14 = _T_4344_14; // @[NV_NVDLA_CSC_wl.scala 835:30:@17426.4]
  assign io_sc2mac_wt_a_bits_data_15 = _T_4344_15; // @[NV_NVDLA_CSC_wl.scala 835:30:@17427.4]
  assign io_sc2mac_wt_a_bits_data_16 = _T_4344_16; // @[NV_NVDLA_CSC_wl.scala 835:30:@17428.4]
  assign io_sc2mac_wt_a_bits_data_17 = _T_4344_17; // @[NV_NVDLA_CSC_wl.scala 835:30:@17429.4]
  assign io_sc2mac_wt_a_bits_data_18 = _T_4344_18; // @[NV_NVDLA_CSC_wl.scala 835:30:@17430.4]
  assign io_sc2mac_wt_a_bits_data_19 = _T_4344_19; // @[NV_NVDLA_CSC_wl.scala 835:30:@17431.4]
  assign io_sc2mac_wt_a_bits_data_20 = _T_4344_20; // @[NV_NVDLA_CSC_wl.scala 835:30:@17432.4]
  assign io_sc2mac_wt_a_bits_data_21 = _T_4344_21; // @[NV_NVDLA_CSC_wl.scala 835:30:@17433.4]
  assign io_sc2mac_wt_a_bits_data_22 = _T_4344_22; // @[NV_NVDLA_CSC_wl.scala 835:30:@17434.4]
  assign io_sc2mac_wt_a_bits_data_23 = _T_4344_23; // @[NV_NVDLA_CSC_wl.scala 835:30:@17435.4]
  assign io_sc2mac_wt_a_bits_data_24 = _T_4344_24; // @[NV_NVDLA_CSC_wl.scala 835:30:@17436.4]
  assign io_sc2mac_wt_a_bits_data_25 = _T_4344_25; // @[NV_NVDLA_CSC_wl.scala 835:30:@17437.4]
  assign io_sc2mac_wt_a_bits_data_26 = _T_4344_26; // @[NV_NVDLA_CSC_wl.scala 835:30:@17438.4]
  assign io_sc2mac_wt_a_bits_data_27 = _T_4344_27; // @[NV_NVDLA_CSC_wl.scala 835:30:@17439.4]
  assign io_sc2mac_wt_a_bits_data_28 = _T_4344_28; // @[NV_NVDLA_CSC_wl.scala 835:30:@17440.4]
  assign io_sc2mac_wt_a_bits_data_29 = _T_4344_29; // @[NV_NVDLA_CSC_wl.scala 835:30:@17441.4]
  assign io_sc2mac_wt_a_bits_data_30 = _T_4344_30; // @[NV_NVDLA_CSC_wl.scala 835:30:@17442.4]
  assign io_sc2mac_wt_a_bits_data_31 = _T_4344_31; // @[NV_NVDLA_CSC_wl.scala 835:30:@17443.4]
  assign io_sc2mac_wt_a_bits_data_32 = _T_4344_32; // @[NV_NVDLA_CSC_wl.scala 835:30:@17444.4]
  assign io_sc2mac_wt_a_bits_data_33 = _T_4344_33; // @[NV_NVDLA_CSC_wl.scala 835:30:@17445.4]
  assign io_sc2mac_wt_a_bits_data_34 = _T_4344_34; // @[NV_NVDLA_CSC_wl.scala 835:30:@17446.4]
  assign io_sc2mac_wt_a_bits_data_35 = _T_4344_35; // @[NV_NVDLA_CSC_wl.scala 835:30:@17447.4]
  assign io_sc2mac_wt_a_bits_data_36 = _T_4344_36; // @[NV_NVDLA_CSC_wl.scala 835:30:@17448.4]
  assign io_sc2mac_wt_a_bits_data_37 = _T_4344_37; // @[NV_NVDLA_CSC_wl.scala 835:30:@17449.4]
  assign io_sc2mac_wt_a_bits_data_38 = _T_4344_38; // @[NV_NVDLA_CSC_wl.scala 835:30:@17450.4]
  assign io_sc2mac_wt_a_bits_data_39 = _T_4344_39; // @[NV_NVDLA_CSC_wl.scala 835:30:@17451.4]
  assign io_sc2mac_wt_a_bits_data_40 = _T_4344_40; // @[NV_NVDLA_CSC_wl.scala 835:30:@17452.4]
  assign io_sc2mac_wt_a_bits_data_41 = _T_4344_41; // @[NV_NVDLA_CSC_wl.scala 835:30:@17453.4]
  assign io_sc2mac_wt_a_bits_data_42 = _T_4344_42; // @[NV_NVDLA_CSC_wl.scala 835:30:@17454.4]
  assign io_sc2mac_wt_a_bits_data_43 = _T_4344_43; // @[NV_NVDLA_CSC_wl.scala 835:30:@17455.4]
  assign io_sc2mac_wt_a_bits_data_44 = _T_4344_44; // @[NV_NVDLA_CSC_wl.scala 835:30:@17456.4]
  assign io_sc2mac_wt_a_bits_data_45 = _T_4344_45; // @[NV_NVDLA_CSC_wl.scala 835:30:@17457.4]
  assign io_sc2mac_wt_a_bits_data_46 = _T_4344_46; // @[NV_NVDLA_CSC_wl.scala 835:30:@17458.4]
  assign io_sc2mac_wt_a_bits_data_47 = _T_4344_47; // @[NV_NVDLA_CSC_wl.scala 835:30:@17459.4]
  assign io_sc2mac_wt_a_bits_data_48 = _T_4344_48; // @[NV_NVDLA_CSC_wl.scala 835:30:@17460.4]
  assign io_sc2mac_wt_a_bits_data_49 = _T_4344_49; // @[NV_NVDLA_CSC_wl.scala 835:30:@17461.4]
  assign io_sc2mac_wt_a_bits_data_50 = _T_4344_50; // @[NV_NVDLA_CSC_wl.scala 835:30:@17462.4]
  assign io_sc2mac_wt_a_bits_data_51 = _T_4344_51; // @[NV_NVDLA_CSC_wl.scala 835:30:@17463.4]
  assign io_sc2mac_wt_a_bits_data_52 = _T_4344_52; // @[NV_NVDLA_CSC_wl.scala 835:30:@17464.4]
  assign io_sc2mac_wt_a_bits_data_53 = _T_4344_53; // @[NV_NVDLA_CSC_wl.scala 835:30:@17465.4]
  assign io_sc2mac_wt_a_bits_data_54 = _T_4344_54; // @[NV_NVDLA_CSC_wl.scala 835:30:@17466.4]
  assign io_sc2mac_wt_a_bits_data_55 = _T_4344_55; // @[NV_NVDLA_CSC_wl.scala 835:30:@17467.4]
  assign io_sc2mac_wt_a_bits_data_56 = _T_4344_56; // @[NV_NVDLA_CSC_wl.scala 835:30:@17468.4]
  assign io_sc2mac_wt_a_bits_data_57 = _T_4344_57; // @[NV_NVDLA_CSC_wl.scala 835:30:@17469.4]
  assign io_sc2mac_wt_a_bits_data_58 = _T_4344_58; // @[NV_NVDLA_CSC_wl.scala 835:30:@17470.4]
  assign io_sc2mac_wt_a_bits_data_59 = _T_4344_59; // @[NV_NVDLA_CSC_wl.scala 835:30:@17471.4]
  assign io_sc2mac_wt_a_bits_data_60 = _T_4344_60; // @[NV_NVDLA_CSC_wl.scala 835:30:@17472.4]
  assign io_sc2mac_wt_a_bits_data_61 = _T_4344_61; // @[NV_NVDLA_CSC_wl.scala 835:30:@17473.4]
  assign io_sc2mac_wt_a_bits_data_62 = _T_4344_62; // @[NV_NVDLA_CSC_wl.scala 835:30:@17474.4]
  assign io_sc2mac_wt_a_bits_data_63 = _T_4344_63; // @[NV_NVDLA_CSC_wl.scala 835:30:@17475.4]
  assign io_sc2mac_wt_b_valid = _T_3160; // @[NV_NVDLA_CSC_wl.scala 830:26:@17251.4]
  assign io_sc2mac_wt_b_bits_sel_0 = _T_4288_0; // @[NV_NVDLA_CSC_wl.scala 834:29:@17396.4]
  assign io_sc2mac_wt_b_bits_sel_1 = _T_4288_1; // @[NV_NVDLA_CSC_wl.scala 834:29:@17397.4]
  assign io_sc2mac_wt_b_bits_sel_2 = _T_4288_2; // @[NV_NVDLA_CSC_wl.scala 834:29:@17398.4]
  assign io_sc2mac_wt_b_bits_sel_3 = _T_4288_3; // @[NV_NVDLA_CSC_wl.scala 834:29:@17399.4]
  assign io_sc2mac_wt_b_bits_sel_4 = _T_4288_4; // @[NV_NVDLA_CSC_wl.scala 834:29:@17400.4]
  assign io_sc2mac_wt_b_bits_sel_5 = _T_4288_5; // @[NV_NVDLA_CSC_wl.scala 834:29:@17401.4]
  assign io_sc2mac_wt_b_bits_sel_6 = _T_4288_6; // @[NV_NVDLA_CSC_wl.scala 834:29:@17402.4]
  assign io_sc2mac_wt_b_bits_sel_7 = _T_4288_7; // @[NV_NVDLA_CSC_wl.scala 834:29:@17403.4]
  assign io_sc2mac_wt_b_bits_sel_8 = _T_4288_8; // @[NV_NVDLA_CSC_wl.scala 834:29:@17404.4]
  assign io_sc2mac_wt_b_bits_sel_9 = _T_4288_9; // @[NV_NVDLA_CSC_wl.scala 834:29:@17405.4]
  assign io_sc2mac_wt_b_bits_sel_10 = _T_4288_10; // @[NV_NVDLA_CSC_wl.scala 834:29:@17406.4]
  assign io_sc2mac_wt_b_bits_sel_11 = _T_4288_11; // @[NV_NVDLA_CSC_wl.scala 834:29:@17407.4]
  assign io_sc2mac_wt_b_bits_sel_12 = _T_4288_12; // @[NV_NVDLA_CSC_wl.scala 834:29:@17408.4]
  assign io_sc2mac_wt_b_bits_sel_13 = _T_4288_13; // @[NV_NVDLA_CSC_wl.scala 834:29:@17409.4]
  assign io_sc2mac_wt_b_bits_sel_14 = _T_4288_14; // @[NV_NVDLA_CSC_wl.scala 834:29:@17410.4]
  assign io_sc2mac_wt_b_bits_sel_15 = _T_4288_15; // @[NV_NVDLA_CSC_wl.scala 834:29:@17411.4]
  assign io_sc2mac_wt_b_bits_mask_0 = _T_3890_0; // @[NV_NVDLA_CSC_wl.scala 832:30:@17316.4]
  assign io_sc2mac_wt_b_bits_mask_1 = _T_3890_1; // @[NV_NVDLA_CSC_wl.scala 832:30:@17317.4]
  assign io_sc2mac_wt_b_bits_mask_2 = _T_3890_2; // @[NV_NVDLA_CSC_wl.scala 832:30:@17318.4]
  assign io_sc2mac_wt_b_bits_mask_3 = _T_3890_3; // @[NV_NVDLA_CSC_wl.scala 832:30:@17319.4]
  assign io_sc2mac_wt_b_bits_mask_4 = _T_3890_4; // @[NV_NVDLA_CSC_wl.scala 832:30:@17320.4]
  assign io_sc2mac_wt_b_bits_mask_5 = _T_3890_5; // @[NV_NVDLA_CSC_wl.scala 832:30:@17321.4]
  assign io_sc2mac_wt_b_bits_mask_6 = _T_3890_6; // @[NV_NVDLA_CSC_wl.scala 832:30:@17322.4]
  assign io_sc2mac_wt_b_bits_mask_7 = _T_3890_7; // @[NV_NVDLA_CSC_wl.scala 832:30:@17323.4]
  assign io_sc2mac_wt_b_bits_mask_8 = _T_3890_8; // @[NV_NVDLA_CSC_wl.scala 832:30:@17324.4]
  assign io_sc2mac_wt_b_bits_mask_9 = _T_3890_9; // @[NV_NVDLA_CSC_wl.scala 832:30:@17325.4]
  assign io_sc2mac_wt_b_bits_mask_10 = _T_3890_10; // @[NV_NVDLA_CSC_wl.scala 832:30:@17326.4]
  assign io_sc2mac_wt_b_bits_mask_11 = _T_3890_11; // @[NV_NVDLA_CSC_wl.scala 832:30:@17327.4]
  assign io_sc2mac_wt_b_bits_mask_12 = _T_3890_12; // @[NV_NVDLA_CSC_wl.scala 832:30:@17328.4]
  assign io_sc2mac_wt_b_bits_mask_13 = _T_3890_13; // @[NV_NVDLA_CSC_wl.scala 832:30:@17329.4]
  assign io_sc2mac_wt_b_bits_mask_14 = _T_3890_14; // @[NV_NVDLA_CSC_wl.scala 832:30:@17330.4]
  assign io_sc2mac_wt_b_bits_mask_15 = _T_3890_15; // @[NV_NVDLA_CSC_wl.scala 832:30:@17331.4]
  assign io_sc2mac_wt_b_bits_mask_16 = _T_3890_16; // @[NV_NVDLA_CSC_wl.scala 832:30:@17332.4]
  assign io_sc2mac_wt_b_bits_mask_17 = _T_3890_17; // @[NV_NVDLA_CSC_wl.scala 832:30:@17333.4]
  assign io_sc2mac_wt_b_bits_mask_18 = _T_3890_18; // @[NV_NVDLA_CSC_wl.scala 832:30:@17334.4]
  assign io_sc2mac_wt_b_bits_mask_19 = _T_3890_19; // @[NV_NVDLA_CSC_wl.scala 832:30:@17335.4]
  assign io_sc2mac_wt_b_bits_mask_20 = _T_3890_20; // @[NV_NVDLA_CSC_wl.scala 832:30:@17336.4]
  assign io_sc2mac_wt_b_bits_mask_21 = _T_3890_21; // @[NV_NVDLA_CSC_wl.scala 832:30:@17337.4]
  assign io_sc2mac_wt_b_bits_mask_22 = _T_3890_22; // @[NV_NVDLA_CSC_wl.scala 832:30:@17338.4]
  assign io_sc2mac_wt_b_bits_mask_23 = _T_3890_23; // @[NV_NVDLA_CSC_wl.scala 832:30:@17339.4]
  assign io_sc2mac_wt_b_bits_mask_24 = _T_3890_24; // @[NV_NVDLA_CSC_wl.scala 832:30:@17340.4]
  assign io_sc2mac_wt_b_bits_mask_25 = _T_3890_25; // @[NV_NVDLA_CSC_wl.scala 832:30:@17341.4]
  assign io_sc2mac_wt_b_bits_mask_26 = _T_3890_26; // @[NV_NVDLA_CSC_wl.scala 832:30:@17342.4]
  assign io_sc2mac_wt_b_bits_mask_27 = _T_3890_27; // @[NV_NVDLA_CSC_wl.scala 832:30:@17343.4]
  assign io_sc2mac_wt_b_bits_mask_28 = _T_3890_28; // @[NV_NVDLA_CSC_wl.scala 832:30:@17344.4]
  assign io_sc2mac_wt_b_bits_mask_29 = _T_3890_29; // @[NV_NVDLA_CSC_wl.scala 832:30:@17345.4]
  assign io_sc2mac_wt_b_bits_mask_30 = _T_3890_30; // @[NV_NVDLA_CSC_wl.scala 832:30:@17346.4]
  assign io_sc2mac_wt_b_bits_mask_31 = _T_3890_31; // @[NV_NVDLA_CSC_wl.scala 832:30:@17347.4]
  assign io_sc2mac_wt_b_bits_mask_32 = _T_3890_32; // @[NV_NVDLA_CSC_wl.scala 832:30:@17348.4]
  assign io_sc2mac_wt_b_bits_mask_33 = _T_3890_33; // @[NV_NVDLA_CSC_wl.scala 832:30:@17349.4]
  assign io_sc2mac_wt_b_bits_mask_34 = _T_3890_34; // @[NV_NVDLA_CSC_wl.scala 832:30:@17350.4]
  assign io_sc2mac_wt_b_bits_mask_35 = _T_3890_35; // @[NV_NVDLA_CSC_wl.scala 832:30:@17351.4]
  assign io_sc2mac_wt_b_bits_mask_36 = _T_3890_36; // @[NV_NVDLA_CSC_wl.scala 832:30:@17352.4]
  assign io_sc2mac_wt_b_bits_mask_37 = _T_3890_37; // @[NV_NVDLA_CSC_wl.scala 832:30:@17353.4]
  assign io_sc2mac_wt_b_bits_mask_38 = _T_3890_38; // @[NV_NVDLA_CSC_wl.scala 832:30:@17354.4]
  assign io_sc2mac_wt_b_bits_mask_39 = _T_3890_39; // @[NV_NVDLA_CSC_wl.scala 832:30:@17355.4]
  assign io_sc2mac_wt_b_bits_mask_40 = _T_3890_40; // @[NV_NVDLA_CSC_wl.scala 832:30:@17356.4]
  assign io_sc2mac_wt_b_bits_mask_41 = _T_3890_41; // @[NV_NVDLA_CSC_wl.scala 832:30:@17357.4]
  assign io_sc2mac_wt_b_bits_mask_42 = _T_3890_42; // @[NV_NVDLA_CSC_wl.scala 832:30:@17358.4]
  assign io_sc2mac_wt_b_bits_mask_43 = _T_3890_43; // @[NV_NVDLA_CSC_wl.scala 832:30:@17359.4]
  assign io_sc2mac_wt_b_bits_mask_44 = _T_3890_44; // @[NV_NVDLA_CSC_wl.scala 832:30:@17360.4]
  assign io_sc2mac_wt_b_bits_mask_45 = _T_3890_45; // @[NV_NVDLA_CSC_wl.scala 832:30:@17361.4]
  assign io_sc2mac_wt_b_bits_mask_46 = _T_3890_46; // @[NV_NVDLA_CSC_wl.scala 832:30:@17362.4]
  assign io_sc2mac_wt_b_bits_mask_47 = _T_3890_47; // @[NV_NVDLA_CSC_wl.scala 832:30:@17363.4]
  assign io_sc2mac_wt_b_bits_mask_48 = _T_3890_48; // @[NV_NVDLA_CSC_wl.scala 832:30:@17364.4]
  assign io_sc2mac_wt_b_bits_mask_49 = _T_3890_49; // @[NV_NVDLA_CSC_wl.scala 832:30:@17365.4]
  assign io_sc2mac_wt_b_bits_mask_50 = _T_3890_50; // @[NV_NVDLA_CSC_wl.scala 832:30:@17366.4]
  assign io_sc2mac_wt_b_bits_mask_51 = _T_3890_51; // @[NV_NVDLA_CSC_wl.scala 832:30:@17367.4]
  assign io_sc2mac_wt_b_bits_mask_52 = _T_3890_52; // @[NV_NVDLA_CSC_wl.scala 832:30:@17368.4]
  assign io_sc2mac_wt_b_bits_mask_53 = _T_3890_53; // @[NV_NVDLA_CSC_wl.scala 832:30:@17369.4]
  assign io_sc2mac_wt_b_bits_mask_54 = _T_3890_54; // @[NV_NVDLA_CSC_wl.scala 832:30:@17370.4]
  assign io_sc2mac_wt_b_bits_mask_55 = _T_3890_55; // @[NV_NVDLA_CSC_wl.scala 832:30:@17371.4]
  assign io_sc2mac_wt_b_bits_mask_56 = _T_3890_56; // @[NV_NVDLA_CSC_wl.scala 832:30:@17372.4]
  assign io_sc2mac_wt_b_bits_mask_57 = _T_3890_57; // @[NV_NVDLA_CSC_wl.scala 832:30:@17373.4]
  assign io_sc2mac_wt_b_bits_mask_58 = _T_3890_58; // @[NV_NVDLA_CSC_wl.scala 832:30:@17374.4]
  assign io_sc2mac_wt_b_bits_mask_59 = _T_3890_59; // @[NV_NVDLA_CSC_wl.scala 832:30:@17375.4]
  assign io_sc2mac_wt_b_bits_mask_60 = _T_3890_60; // @[NV_NVDLA_CSC_wl.scala 832:30:@17376.4]
  assign io_sc2mac_wt_b_bits_mask_61 = _T_3890_61; // @[NV_NVDLA_CSC_wl.scala 832:30:@17377.4]
  assign io_sc2mac_wt_b_bits_mask_62 = _T_3890_62; // @[NV_NVDLA_CSC_wl.scala 832:30:@17378.4]
  assign io_sc2mac_wt_b_bits_mask_63 = _T_3890_63; // @[NV_NVDLA_CSC_wl.scala 832:30:@17379.4]
  assign io_sc2mac_wt_b_bits_data_0 = _T_4414_0; // @[NV_NVDLA_CSC_wl.scala 836:30:@17476.4]
  assign io_sc2mac_wt_b_bits_data_1 = _T_4414_1; // @[NV_NVDLA_CSC_wl.scala 836:30:@17477.4]
  assign io_sc2mac_wt_b_bits_data_2 = _T_4414_2; // @[NV_NVDLA_CSC_wl.scala 836:30:@17478.4]
  assign io_sc2mac_wt_b_bits_data_3 = _T_4414_3; // @[NV_NVDLA_CSC_wl.scala 836:30:@17479.4]
  assign io_sc2mac_wt_b_bits_data_4 = _T_4414_4; // @[NV_NVDLA_CSC_wl.scala 836:30:@17480.4]
  assign io_sc2mac_wt_b_bits_data_5 = _T_4414_5; // @[NV_NVDLA_CSC_wl.scala 836:30:@17481.4]
  assign io_sc2mac_wt_b_bits_data_6 = _T_4414_6; // @[NV_NVDLA_CSC_wl.scala 836:30:@17482.4]
  assign io_sc2mac_wt_b_bits_data_7 = _T_4414_7; // @[NV_NVDLA_CSC_wl.scala 836:30:@17483.4]
  assign io_sc2mac_wt_b_bits_data_8 = _T_4414_8; // @[NV_NVDLA_CSC_wl.scala 836:30:@17484.4]
  assign io_sc2mac_wt_b_bits_data_9 = _T_4414_9; // @[NV_NVDLA_CSC_wl.scala 836:30:@17485.4]
  assign io_sc2mac_wt_b_bits_data_10 = _T_4414_10; // @[NV_NVDLA_CSC_wl.scala 836:30:@17486.4]
  assign io_sc2mac_wt_b_bits_data_11 = _T_4414_11; // @[NV_NVDLA_CSC_wl.scala 836:30:@17487.4]
  assign io_sc2mac_wt_b_bits_data_12 = _T_4414_12; // @[NV_NVDLA_CSC_wl.scala 836:30:@17488.4]
  assign io_sc2mac_wt_b_bits_data_13 = _T_4414_13; // @[NV_NVDLA_CSC_wl.scala 836:30:@17489.4]
  assign io_sc2mac_wt_b_bits_data_14 = _T_4414_14; // @[NV_NVDLA_CSC_wl.scala 836:30:@17490.4]
  assign io_sc2mac_wt_b_bits_data_15 = _T_4414_15; // @[NV_NVDLA_CSC_wl.scala 836:30:@17491.4]
  assign io_sc2mac_wt_b_bits_data_16 = _T_4414_16; // @[NV_NVDLA_CSC_wl.scala 836:30:@17492.4]
  assign io_sc2mac_wt_b_bits_data_17 = _T_4414_17; // @[NV_NVDLA_CSC_wl.scala 836:30:@17493.4]
  assign io_sc2mac_wt_b_bits_data_18 = _T_4414_18; // @[NV_NVDLA_CSC_wl.scala 836:30:@17494.4]
  assign io_sc2mac_wt_b_bits_data_19 = _T_4414_19; // @[NV_NVDLA_CSC_wl.scala 836:30:@17495.4]
  assign io_sc2mac_wt_b_bits_data_20 = _T_4414_20; // @[NV_NVDLA_CSC_wl.scala 836:30:@17496.4]
  assign io_sc2mac_wt_b_bits_data_21 = _T_4414_21; // @[NV_NVDLA_CSC_wl.scala 836:30:@17497.4]
  assign io_sc2mac_wt_b_bits_data_22 = _T_4414_22; // @[NV_NVDLA_CSC_wl.scala 836:30:@17498.4]
  assign io_sc2mac_wt_b_bits_data_23 = _T_4414_23; // @[NV_NVDLA_CSC_wl.scala 836:30:@17499.4]
  assign io_sc2mac_wt_b_bits_data_24 = _T_4414_24; // @[NV_NVDLA_CSC_wl.scala 836:30:@17500.4]
  assign io_sc2mac_wt_b_bits_data_25 = _T_4414_25; // @[NV_NVDLA_CSC_wl.scala 836:30:@17501.4]
  assign io_sc2mac_wt_b_bits_data_26 = _T_4414_26; // @[NV_NVDLA_CSC_wl.scala 836:30:@17502.4]
  assign io_sc2mac_wt_b_bits_data_27 = _T_4414_27; // @[NV_NVDLA_CSC_wl.scala 836:30:@17503.4]
  assign io_sc2mac_wt_b_bits_data_28 = _T_4414_28; // @[NV_NVDLA_CSC_wl.scala 836:30:@17504.4]
  assign io_sc2mac_wt_b_bits_data_29 = _T_4414_29; // @[NV_NVDLA_CSC_wl.scala 836:30:@17505.4]
  assign io_sc2mac_wt_b_bits_data_30 = _T_4414_30; // @[NV_NVDLA_CSC_wl.scala 836:30:@17506.4]
  assign io_sc2mac_wt_b_bits_data_31 = _T_4414_31; // @[NV_NVDLA_CSC_wl.scala 836:30:@17507.4]
  assign io_sc2mac_wt_b_bits_data_32 = _T_4414_32; // @[NV_NVDLA_CSC_wl.scala 836:30:@17508.4]
  assign io_sc2mac_wt_b_bits_data_33 = _T_4414_33; // @[NV_NVDLA_CSC_wl.scala 836:30:@17509.4]
  assign io_sc2mac_wt_b_bits_data_34 = _T_4414_34; // @[NV_NVDLA_CSC_wl.scala 836:30:@17510.4]
  assign io_sc2mac_wt_b_bits_data_35 = _T_4414_35; // @[NV_NVDLA_CSC_wl.scala 836:30:@17511.4]
  assign io_sc2mac_wt_b_bits_data_36 = _T_4414_36; // @[NV_NVDLA_CSC_wl.scala 836:30:@17512.4]
  assign io_sc2mac_wt_b_bits_data_37 = _T_4414_37; // @[NV_NVDLA_CSC_wl.scala 836:30:@17513.4]
  assign io_sc2mac_wt_b_bits_data_38 = _T_4414_38; // @[NV_NVDLA_CSC_wl.scala 836:30:@17514.4]
  assign io_sc2mac_wt_b_bits_data_39 = _T_4414_39; // @[NV_NVDLA_CSC_wl.scala 836:30:@17515.4]
  assign io_sc2mac_wt_b_bits_data_40 = _T_4414_40; // @[NV_NVDLA_CSC_wl.scala 836:30:@17516.4]
  assign io_sc2mac_wt_b_bits_data_41 = _T_4414_41; // @[NV_NVDLA_CSC_wl.scala 836:30:@17517.4]
  assign io_sc2mac_wt_b_bits_data_42 = _T_4414_42; // @[NV_NVDLA_CSC_wl.scala 836:30:@17518.4]
  assign io_sc2mac_wt_b_bits_data_43 = _T_4414_43; // @[NV_NVDLA_CSC_wl.scala 836:30:@17519.4]
  assign io_sc2mac_wt_b_bits_data_44 = _T_4414_44; // @[NV_NVDLA_CSC_wl.scala 836:30:@17520.4]
  assign io_sc2mac_wt_b_bits_data_45 = _T_4414_45; // @[NV_NVDLA_CSC_wl.scala 836:30:@17521.4]
  assign io_sc2mac_wt_b_bits_data_46 = _T_4414_46; // @[NV_NVDLA_CSC_wl.scala 836:30:@17522.4]
  assign io_sc2mac_wt_b_bits_data_47 = _T_4414_47; // @[NV_NVDLA_CSC_wl.scala 836:30:@17523.4]
  assign io_sc2mac_wt_b_bits_data_48 = _T_4414_48; // @[NV_NVDLA_CSC_wl.scala 836:30:@17524.4]
  assign io_sc2mac_wt_b_bits_data_49 = _T_4414_49; // @[NV_NVDLA_CSC_wl.scala 836:30:@17525.4]
  assign io_sc2mac_wt_b_bits_data_50 = _T_4414_50; // @[NV_NVDLA_CSC_wl.scala 836:30:@17526.4]
  assign io_sc2mac_wt_b_bits_data_51 = _T_4414_51; // @[NV_NVDLA_CSC_wl.scala 836:30:@17527.4]
  assign io_sc2mac_wt_b_bits_data_52 = _T_4414_52; // @[NV_NVDLA_CSC_wl.scala 836:30:@17528.4]
  assign io_sc2mac_wt_b_bits_data_53 = _T_4414_53; // @[NV_NVDLA_CSC_wl.scala 836:30:@17529.4]
  assign io_sc2mac_wt_b_bits_data_54 = _T_4414_54; // @[NV_NVDLA_CSC_wl.scala 836:30:@17530.4]
  assign io_sc2mac_wt_b_bits_data_55 = _T_4414_55; // @[NV_NVDLA_CSC_wl.scala 836:30:@17531.4]
  assign io_sc2mac_wt_b_bits_data_56 = _T_4414_56; // @[NV_NVDLA_CSC_wl.scala 836:30:@17532.4]
  assign io_sc2mac_wt_b_bits_data_57 = _T_4414_57; // @[NV_NVDLA_CSC_wl.scala 836:30:@17533.4]
  assign io_sc2mac_wt_b_bits_data_58 = _T_4414_58; // @[NV_NVDLA_CSC_wl.scala 836:30:@17534.4]
  assign io_sc2mac_wt_b_bits_data_59 = _T_4414_59; // @[NV_NVDLA_CSC_wl.scala 836:30:@17535.4]
  assign io_sc2mac_wt_b_bits_data_60 = _T_4414_60; // @[NV_NVDLA_CSC_wl.scala 836:30:@17536.4]
  assign io_sc2mac_wt_b_bits_data_61 = _T_4414_61; // @[NV_NVDLA_CSC_wl.scala 836:30:@17537.4]
  assign io_sc2mac_wt_b_bits_data_62 = _T_4414_62; // @[NV_NVDLA_CSC_wl.scala 836:30:@17538.4]
  assign io_sc2mac_wt_b_bits_data_63 = _T_4414_63; // @[NV_NVDLA_CSC_wl.scala 836:30:@17539.4]
  assign NV_NVDLA_CSC_WL_dec_reset = reset; // @[:@15838.4]
  assign NV_NVDLA_CSC_WL_dec_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CSC_wl.scala 779:29:@15839.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_valid = _T_2472; // @[NV_NVDLA_CSC_wl.scala 783:26:@15969.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_0 = _T_2739_0; // @[NV_NVDLA_CSC_wl.scala 781:30:@15904.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_1 = _T_2739_1; // @[NV_NVDLA_CSC_wl.scala 781:30:@15905.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_2 = _T_2739_2; // @[NV_NVDLA_CSC_wl.scala 781:30:@15906.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_3 = _T_2739_3; // @[NV_NVDLA_CSC_wl.scala 781:30:@15907.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_4 = _T_2739_4; // @[NV_NVDLA_CSC_wl.scala 781:30:@15908.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_5 = _T_2739_5; // @[NV_NVDLA_CSC_wl.scala 781:30:@15909.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_6 = _T_2739_6; // @[NV_NVDLA_CSC_wl.scala 781:30:@15910.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_7 = _T_2739_7; // @[NV_NVDLA_CSC_wl.scala 781:30:@15911.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_8 = _T_2739_8; // @[NV_NVDLA_CSC_wl.scala 781:30:@15912.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_9 = _T_2739_9; // @[NV_NVDLA_CSC_wl.scala 781:30:@15913.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_10 = _T_2739_10; // @[NV_NVDLA_CSC_wl.scala 781:30:@15914.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_11 = _T_2739_11; // @[NV_NVDLA_CSC_wl.scala 781:30:@15915.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_12 = _T_2739_12; // @[NV_NVDLA_CSC_wl.scala 781:30:@15916.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_13 = _T_2739_13; // @[NV_NVDLA_CSC_wl.scala 781:30:@15917.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_14 = _T_2739_14; // @[NV_NVDLA_CSC_wl.scala 781:30:@15918.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_15 = _T_2739_15; // @[NV_NVDLA_CSC_wl.scala 781:30:@15919.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_16 = _T_2739_16; // @[NV_NVDLA_CSC_wl.scala 781:30:@15920.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_17 = _T_2739_17; // @[NV_NVDLA_CSC_wl.scala 781:30:@15921.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_18 = _T_2739_18; // @[NV_NVDLA_CSC_wl.scala 781:30:@15922.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_19 = _T_2739_19; // @[NV_NVDLA_CSC_wl.scala 781:30:@15923.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_20 = _T_2739_20; // @[NV_NVDLA_CSC_wl.scala 781:30:@15924.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_21 = _T_2739_21; // @[NV_NVDLA_CSC_wl.scala 781:30:@15925.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_22 = _T_2739_22; // @[NV_NVDLA_CSC_wl.scala 781:30:@15926.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_23 = _T_2739_23; // @[NV_NVDLA_CSC_wl.scala 781:30:@15927.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_24 = _T_2739_24; // @[NV_NVDLA_CSC_wl.scala 781:30:@15928.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_25 = _T_2739_25; // @[NV_NVDLA_CSC_wl.scala 781:30:@15929.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_26 = _T_2739_26; // @[NV_NVDLA_CSC_wl.scala 781:30:@15930.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_27 = _T_2739_27; // @[NV_NVDLA_CSC_wl.scala 781:30:@15931.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_28 = _T_2739_28; // @[NV_NVDLA_CSC_wl.scala 781:30:@15932.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_29 = _T_2739_29; // @[NV_NVDLA_CSC_wl.scala 781:30:@15933.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_30 = _T_2739_30; // @[NV_NVDLA_CSC_wl.scala 781:30:@15934.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_31 = _T_2739_31; // @[NV_NVDLA_CSC_wl.scala 781:30:@15935.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_32 = _T_2739_32; // @[NV_NVDLA_CSC_wl.scala 781:30:@15936.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_33 = _T_2739_33; // @[NV_NVDLA_CSC_wl.scala 781:30:@15937.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_34 = _T_2739_34; // @[NV_NVDLA_CSC_wl.scala 781:30:@15938.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_35 = _T_2739_35; // @[NV_NVDLA_CSC_wl.scala 781:30:@15939.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_36 = _T_2739_36; // @[NV_NVDLA_CSC_wl.scala 781:30:@15940.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_37 = _T_2739_37; // @[NV_NVDLA_CSC_wl.scala 781:30:@15941.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_38 = _T_2739_38; // @[NV_NVDLA_CSC_wl.scala 781:30:@15942.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_39 = _T_2739_39; // @[NV_NVDLA_CSC_wl.scala 781:30:@15943.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_40 = _T_2739_40; // @[NV_NVDLA_CSC_wl.scala 781:30:@15944.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_41 = _T_2739_41; // @[NV_NVDLA_CSC_wl.scala 781:30:@15945.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_42 = _T_2739_42; // @[NV_NVDLA_CSC_wl.scala 781:30:@15946.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_43 = _T_2739_43; // @[NV_NVDLA_CSC_wl.scala 781:30:@15947.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_44 = _T_2739_44; // @[NV_NVDLA_CSC_wl.scala 781:30:@15948.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_45 = _T_2739_45; // @[NV_NVDLA_CSC_wl.scala 781:30:@15949.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_46 = _T_2739_46; // @[NV_NVDLA_CSC_wl.scala 781:30:@15950.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_47 = _T_2739_47; // @[NV_NVDLA_CSC_wl.scala 781:30:@15951.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_48 = _T_2739_48; // @[NV_NVDLA_CSC_wl.scala 781:30:@15952.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_49 = _T_2739_49; // @[NV_NVDLA_CSC_wl.scala 781:30:@15953.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_50 = _T_2739_50; // @[NV_NVDLA_CSC_wl.scala 781:30:@15954.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_51 = _T_2739_51; // @[NV_NVDLA_CSC_wl.scala 781:30:@15955.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_52 = _T_2739_52; // @[NV_NVDLA_CSC_wl.scala 781:30:@15956.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_53 = _T_2739_53; // @[NV_NVDLA_CSC_wl.scala 781:30:@15957.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_54 = _T_2739_54; // @[NV_NVDLA_CSC_wl.scala 781:30:@15958.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_55 = _T_2739_55; // @[NV_NVDLA_CSC_wl.scala 781:30:@15959.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_56 = _T_2739_56; // @[NV_NVDLA_CSC_wl.scala 781:30:@15960.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_57 = _T_2739_57; // @[NV_NVDLA_CSC_wl.scala 781:30:@15961.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_58 = _T_2739_58; // @[NV_NVDLA_CSC_wl.scala 781:30:@15962.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_59 = _T_2739_59; // @[NV_NVDLA_CSC_wl.scala 781:30:@15963.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_60 = _T_2739_60; // @[NV_NVDLA_CSC_wl.scala 781:30:@15964.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_61 = _T_2739_61; // @[NV_NVDLA_CSC_wl.scala 781:30:@15965.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_62 = _T_2739_62; // @[NV_NVDLA_CSC_wl.scala 781:30:@15966.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_mask_63 = _T_2739_63; // @[NV_NVDLA_CSC_wl.scala 781:30:@15967.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_0 = _T_2095_0; // @[NV_NVDLA_CSC_wl.scala 780:30:@15840.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_1 = _T_2095_1; // @[NV_NVDLA_CSC_wl.scala 780:30:@15841.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_2 = _T_2095_2; // @[NV_NVDLA_CSC_wl.scala 780:30:@15842.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_3 = _T_2095_3; // @[NV_NVDLA_CSC_wl.scala 780:30:@15843.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_4 = _T_2095_4; // @[NV_NVDLA_CSC_wl.scala 780:30:@15844.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_5 = _T_2095_5; // @[NV_NVDLA_CSC_wl.scala 780:30:@15845.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_6 = _T_2095_6; // @[NV_NVDLA_CSC_wl.scala 780:30:@15846.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_7 = _T_2095_7; // @[NV_NVDLA_CSC_wl.scala 780:30:@15847.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_8 = _T_2095_8; // @[NV_NVDLA_CSC_wl.scala 780:30:@15848.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_9 = _T_2095_9; // @[NV_NVDLA_CSC_wl.scala 780:30:@15849.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_10 = _T_2095_10; // @[NV_NVDLA_CSC_wl.scala 780:30:@15850.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_11 = _T_2095_11; // @[NV_NVDLA_CSC_wl.scala 780:30:@15851.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_12 = _T_2095_12; // @[NV_NVDLA_CSC_wl.scala 780:30:@15852.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_13 = _T_2095_13; // @[NV_NVDLA_CSC_wl.scala 780:30:@15853.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_14 = _T_2095_14; // @[NV_NVDLA_CSC_wl.scala 780:30:@15854.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_15 = _T_2095_15; // @[NV_NVDLA_CSC_wl.scala 780:30:@15855.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_16 = _T_2095_16; // @[NV_NVDLA_CSC_wl.scala 780:30:@15856.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_17 = _T_2095_17; // @[NV_NVDLA_CSC_wl.scala 780:30:@15857.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_18 = _T_2095_18; // @[NV_NVDLA_CSC_wl.scala 780:30:@15858.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_19 = _T_2095_19; // @[NV_NVDLA_CSC_wl.scala 780:30:@15859.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_20 = _T_2095_20; // @[NV_NVDLA_CSC_wl.scala 780:30:@15860.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_21 = _T_2095_21; // @[NV_NVDLA_CSC_wl.scala 780:30:@15861.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_22 = _T_2095_22; // @[NV_NVDLA_CSC_wl.scala 780:30:@15862.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_23 = _T_2095_23; // @[NV_NVDLA_CSC_wl.scala 780:30:@15863.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_24 = _T_2095_24; // @[NV_NVDLA_CSC_wl.scala 780:30:@15864.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_25 = _T_2095_25; // @[NV_NVDLA_CSC_wl.scala 780:30:@15865.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_26 = _T_2095_26; // @[NV_NVDLA_CSC_wl.scala 780:30:@15866.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_27 = _T_2095_27; // @[NV_NVDLA_CSC_wl.scala 780:30:@15867.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_28 = _T_2095_28; // @[NV_NVDLA_CSC_wl.scala 780:30:@15868.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_29 = _T_2095_29; // @[NV_NVDLA_CSC_wl.scala 780:30:@15869.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_30 = _T_2095_30; // @[NV_NVDLA_CSC_wl.scala 780:30:@15870.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_31 = _T_2095_31; // @[NV_NVDLA_CSC_wl.scala 780:30:@15871.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_32 = _T_2095_32; // @[NV_NVDLA_CSC_wl.scala 780:30:@15872.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_33 = _T_2095_33; // @[NV_NVDLA_CSC_wl.scala 780:30:@15873.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_34 = _T_2095_34; // @[NV_NVDLA_CSC_wl.scala 780:30:@15874.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_35 = _T_2095_35; // @[NV_NVDLA_CSC_wl.scala 780:30:@15875.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_36 = _T_2095_36; // @[NV_NVDLA_CSC_wl.scala 780:30:@15876.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_37 = _T_2095_37; // @[NV_NVDLA_CSC_wl.scala 780:30:@15877.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_38 = _T_2095_38; // @[NV_NVDLA_CSC_wl.scala 780:30:@15878.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_39 = _T_2095_39; // @[NV_NVDLA_CSC_wl.scala 780:30:@15879.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_40 = _T_2095_40; // @[NV_NVDLA_CSC_wl.scala 780:30:@15880.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_41 = _T_2095_41; // @[NV_NVDLA_CSC_wl.scala 780:30:@15881.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_42 = _T_2095_42; // @[NV_NVDLA_CSC_wl.scala 780:30:@15882.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_43 = _T_2095_43; // @[NV_NVDLA_CSC_wl.scala 780:30:@15883.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_44 = _T_2095_44; // @[NV_NVDLA_CSC_wl.scala 780:30:@15884.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_45 = _T_2095_45; // @[NV_NVDLA_CSC_wl.scala 780:30:@15885.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_46 = _T_2095_46; // @[NV_NVDLA_CSC_wl.scala 780:30:@15886.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_47 = _T_2095_47; // @[NV_NVDLA_CSC_wl.scala 780:30:@15887.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_48 = _T_2095_48; // @[NV_NVDLA_CSC_wl.scala 780:30:@15888.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_49 = _T_2095_49; // @[NV_NVDLA_CSC_wl.scala 780:30:@15889.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_50 = _T_2095_50; // @[NV_NVDLA_CSC_wl.scala 780:30:@15890.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_51 = _T_2095_51; // @[NV_NVDLA_CSC_wl.scala 780:30:@15891.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_52 = _T_2095_52; // @[NV_NVDLA_CSC_wl.scala 780:30:@15892.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_53 = _T_2095_53; // @[NV_NVDLA_CSC_wl.scala 780:30:@15893.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_54 = _T_2095_54; // @[NV_NVDLA_CSC_wl.scala 780:30:@15894.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_55 = _T_2095_55; // @[NV_NVDLA_CSC_wl.scala 780:30:@15895.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_56 = _T_2095_56; // @[NV_NVDLA_CSC_wl.scala 780:30:@15896.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_57 = _T_2095_57; // @[NV_NVDLA_CSC_wl.scala 780:30:@15897.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_58 = _T_2095_58; // @[NV_NVDLA_CSC_wl.scala 780:30:@15898.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_59 = _T_2095_59; // @[NV_NVDLA_CSC_wl.scala 780:30:@15899.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_60 = _T_2095_60; // @[NV_NVDLA_CSC_wl.scala 780:30:@15900.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_61 = _T_2095_61; // @[NV_NVDLA_CSC_wl.scala 780:30:@15901.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_62 = _T_2095_62; // @[NV_NVDLA_CSC_wl.scala 780:30:@15902.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_data_63 = _T_2095_63; // @[NV_NVDLA_CSC_wl.scala 780:30:@15903.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_0 = _T_2362[0]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15970.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_1 = _T_2362[1]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15971.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_2 = _T_2362[2]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15972.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_3 = _T_2362[3]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15973.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_4 = _T_2362[4]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15974.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_5 = _T_2362[5]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15975.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_6 = _T_2362[6]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15976.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_7 = _T_2362[7]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15977.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_8 = _T_2362[8]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15978.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_9 = _T_2362[9]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15979.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_10 = _T_2362[10]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15980.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_11 = _T_2362[11]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15981.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_12 = _T_2362[12]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15982.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_13 = _T_2362[13]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15983.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_14 = _T_2362[14]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15984.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_15 = _T_2362[15]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15985.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_16 = _T_2362[16]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15986.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_17 = _T_2362[17]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15987.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_18 = _T_2362[18]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15988.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_19 = _T_2362[19]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15989.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_20 = _T_2362[20]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15990.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_21 = _T_2362[21]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15991.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_22 = _T_2362[22]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15992.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_23 = _T_2362[23]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15993.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_24 = _T_2362[24]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15994.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_25 = _T_2362[25]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15995.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_26 = _T_2362[26]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15996.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_27 = _T_2362[27]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15997.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_28 = _T_2362[28]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15998.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_29 = _T_2362[29]; // @[NV_NVDLA_CSC_wl.scala 784:29:@15999.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_30 = _T_2362[30]; // @[NV_NVDLA_CSC_wl.scala 784:29:@16000.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_bits_sel_31 = _T_2362[31]; // @[NV_NVDLA_CSC_wl.scala 784:29:@16001.4]
  assign NV_NVDLA_CSC_WL_dec_io_input_mask_en = _T_2938; // @[NV_NVDLA_CSC_wl.scala 782:28:@15968.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_698 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_715 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_722 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_729 = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_736 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_739 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_742 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1692 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_1712 = _RAND_8[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_798 = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_863 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_867 = _RAND_11[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_871 = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_877 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_882 = _RAND_14[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_893 = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_896 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_920 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_923 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1003 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1006 = _RAND_20[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1041 = _RAND_21[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1044 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1047 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1050 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1053 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1056 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1059 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1062 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1081 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1084 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1087 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1090 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_1093 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1096 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_1101 = _RAND_35[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_1104 = _RAND_36[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_1107 = _RAND_37[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_1110 = _RAND_38[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_1113 = _RAND_39[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1116 = _RAND_40[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {10{`RANDOM}};
  _T_1156 = _RAND_41[318:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {16{`RANDOM}};
  _T_1163 = _RAND_42[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {16{`RANDOM}};
  _T_1193 = _RAND_43[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1223 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1226 = _RAND_45[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1229 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1232 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1235 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1238 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1241 = _RAND_50[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1244 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1247 = _RAND_52[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  _T_1447 = _RAND_53[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1537 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1540 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1563 = _RAND_56[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1566 = _RAND_57[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1605 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1608 = _RAND_59[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1631 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1634 = _RAND_61[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1637 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1640 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1643 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1646 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1649 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1652 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1655 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1658 = _RAND_69[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1661 = _RAND_70[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1677 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1680 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1683 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1686 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1689 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {2{`RANDOM}};
  _T_1697 = _RAND_76[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {2{`RANDOM}};
  _T_1700 = _RAND_77[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {2{`RANDOM}};
  _T_1703 = _RAND_78[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {2{`RANDOM}};
  _T_1706 = _RAND_79[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {2{`RANDOM}};
  _T_1709 = _RAND_80[35:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1717 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1720 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1723 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1726 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1729 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1732 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {2{`RANDOM}};
  _T_1737 = _RAND_87[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {2{`RANDOM}};
  _T_1740 = _RAND_88[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {2{`RANDOM}};
  _T_1743 = _RAND_89[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {2{`RANDOM}};
  _T_1746 = _RAND_90[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {2{`RANDOM}};
  _T_1749 = _RAND_91[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {2{`RANDOM}};
  _T_1752 = _RAND_92[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1762 = _RAND_93[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1765 = _RAND_94[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {16{`RANDOM}};
  _T_1786 = _RAND_95[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {16{`RANDOM}};
  _T_1788 = _RAND_96[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_2095_0 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_2095_1 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_2095_2 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_2095_3 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_2095_4 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_2095_5 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_2095_6 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_2095_7 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_2095_8 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_2095_9 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_2095_10 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_2095_11 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_2095_12 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_2095_13 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_2095_14 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_2095_15 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_2095_16 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_2095_17 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_2095_18 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_2095_19 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_2095_20 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_2095_21 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_2095_22 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_2095_23 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_2095_24 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_2095_25 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_2095_26 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_2095_27 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_2095_28 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_2095_29 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_2095_30 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_2095_31 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_2095_32 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_2095_33 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_2095_34 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_2095_35 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_2095_36 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_2095_37 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_2095_38 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_2095_39 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_2095_40 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_2095_41 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_2095_42 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_2095_43 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_2095_44 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_2095_45 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_2095_46 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_2095_47 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2095_48 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2095_49 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_2095_50 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_2095_51 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_2095_52 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_2095_53 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_2095_54 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_2095_55 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_2095_56 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_2095_57 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_2095_58 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_2095_59 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_2095_60 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_2095_61 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_2095_62 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_2095_63 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_2359 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_2362 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_2472 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_2739_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_2739_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_2739_2 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_2739_3 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_2739_4 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_2739_5 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_2739_6 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_2739_7 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_2739_8 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_2739_9 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_2739_10 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_2739_11 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_2739_12 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_2739_13 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_2739_14 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_2739_15 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_2739_16 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_2739_17 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_2739_18 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_2739_19 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_2739_20 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_2739_21 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_2739_22 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_2739_23 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_2739_24 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_2739_25 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_2739_26 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_2739_27 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_2739_28 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_2739_29 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_2739_30 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_2739_31 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_2739_32 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_2739_33 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_2739_34 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_2739_35 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_2739_36 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_2739_37 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_2739_38 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_2739_39 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_2739_40 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_2739_41 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_2739_42 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_2739_43 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_2739_44 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_2739_45 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_2739_46 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_2739_47 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_2739_48 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_2739_49 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_2739_50 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_2739_51 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_2739_52 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_2739_53 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_2739_54 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_2739_55 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_2739_56 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_2739_57 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_2739_58 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_2739_59 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_2739_60 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_2739_61 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_2739_62 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_2739_63 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_2938 = _RAND_228[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3157 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3160 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3427_0 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3427_1 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3427_2 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3427_3 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3427_4 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3427_5 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3427_6 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3427_7 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3427_8 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3427_9 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3427_10 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3427_11 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3427_12 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3427_13 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3427_14 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3427_15 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3427_16 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3427_17 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3427_18 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3427_19 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3427_20 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3427_21 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3427_22 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3427_23 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3427_24 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3427_25 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3427_26 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3427_27 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3427_28 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3427_29 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3427_30 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3427_31 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3427_32 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3427_33 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3427_34 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3427_35 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3427_36 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3427_37 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3427_38 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3427_39 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3427_40 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3427_41 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3427_42 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3427_43 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3427_44 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3427_45 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3427_46 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3427_47 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3427_48 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3427_49 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3427_50 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_3427_51 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_3427_52 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_3427_53 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_3427_54 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_3427_55 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_3427_56 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_3427_57 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_3427_58 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_3427_59 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_3427_60 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_3427_61 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_3427_62 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_3427_63 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_3890_0 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_3890_1 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_3890_2 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_3890_3 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_3890_4 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_3890_5 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_3890_6 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_3890_7 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_3890_8 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_3890_9 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_3890_10 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_3890_11 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_3890_12 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_3890_13 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_3890_14 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_3890_15 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_3890_16 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_3890_17 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_3890_18 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_3890_19 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_3890_20 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_3890_21 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_3890_22 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_3890_23 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_3890_24 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_3890_25 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_3890_26 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_3890_27 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_3890_28 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_3890_29 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_3890_30 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_3890_31 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_3890_32 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_3890_33 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_3890_34 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_3890_35 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_3890_36 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_3890_37 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_3890_38 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_3890_39 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_3890_40 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_3890_41 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_3890_42 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_3890_43 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_3890_44 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_3890_45 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_3890_46 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_3890_47 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_3890_48 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_3890_49 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_3890_50 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_3890_51 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_3890_52 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_3890_53 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_3890_54 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_3890_55 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_3890_56 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_3890_57 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_3890_58 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_3890_59 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_3890_60 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_3890_61 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_3890_62 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_3890_63 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4161_0 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4161_1 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4161_2 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4161_3 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4161_4 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4161_5 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4161_6 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4161_7 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4161_8 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4161_9 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4161_10 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4161_11 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4161_12 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4161_13 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4161_14 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4161_15 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4288_0 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4288_1 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4288_2 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4288_3 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4288_4 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4288_5 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4288_6 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4288_7 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4288_8 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4288_9 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4288_10 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4288_11 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4288_12 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4288_13 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4288_14 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4288_15 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4344_0 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4344_1 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4344_2 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4344_3 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4344_4 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4344_5 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4344_6 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4344_7 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4344_8 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4344_9 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4344_10 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4344_11 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4344_12 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4344_13 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4344_14 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4344_15 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4344_16 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4344_17 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4344_18 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4344_19 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4344_20 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4344_21 = _RAND_412[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4344_22 = _RAND_413[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4344_23 = _RAND_414[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4344_24 = _RAND_415[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4344_25 = _RAND_416[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_4344_26 = _RAND_417[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_4344_27 = _RAND_418[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_4344_28 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_4344_29 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_4344_30 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_4344_31 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_4344_32 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_4344_33 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_4344_34 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_4344_35 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_4344_36 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_4344_37 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_4344_38 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_4344_39 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_4344_40 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_4344_41 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_4344_42 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_4344_43 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_4344_44 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_4344_45 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_4344_46 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_4344_47 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_4344_48 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_4344_49 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_4344_50 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_4344_51 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_4344_52 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_4344_53 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_4344_54 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_4344_55 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_4344_56 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_4344_57 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_4344_58 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_4344_59 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_4344_60 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_4344_61 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_4344_62 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_4344_63 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_4414_0 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_4414_1 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_4414_2 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_4414_3 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_4414_4 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_4414_5 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_4414_6 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_4414_7 = _RAND_462[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_4414_8 = _RAND_463[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_4414_9 = _RAND_464[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_4414_10 = _RAND_465[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_4414_11 = _RAND_466[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_4414_12 = _RAND_467[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_4414_13 = _RAND_468[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_4414_14 = _RAND_469[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_4414_15 = _RAND_470[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_4414_16 = _RAND_471[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_4414_17 = _RAND_472[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_4414_18 = _RAND_473[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_4414_19 = _RAND_474[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_4414_20 = _RAND_475[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_4414_21 = _RAND_476[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_4414_22 = _RAND_477[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_4414_23 = _RAND_478[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_4414_24 = _RAND_479[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_4414_25 = _RAND_480[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_4414_26 = _RAND_481[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_4414_27 = _RAND_482[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_4414_28 = _RAND_483[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_4414_29 = _RAND_484[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_4414_30 = _RAND_485[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_4414_31 = _RAND_486[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_4414_32 = _RAND_487[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_4414_33 = _RAND_488[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_4414_34 = _RAND_489[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_4414_35 = _RAND_490[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_4414_36 = _RAND_491[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_4414_37 = _RAND_492[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_4414_38 = _RAND_493[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_4414_39 = _RAND_494[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_4414_40 = _RAND_495[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_4414_41 = _RAND_496[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_4414_42 = _RAND_497[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_4414_43 = _RAND_498[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_4414_44 = _RAND_499[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_4414_45 = _RAND_500[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_4414_46 = _RAND_501[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_4414_47 = _RAND_502[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_4414_48 = _RAND_503[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_4414_49 = _RAND_504[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_4414_50 = _RAND_505[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_4414_51 = _RAND_506[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_4414_52 = _RAND_507[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_4414_53 = _RAND_508[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_4414_54 = _RAND_509[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_4414_55 = _RAND_510[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_4414_56 = _RAND_511[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_4414_57 = _RAND_512[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_4414_58 = _RAND_513[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_4414_59 = _RAND_514[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_4414_60 = _RAND_515[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_4414_61 = _RAND_516[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_4414_62 = _RAND_517[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_4414_63 = _RAND_518[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_698 <= 1'h0;
    end else begin
      _T_698 <= _T_704;
    end
    if (reset) begin
      _T_715 <= 5'h0;
    end else begin
      if (_T_743) begin
        _T_715 <= _T_750;
      end
    end
    if (reset) begin
      _T_722 <= 5'h0;
    end else begin
      if (_T_743) begin
        _T_722 <= _T_753;
      end
    end
    if (reset) begin
      _T_729 <= 15'h0;
    end else begin
      if (_T_757) begin
        _T_729 <= _T_758;
      end
    end
    if (reset) begin
      _T_736 <= 9'h0;
    end else begin
      if (_T_757) begin
        if (_T_742) begin
          _T_736 <= _T_759;
        end else begin
          _T_736 <= 9'h0;
        end
      end
    end
    if (reset) begin
      _T_739 <= 3'h1;
    end else begin
      if (_T_743) begin
        _T_739 <= _T_756;
      end
    end
    if (reset) begin
      _T_742 <= 1'h0;
    end else begin
      if (_T_743) begin
        _T_742 <= io_reg2dp_weight_format;
      end
    end
    if (reset) begin
      _T_1692 <= 1'h0;
    end else begin
      _T_1692 <= _T_1689;
    end
    if (reset) begin
      _T_1712 <= 36'h0;
    end else begin
      if (_T_1689) begin
        _T_1712 <= _T_1709;
      end
    end
    if (reset) begin
      _T_863 <= 1'h0;
    end else begin
      _T_863 <= _T_858;
    end
    if (reset) begin
      _T_867 <= 15'h0;
    end else begin
      if (_T_858) begin
        if (io_sg2wl_reuse_rls) begin
          _T_867 <= _T_729;
        end else begin
          _T_867 <= _T_1755;
        end
      end
    end
    if (reset) begin
      _T_871 <= 9'h0;
    end else begin
      if (_T_858) begin
        if (io_sg2wl_reuse_rls) begin
          _T_871 <= _T_736;
        end else begin
          _T_871 <= _T_1754;
        end
      end
    end
    if (reset) begin
      _T_877 <= 1'h0;
    end else begin
      _T_877 <= io_sg2wl_pd_valid;
    end
    if (reset) begin
      _T_882 <= 18'h0;
    end else begin
      if (io_sg2wl_pd_valid) begin
        _T_882 <= {{17'd0}, _T_879};
      end
    end
    if (reset) begin
      _T_893 <= 5'h0;
    end else begin
      if (_T_913) begin
        if (_T_743) begin
          _T_893 <= 5'h0;
        end else begin
          if (_T_905) begin
            _T_893 <= 5'h0;
          end else begin
            _T_893 <= _T_899;
          end
        end
      end
    end
    if (reset) begin
      _T_896 <= 1'h0;
    end else begin
      if (_T_877) begin
        _T_896 <= 1'h1;
      end else begin
        if (_T_909) begin
          _T_896 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_920 <= 11'h0;
    end else begin
      if (_T_972) begin
        if (_T_743) begin
          _T_920 <= 11'h0;
        end else begin
          if (_T_938) begin
            _T_920 <= _T_923;
          end else begin
            _T_920 <= _T_934;
          end
        end
      end
    end
    if (reset) begin
      _T_923 <= 11'h0;
    end else begin
      if (_T_976) begin
        if (_T_743) begin
          _T_923 <= 11'h0;
        end else begin
          if (!(_T_938)) begin
            _T_923 <= _T_934;
          end
        end
      end
    end
    if (reset) begin
      _T_1003 <= 1'h0;
    end else begin
      if (_T_1008) begin
        _T_1003 <= 1'h0;
      end else begin
        if (_T_1010) begin
          _T_1003 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1006 <= 9'h0;
    end else begin
      if (_T_1029) begin
        if (_T_743) begin
          _T_1006 <= 9'h0;
        end else begin
          if (_T_1018) begin
            _T_1006 <= 9'h0;
          end else begin
            _T_1006 <= _T_1016;
          end
        end
      end
    end
    if (reset) begin
      _T_1041 <= 7'h0;
    end else begin
      if (_T_912) begin
        _T_1041 <= _T_883;
      end
    end
    if (reset) begin
      _T_1044 <= 8'h0;
    end else begin
      if (_T_912) begin
        _T_1044 <= _T_917;
      end
    end
    if (reset) begin
      _T_1047 <= 9'h0;
    end else begin
      if (_T_1064) begin
        if (_T_1031) begin
          _T_1047 <= _T_1006;
        end else begin
          _T_1047 <= _T_1016;
        end
      end
    end
    if (reset) begin
      _T_1050 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1050 <= _T_905;
      end
    end
    if (reset) begin
      _T_1053 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1053 <= _T_1010;
      end
    end
    if (reset) begin
      _T_1056 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1056 <= _T_1007;
      end
    end
    if (reset) begin
      _T_1059 <= 1'h0;
    end else begin
      if (_T_912) begin
        _T_1059 <= _T_1067;
      end
    end
    if (reset) begin
      _T_1062 <= 2'h0;
    end else begin
      if (_T_912) begin
        _T_1062 <= _T_885;
      end
    end
    if (reset) begin
      _T_1081 <= 1'h0;
    end else begin
      _T_1081 <= _T_896;
    end
    if (reset) begin
      _T_1084 <= 1'h0;
    end else begin
      _T_1084 <= _T_1081;
    end
    if (reset) begin
      _T_1087 <= 1'h0;
    end else begin
      _T_1087 <= _T_1084;
    end
    if (reset) begin
      _T_1090 <= 1'h0;
    end else begin
      _T_1090 <= _T_1087;
    end
    if (reset) begin
      _T_1093 <= 1'h0;
    end else begin
      _T_1093 <= _T_1090;
    end
    if (reset) begin
      _T_1096 <= 1'h0;
    end else begin
      _T_1096 <= _T_1093;
    end
    if (reset) begin
      _T_1101 <= 31'h0;
    end else begin
      if (_T_896) begin
        _T_1101 <= _T_1076;
      end
    end
    if (reset) begin
      _T_1104 <= 31'h0;
    end else begin
      if (_T_1081) begin
        _T_1104 <= _T_1101;
      end
    end
    if (reset) begin
      _T_1107 <= 31'h0;
    end else begin
      if (_T_1084) begin
        _T_1107 <= _T_1104;
      end
    end
    if (reset) begin
      _T_1110 <= 31'h0;
    end else begin
      if (_T_1087) begin
        _T_1110 <= _T_1107;
      end
    end
    if (reset) begin
      _T_1113 <= 31'h0;
    end else begin
      if (_T_1090) begin
        _T_1113 <= _T_1110;
      end
    end
    if (reset) begin
      _T_1116 <= 31'h0;
    end else begin
      if (_T_1093) begin
        _T_1116 <= _T_1113;
      end
    end
    if (reset) begin
      _T_1156 <= 319'h0;
    end else begin
      if (_T_1096) begin
        _T_1156 <= _T_1186;
      end
    end
    if (reset) begin
      _T_1163 <= 512'h0;
    end else begin
      if (_T_1149) begin
        if (_T_743) begin
          _T_1163 <= 512'h0;
        end else begin
          if (_T_1138) begin
            _T_1163 <= _T_1193;
          end else begin
            _T_1163 <= _T_1199;
          end
        end
      end
    end
    if (reset) begin
      _T_1193 <= 512'h0;
    end else begin
      if (_T_1147) begin
        if (_T_743) begin
          _T_1193 <= 512'h0;
        end else begin
          if (!(_T_1138)) begin
            _T_1193 <= _T_1199;
          end
        end
      end
    end
    if (reset) begin
      _T_1223 <= 1'h0;
    end else begin
      _T_1223 <= _T_1096;
    end
    if (reset) begin
      _T_1226 <= 7'h0;
    end else begin
      if (_T_1096) begin
        _T_1226 <= _T_1117;
      end
    end
    if (reset) begin
      _T_1229 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1229 <= _T_1120;
      end
    end
    if (reset) begin
      _T_1232 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1232 <= _T_1121;
      end
    end
    if (reset) begin
      _T_1235 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1235 <= _T_1122;
      end
    end
    if (reset) begin
      _T_1238 <= 1'h0;
    end else begin
      if (_T_1096) begin
        _T_1238 <= _T_1123;
      end
    end
    if (reset) begin
      _T_1241 <= 9'h0;
    end else begin
      if (_T_1096) begin
        _T_1241 <= _T_1119;
      end
    end
    if (reset) begin
      _T_1244 <= 2'h0;
    end else begin
      if (_T_1096) begin
        _T_1244 <= _T_1124;
      end
    end
    if (reset) begin
      _T_1247 <= 7'h0;
    end else begin
      if (_T_1096) begin
        _T_1247 <= {{1'd0}, _T_1220};
      end
    end
    if (reset) begin
      _T_1447 <= 64'h0;
    end else begin
      _T_1447 <= _GEN_60[63:0];
    end
    if (reset) begin
      _T_1537 <= 8'h0;
    end else begin
      _T_1537 <= _GEN_49[7:0];
    end
    if (reset) begin
      _T_1540 <= 8'h0;
    end else begin
      _T_1540 <= _GEN_50[7:0];
    end
    if (reset) begin
      _T_1563 <= 13'h0;
    end else begin
      if (_T_1591) begin
        if (_T_708) begin
          _T_1563 <= _T_1583;
        end else begin
          if (_T_1554) begin
            _T_1563 <= _T_1566;
          end else begin
            if (_T_1542) begin
              if (_T_1576) begin
                _T_1563 <= 13'h0;
              end else begin
                _T_1563 <= _T_1569;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1566 <= 13'h0;
    end else begin
      if (_T_1594) begin
        if (_T_708) begin
          _T_1566 <= _T_1583;
        end else begin
          if (!(_T_1554)) begin
            if (_T_1542) begin
              if (_T_1576) begin
                _T_1566 <= 13'h0;
              end else begin
                _T_1566 <= _T_1569;
              end
            end else begin
              _T_1566 <= _T_1563;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1605 <= 1'h0;
    end else begin
      if (_T_1609) begin
        _T_1605 <= 1'h0;
      end else begin
        if (_T_1232) begin
          _T_1605 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1608 <= 15'h0;
    end else begin
      if (_T_1625) begin
        if (_T_743) begin
          _T_1608 <= 15'h0;
        end else begin
          if (_T_1235) begin
            _T_1608 <= 15'h0;
          end else begin
            _T_1608 <= _T_1616;
          end
        end
      end
    end
    if (reset) begin
      _T_1631 <= 1'h0;
    end else begin
      _T_1631 <= _T_1542;
    end
    if (reset) begin
      _T_1634 <= 13'h0;
    end else begin
      _T_1634 <= _GEN_54[12:0];
    end
    if (reset) begin
      _T_1637 <= 1'h0;
    end else begin
      _T_1637 <= _T_1223;
    end
    if (reset) begin
      _T_1640 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1640 <= _T_1229;
      end
    end
    if (reset) begin
      _T_1643 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1643 <= _T_1232;
      end
    end
    if (reset) begin
      _T_1646 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1646 <= _T_1235;
      end
    end
    if (reset) begin
      _T_1649 <= 1'h0;
    end else begin
      if (_T_1223) begin
        _T_1649 <= _T_1238;
      end
    end
    if (reset) begin
      _T_1652 <= 8'h0;
    end else begin
      _T_1652 <= _GEN_59[7:0];
    end
    if (reset) begin
      _T_1655 <= 1'h0;
    end else begin
      _T_1655 <= _T_1534;
    end
    if (reset) begin
      _T_1658 <= 9'h0;
    end else begin
      if (_T_1223) begin
        _T_1658 <= _T_1241;
      end
    end
    if (reset) begin
      _T_1661 <= 15'h0;
    end else begin
      if (_T_1663) begin
        if (_T_1627) begin
          _T_1661 <= _T_1608;
        end else begin
          _T_1661 <= _T_1616;
        end
      end
    end
    if (reset) begin
      _T_1677 <= 1'h0;
    end else begin
      _T_1677 <= _T_1637;
    end
    if (reset) begin
      _T_1680 <= 1'h0;
    end else begin
      _T_1680 <= _T_1677;
    end
    if (reset) begin
      _T_1683 <= 1'h0;
    end else begin
      _T_1683 <= _T_1680;
    end
    if (reset) begin
      _T_1686 <= 1'h0;
    end else begin
      _T_1686 <= _T_1683;
    end
    if (reset) begin
      _T_1689 <= 1'h0;
    end else begin
      _T_1689 <= _T_1686;
    end
    if (reset) begin
      _T_1697 <= 36'h0;
    end else begin
      if (_T_1637) begin
        _T_1697 <= _T_1672;
      end
    end
    if (reset) begin
      _T_1700 <= 36'h0;
    end else begin
      if (_T_1677) begin
        _T_1700 <= _T_1697;
      end
    end
    if (reset) begin
      _T_1703 <= 36'h0;
    end else begin
      if (_T_1680) begin
        _T_1703 <= _T_1700;
      end
    end
    if (reset) begin
      _T_1706 <= 36'h0;
    end else begin
      if (_T_1683) begin
        _T_1706 <= _T_1703;
      end
    end
    if (reset) begin
      _T_1709 <= 36'h0;
    end else begin
      if (_T_1686) begin
        _T_1709 <= _T_1706;
      end
    end
    if (reset) begin
      _T_1717 <= 1'h0;
    end else begin
      _T_1717 <= _T_1655;
    end
    if (reset) begin
      _T_1720 <= 1'h0;
    end else begin
      _T_1720 <= _T_1717;
    end
    if (reset) begin
      _T_1723 <= 1'h0;
    end else begin
      _T_1723 <= _T_1720;
    end
    if (reset) begin
      _T_1726 <= 1'h0;
    end else begin
      _T_1726 <= _T_1723;
    end
    if (reset) begin
      _T_1729 <= 1'h0;
    end else begin
      _T_1729 <= _T_1726;
    end
    if (reset) begin
      _T_1732 <= 1'h0;
    end else begin
      _T_1732 <= _T_1729;
    end
    if (reset) begin
      _T_1737 <= 64'h0;
    end else begin
      if (_T_1655) begin
        _T_1737 <= _T_1447;
      end
    end
    if (reset) begin
      _T_1740 <= 64'h0;
    end else begin
      if (_T_1717) begin
        _T_1740 <= _T_1737;
      end
    end
    if (reset) begin
      _T_1743 <= 64'h0;
    end else begin
      if (_T_1720) begin
        _T_1743 <= _T_1740;
      end
    end
    if (reset) begin
      _T_1746 <= 64'h0;
    end else begin
      if (_T_1723) begin
        _T_1746 <= _T_1743;
      end
    end
    if (reset) begin
      _T_1749 <= 64'h0;
    end else begin
      if (_T_1726) begin
        _T_1749 <= _T_1746;
      end
    end
    if (reset) begin
      _T_1752 <= 64'h0;
    end else begin
      if (_T_1729) begin
        _T_1752 <= _T_1749;
      end
    end
    if (reset) begin
      _T_1762 <= 7'h0;
    end else begin
      if (_T_1782) begin
        _T_1762 <= _T_1781;
      end
    end
    if (reset) begin
      _T_1765 <= 7'h0;
    end else begin
      if (_T_1784) begin
        _T_1765 <= _T_1781;
      end
    end
    if (_T_1817) begin
      if (_T_743) begin
        _T_1786 <= 512'h0;
      end else begin
        if (_T_1810) begin
          _T_1786 <= _T_1788;
        end else begin
          if (io_sc2buf_wt_rd_data_valid) begin
            _T_1786 <= _T_1796;
          end else begin
            _T_1786 <= _T_1804;
          end
        end
      end
    end
    if (_T_1822) begin
      if (_T_743) begin
        _T_1788 <= 512'h0;
      end else begin
        if (!(_T_1810)) begin
          if (io_sc2buf_wt_rd_data_valid) begin
            _T_1788 <= _T_1796;
          end else begin
            _T_1788 <= _T_1804;
          end
        end
      end
    end
    if (reset) begin
      _T_2095_0 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_0 <= _T_2293;
      end
    end
    if (reset) begin
      _T_2095_1 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_1 <= _T_2294;
      end
    end
    if (reset) begin
      _T_2095_2 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_2 <= _T_2295;
      end
    end
    if (reset) begin
      _T_2095_3 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_3 <= _T_2296;
      end
    end
    if (reset) begin
      _T_2095_4 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_4 <= _T_2297;
      end
    end
    if (reset) begin
      _T_2095_5 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_5 <= _T_2298;
      end
    end
    if (reset) begin
      _T_2095_6 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_6 <= _T_2299;
      end
    end
    if (reset) begin
      _T_2095_7 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_7 <= _T_2300;
      end
    end
    if (reset) begin
      _T_2095_8 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_8 <= _T_2301;
      end
    end
    if (reset) begin
      _T_2095_9 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_9 <= _T_2302;
      end
    end
    if (reset) begin
      _T_2095_10 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_10 <= _T_2303;
      end
    end
    if (reset) begin
      _T_2095_11 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_11 <= _T_2304;
      end
    end
    if (reset) begin
      _T_2095_12 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_12 <= _T_2305;
      end
    end
    if (reset) begin
      _T_2095_13 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_13 <= _T_2306;
      end
    end
    if (reset) begin
      _T_2095_14 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_14 <= _T_2307;
      end
    end
    if (reset) begin
      _T_2095_15 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_15 <= _T_2308;
      end
    end
    if (reset) begin
      _T_2095_16 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_16 <= _T_2309;
      end
    end
    if (reset) begin
      _T_2095_17 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_17 <= _T_2310;
      end
    end
    if (reset) begin
      _T_2095_18 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_18 <= _T_2311;
      end
    end
    if (reset) begin
      _T_2095_19 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_19 <= _T_2312;
      end
    end
    if (reset) begin
      _T_2095_20 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_20 <= _T_2313;
      end
    end
    if (reset) begin
      _T_2095_21 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_21 <= _T_2314;
      end
    end
    if (reset) begin
      _T_2095_22 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_22 <= _T_2315;
      end
    end
    if (reset) begin
      _T_2095_23 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_23 <= _T_2316;
      end
    end
    if (reset) begin
      _T_2095_24 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_24 <= _T_2317;
      end
    end
    if (reset) begin
      _T_2095_25 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_25 <= _T_2318;
      end
    end
    if (reset) begin
      _T_2095_26 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_26 <= _T_2319;
      end
    end
    if (reset) begin
      _T_2095_27 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_27 <= _T_2320;
      end
    end
    if (reset) begin
      _T_2095_28 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_28 <= _T_2321;
      end
    end
    if (reset) begin
      _T_2095_29 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_29 <= _T_2322;
      end
    end
    if (reset) begin
      _T_2095_30 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_30 <= _T_2323;
      end
    end
    if (reset) begin
      _T_2095_31 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_31 <= _T_2324;
      end
    end
    if (reset) begin
      _T_2095_32 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_32 <= _T_2325;
      end
    end
    if (reset) begin
      _T_2095_33 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_33 <= _T_2326;
      end
    end
    if (reset) begin
      _T_2095_34 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_34 <= _T_2327;
      end
    end
    if (reset) begin
      _T_2095_35 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_35 <= _T_2328;
      end
    end
    if (reset) begin
      _T_2095_36 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_36 <= _T_2329;
      end
    end
    if (reset) begin
      _T_2095_37 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_37 <= _T_2330;
      end
    end
    if (reset) begin
      _T_2095_38 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_38 <= _T_2331;
      end
    end
    if (reset) begin
      _T_2095_39 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_39 <= _T_2332;
      end
    end
    if (reset) begin
      _T_2095_40 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_40 <= _T_2333;
      end
    end
    if (reset) begin
      _T_2095_41 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_41 <= _T_2334;
      end
    end
    if (reset) begin
      _T_2095_42 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_42 <= _T_2335;
      end
    end
    if (reset) begin
      _T_2095_43 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_43 <= _T_2336;
      end
    end
    if (reset) begin
      _T_2095_44 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_44 <= _T_2337;
      end
    end
    if (reset) begin
      _T_2095_45 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_45 <= _T_2338;
      end
    end
    if (reset) begin
      _T_2095_46 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_46 <= _T_2339;
      end
    end
    if (reset) begin
      _T_2095_47 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_47 <= _T_2340;
      end
    end
    if (reset) begin
      _T_2095_48 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_48 <= _T_2341;
      end
    end
    if (reset) begin
      _T_2095_49 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_49 <= _T_2342;
      end
    end
    if (reset) begin
      _T_2095_50 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_50 <= _T_2343;
      end
    end
    if (reset) begin
      _T_2095_51 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_51 <= _T_2344;
      end
    end
    if (reset) begin
      _T_2095_52 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_52 <= _T_2345;
      end
    end
    if (reset) begin
      _T_2095_53 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_53 <= _T_2346;
      end
    end
    if (reset) begin
      _T_2095_54 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_54 <= _T_2347;
      end
    end
    if (reset) begin
      _T_2095_55 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_55 <= _T_2348;
      end
    end
    if (reset) begin
      _T_2095_56 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_56 <= _T_2349;
      end
    end
    if (reset) begin
      _T_2095_57 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_57 <= _T_2350;
      end
    end
    if (reset) begin
      _T_2095_58 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_58 <= _T_2351;
      end
    end
    if (reset) begin
      _T_2095_59 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_59 <= _T_2352;
      end
    end
    if (reset) begin
      _T_2095_60 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_60 <= _T_2353;
      end
    end
    if (reset) begin
      _T_2095_61 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_61 <= _T_2354;
      end
    end
    if (reset) begin
      _T_2095_62 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_62 <= _T_2355;
      end
    end
    if (reset) begin
      _T_2095_63 <= 8'h0;
    end else begin
      if (_T_1692) begin
        _T_2095_63 <= _T_2356;
      end
    end
    if (reset) begin
      _T_2359 <= 1'h0;
    end else begin
      if (_T_1692) begin
        _T_2359 <= _T_1756;
      end
    end
    if (reset) begin
      _T_2362 <= 32'h1;
    end else begin
      if (_T_1692) begin
        if (_T_2359) begin
          _T_2362 <= 32'h1;
        end else begin
          _T_2362 <= _T_2366;
        end
      end
    end
    if (reset) begin
      _T_2472 <= 1'h0;
    end else begin
      _T_2472 <= _T_1692;
    end
    if (reset) begin
      _T_2739_0 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_0 <= _T_2939;
      end
    end
    if (reset) begin
      _T_2739_1 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_1 <= _T_2940;
      end
    end
    if (reset) begin
      _T_2739_2 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_2 <= _T_2941;
      end
    end
    if (reset) begin
      _T_2739_3 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_3 <= _T_2942;
      end
    end
    if (reset) begin
      _T_2739_4 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_4 <= _T_2943;
      end
    end
    if (reset) begin
      _T_2739_5 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_5 <= _T_2944;
      end
    end
    if (reset) begin
      _T_2739_6 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_6 <= _T_2945;
      end
    end
    if (reset) begin
      _T_2739_7 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_7 <= _T_2946;
      end
    end
    if (reset) begin
      _T_2739_8 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_8 <= _T_2947;
      end
    end
    if (reset) begin
      _T_2739_9 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_9 <= _T_2948;
      end
    end
    if (reset) begin
      _T_2739_10 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_10 <= _T_2949;
      end
    end
    if (reset) begin
      _T_2739_11 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_11 <= _T_2950;
      end
    end
    if (reset) begin
      _T_2739_12 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_12 <= _T_2951;
      end
    end
    if (reset) begin
      _T_2739_13 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_13 <= _T_2952;
      end
    end
    if (reset) begin
      _T_2739_14 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_14 <= _T_2953;
      end
    end
    if (reset) begin
      _T_2739_15 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_15 <= _T_2954;
      end
    end
    if (reset) begin
      _T_2739_16 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_16 <= _T_2955;
      end
    end
    if (reset) begin
      _T_2739_17 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_17 <= _T_2956;
      end
    end
    if (reset) begin
      _T_2739_18 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_18 <= _T_2957;
      end
    end
    if (reset) begin
      _T_2739_19 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_19 <= _T_2958;
      end
    end
    if (reset) begin
      _T_2739_20 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_20 <= _T_2959;
      end
    end
    if (reset) begin
      _T_2739_21 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_21 <= _T_2960;
      end
    end
    if (reset) begin
      _T_2739_22 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_22 <= _T_2961;
      end
    end
    if (reset) begin
      _T_2739_23 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_23 <= _T_2962;
      end
    end
    if (reset) begin
      _T_2739_24 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_24 <= _T_2963;
      end
    end
    if (reset) begin
      _T_2739_25 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_25 <= _T_2964;
      end
    end
    if (reset) begin
      _T_2739_26 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_26 <= _T_2965;
      end
    end
    if (reset) begin
      _T_2739_27 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_27 <= _T_2966;
      end
    end
    if (reset) begin
      _T_2739_28 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_28 <= _T_2967;
      end
    end
    if (reset) begin
      _T_2739_29 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_29 <= _T_2968;
      end
    end
    if (reset) begin
      _T_2739_30 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_30 <= _T_2969;
      end
    end
    if (reset) begin
      _T_2739_31 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_31 <= _T_2970;
      end
    end
    if (reset) begin
      _T_2739_32 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_32 <= _T_2971;
      end
    end
    if (reset) begin
      _T_2739_33 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_33 <= _T_2972;
      end
    end
    if (reset) begin
      _T_2739_34 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_34 <= _T_2973;
      end
    end
    if (reset) begin
      _T_2739_35 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_35 <= _T_2974;
      end
    end
    if (reset) begin
      _T_2739_36 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_36 <= _T_2975;
      end
    end
    if (reset) begin
      _T_2739_37 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_37 <= _T_2976;
      end
    end
    if (reset) begin
      _T_2739_38 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_38 <= _T_2977;
      end
    end
    if (reset) begin
      _T_2739_39 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_39 <= _T_2978;
      end
    end
    if (reset) begin
      _T_2739_40 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_40 <= _T_2979;
      end
    end
    if (reset) begin
      _T_2739_41 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_41 <= _T_2980;
      end
    end
    if (reset) begin
      _T_2739_42 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_42 <= _T_2981;
      end
    end
    if (reset) begin
      _T_2739_43 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_43 <= _T_2982;
      end
    end
    if (reset) begin
      _T_2739_44 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_44 <= _T_2983;
      end
    end
    if (reset) begin
      _T_2739_45 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_45 <= _T_2984;
      end
    end
    if (reset) begin
      _T_2739_46 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_46 <= _T_2985;
      end
    end
    if (reset) begin
      _T_2739_47 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_47 <= _T_2986;
      end
    end
    if (reset) begin
      _T_2739_48 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_48 <= _T_2987;
      end
    end
    if (reset) begin
      _T_2739_49 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_49 <= _T_2988;
      end
    end
    if (reset) begin
      _T_2739_50 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_50 <= _T_2989;
      end
    end
    if (reset) begin
      _T_2739_51 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_51 <= _T_2990;
      end
    end
    if (reset) begin
      _T_2739_52 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_52 <= _T_2991;
      end
    end
    if (reset) begin
      _T_2739_53 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_53 <= _T_2992;
      end
    end
    if (reset) begin
      _T_2739_54 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_54 <= _T_2993;
      end
    end
    if (reset) begin
      _T_2739_55 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_55 <= _T_2994;
      end
    end
    if (reset) begin
      _T_2739_56 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_56 <= _T_2995;
      end
    end
    if (reset) begin
      _T_2739_57 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_57 <= _T_2996;
      end
    end
    if (reset) begin
      _T_2739_58 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_58 <= _T_2997;
      end
    end
    if (reset) begin
      _T_2739_59 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_59 <= _T_2998;
      end
    end
    if (reset) begin
      _T_2739_60 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_60 <= _T_2999;
      end
    end
    if (reset) begin
      _T_2739_61 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_61 <= _T_3000;
      end
    end
    if (reset) begin
      _T_2739_62 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_62 <= _T_3001;
      end
    end
    if (reset) begin
      _T_2739_63 <= 1'h0;
    end else begin
      if (_T_1732) begin
        _T_2739_63 <= _T_3002;
      end
    end
    if (reset) begin
      _T_2938 <= 10'h0;
    end else begin
      if (_T_1732) begin
        _T_2938 <= 10'h3ff;
      end else begin
        _T_2938 <= 10'h0;
      end
    end
    if (reset) begin
      _T_3157 <= 1'h0;
    end else begin
      _T_3157 <= _T_3152;
    end
    if (reset) begin
      _T_3160 <= 1'h0;
    end else begin
      _T_3160 <= _T_3154;
    end
    if (reset) begin
      _T_3427_0 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_0 <= _T_4482;
      end
    end
    if (reset) begin
      _T_3427_1 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_1 <= _T_4484;
      end
    end
    if (reset) begin
      _T_3427_2 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_2 <= _T_4486;
      end
    end
    if (reset) begin
      _T_3427_3 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_3 <= _T_4488;
      end
    end
    if (reset) begin
      _T_3427_4 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_4 <= _T_4490;
      end
    end
    if (reset) begin
      _T_3427_5 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_5 <= _T_4492;
      end
    end
    if (reset) begin
      _T_3427_6 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_6 <= _T_4494;
      end
    end
    if (reset) begin
      _T_3427_7 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_7 <= _T_4496;
      end
    end
    if (reset) begin
      _T_3427_8 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_8 <= _T_4498;
      end
    end
    if (reset) begin
      _T_3427_9 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_9 <= _T_4500;
      end
    end
    if (reset) begin
      _T_3427_10 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_10 <= _T_4502;
      end
    end
    if (reset) begin
      _T_3427_11 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_11 <= _T_4504;
      end
    end
    if (reset) begin
      _T_3427_12 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_12 <= _T_4506;
      end
    end
    if (reset) begin
      _T_3427_13 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_13 <= _T_4508;
      end
    end
    if (reset) begin
      _T_3427_14 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_14 <= _T_4510;
      end
    end
    if (reset) begin
      _T_3427_15 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_15 <= _T_4512;
      end
    end
    if (reset) begin
      _T_3427_16 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_16 <= _T_4514;
      end
    end
    if (reset) begin
      _T_3427_17 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_17 <= _T_4516;
      end
    end
    if (reset) begin
      _T_3427_18 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_18 <= _T_4518;
      end
    end
    if (reset) begin
      _T_3427_19 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_19 <= _T_4520;
      end
    end
    if (reset) begin
      _T_3427_20 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_20 <= _T_4522;
      end
    end
    if (reset) begin
      _T_3427_21 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_21 <= _T_4524;
      end
    end
    if (reset) begin
      _T_3427_22 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_22 <= _T_4526;
      end
    end
    if (reset) begin
      _T_3427_23 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_23 <= _T_4528;
      end
    end
    if (reset) begin
      _T_3427_24 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_24 <= _T_4530;
      end
    end
    if (reset) begin
      _T_3427_25 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_25 <= _T_4532;
      end
    end
    if (reset) begin
      _T_3427_26 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_26 <= _T_4534;
      end
    end
    if (reset) begin
      _T_3427_27 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_27 <= _T_4536;
      end
    end
    if (reset) begin
      _T_3427_28 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_28 <= _T_4538;
      end
    end
    if (reset) begin
      _T_3427_29 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_29 <= _T_4540;
      end
    end
    if (reset) begin
      _T_3427_30 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_30 <= _T_4542;
      end
    end
    if (reset) begin
      _T_3427_31 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_31 <= _T_4544;
      end
    end
    if (reset) begin
      _T_3427_32 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_32 <= _T_4546;
      end
    end
    if (reset) begin
      _T_3427_33 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_33 <= _T_4548;
      end
    end
    if (reset) begin
      _T_3427_34 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_34 <= _T_4550;
      end
    end
    if (reset) begin
      _T_3427_35 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_35 <= _T_4552;
      end
    end
    if (reset) begin
      _T_3427_36 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_36 <= _T_4554;
      end
    end
    if (reset) begin
      _T_3427_37 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_37 <= _T_4556;
      end
    end
    if (reset) begin
      _T_3427_38 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_38 <= _T_4558;
      end
    end
    if (reset) begin
      _T_3427_39 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_39 <= _T_4560;
      end
    end
    if (reset) begin
      _T_3427_40 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_40 <= _T_4562;
      end
    end
    if (reset) begin
      _T_3427_41 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_41 <= _T_4564;
      end
    end
    if (reset) begin
      _T_3427_42 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_42 <= _T_4566;
      end
    end
    if (reset) begin
      _T_3427_43 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_43 <= _T_4568;
      end
    end
    if (reset) begin
      _T_3427_44 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_44 <= _T_4570;
      end
    end
    if (reset) begin
      _T_3427_45 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_45 <= _T_4572;
      end
    end
    if (reset) begin
      _T_3427_46 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_46 <= _T_4574;
      end
    end
    if (reset) begin
      _T_3427_47 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_47 <= _T_4576;
      end
    end
    if (reset) begin
      _T_3427_48 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_48 <= _T_4578;
      end
    end
    if (reset) begin
      _T_3427_49 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_49 <= _T_4580;
      end
    end
    if (reset) begin
      _T_3427_50 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_50 <= _T_4582;
      end
    end
    if (reset) begin
      _T_3427_51 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_51 <= _T_4584;
      end
    end
    if (reset) begin
      _T_3427_52 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_52 <= _T_4586;
      end
    end
    if (reset) begin
      _T_3427_53 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_53 <= _T_4588;
      end
    end
    if (reset) begin
      _T_3427_54 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_54 <= _T_4590;
      end
    end
    if (reset) begin
      _T_3427_55 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_55 <= _T_4592;
      end
    end
    if (reset) begin
      _T_3427_56 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_56 <= _T_4594;
      end
    end
    if (reset) begin
      _T_3427_57 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_57 <= _T_4596;
      end
    end
    if (reset) begin
      _T_3427_58 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_58 <= _T_4598;
      end
    end
    if (reset) begin
      _T_3427_59 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_59 <= _T_4600;
      end
    end
    if (reset) begin
      _T_3427_60 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_60 <= _T_4602;
      end
    end
    if (reset) begin
      _T_3427_61 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_61 <= _T_4604;
      end
    end
    if (reset) begin
      _T_3427_62 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_62 <= _T_4606;
      end
    end
    if (reset) begin
      _T_3427_63 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_3427_63 <= _T_4608;
      end
    end
    if (reset) begin
      _T_3890_0 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_0 <= _T_4680;
      end
    end
    if (reset) begin
      _T_3890_1 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_1 <= _T_4682;
      end
    end
    if (reset) begin
      _T_3890_2 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_2 <= _T_4684;
      end
    end
    if (reset) begin
      _T_3890_3 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_3 <= _T_4686;
      end
    end
    if (reset) begin
      _T_3890_4 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_4 <= _T_4688;
      end
    end
    if (reset) begin
      _T_3890_5 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_5 <= _T_4690;
      end
    end
    if (reset) begin
      _T_3890_6 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_6 <= _T_4692;
      end
    end
    if (reset) begin
      _T_3890_7 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_7 <= _T_4694;
      end
    end
    if (reset) begin
      _T_3890_8 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_8 <= _T_4696;
      end
    end
    if (reset) begin
      _T_3890_9 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_9 <= _T_4698;
      end
    end
    if (reset) begin
      _T_3890_10 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_10 <= _T_4700;
      end
    end
    if (reset) begin
      _T_3890_11 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_11 <= _T_4702;
      end
    end
    if (reset) begin
      _T_3890_12 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_12 <= _T_4704;
      end
    end
    if (reset) begin
      _T_3890_13 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_13 <= _T_4706;
      end
    end
    if (reset) begin
      _T_3890_14 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_14 <= _T_4708;
      end
    end
    if (reset) begin
      _T_3890_15 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_15 <= _T_4710;
      end
    end
    if (reset) begin
      _T_3890_16 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_16 <= _T_4712;
      end
    end
    if (reset) begin
      _T_3890_17 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_17 <= _T_4714;
      end
    end
    if (reset) begin
      _T_3890_18 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_18 <= _T_4716;
      end
    end
    if (reset) begin
      _T_3890_19 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_19 <= _T_4718;
      end
    end
    if (reset) begin
      _T_3890_20 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_20 <= _T_4720;
      end
    end
    if (reset) begin
      _T_3890_21 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_21 <= _T_4722;
      end
    end
    if (reset) begin
      _T_3890_22 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_22 <= _T_4724;
      end
    end
    if (reset) begin
      _T_3890_23 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_23 <= _T_4726;
      end
    end
    if (reset) begin
      _T_3890_24 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_24 <= _T_4728;
      end
    end
    if (reset) begin
      _T_3890_25 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_25 <= _T_4730;
      end
    end
    if (reset) begin
      _T_3890_26 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_26 <= _T_4732;
      end
    end
    if (reset) begin
      _T_3890_27 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_27 <= _T_4734;
      end
    end
    if (reset) begin
      _T_3890_28 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_28 <= _T_4736;
      end
    end
    if (reset) begin
      _T_3890_29 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_29 <= _T_4738;
      end
    end
    if (reset) begin
      _T_3890_30 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_30 <= _T_4740;
      end
    end
    if (reset) begin
      _T_3890_31 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_31 <= _T_4742;
      end
    end
    if (reset) begin
      _T_3890_32 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_32 <= _T_4744;
      end
    end
    if (reset) begin
      _T_3890_33 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_33 <= _T_4746;
      end
    end
    if (reset) begin
      _T_3890_34 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_34 <= _T_4748;
      end
    end
    if (reset) begin
      _T_3890_35 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_35 <= _T_4750;
      end
    end
    if (reset) begin
      _T_3890_36 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_36 <= _T_4752;
      end
    end
    if (reset) begin
      _T_3890_37 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_37 <= _T_4754;
      end
    end
    if (reset) begin
      _T_3890_38 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_38 <= _T_4756;
      end
    end
    if (reset) begin
      _T_3890_39 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_39 <= _T_4758;
      end
    end
    if (reset) begin
      _T_3890_40 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_40 <= _T_4760;
      end
    end
    if (reset) begin
      _T_3890_41 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_41 <= _T_4762;
      end
    end
    if (reset) begin
      _T_3890_42 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_42 <= _T_4764;
      end
    end
    if (reset) begin
      _T_3890_43 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_43 <= _T_4766;
      end
    end
    if (reset) begin
      _T_3890_44 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_44 <= _T_4768;
      end
    end
    if (reset) begin
      _T_3890_45 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_45 <= _T_4770;
      end
    end
    if (reset) begin
      _T_3890_46 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_46 <= _T_4772;
      end
    end
    if (reset) begin
      _T_3890_47 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_47 <= _T_4774;
      end
    end
    if (reset) begin
      _T_3890_48 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_48 <= _T_4776;
      end
    end
    if (reset) begin
      _T_3890_49 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_49 <= _T_4778;
      end
    end
    if (reset) begin
      _T_3890_50 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_50 <= _T_4780;
      end
    end
    if (reset) begin
      _T_3890_51 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_51 <= _T_4782;
      end
    end
    if (reset) begin
      _T_3890_52 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_52 <= _T_4784;
      end
    end
    if (reset) begin
      _T_3890_53 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_53 <= _T_4786;
      end
    end
    if (reset) begin
      _T_3890_54 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_54 <= _T_4788;
      end
    end
    if (reset) begin
      _T_3890_55 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_55 <= _T_4790;
      end
    end
    if (reset) begin
      _T_3890_56 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_56 <= _T_4792;
      end
    end
    if (reset) begin
      _T_3890_57 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_57 <= _T_4794;
      end
    end
    if (reset) begin
      _T_3890_58 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_58 <= _T_4796;
      end
    end
    if (reset) begin
      _T_3890_59 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_59 <= _T_4798;
      end
    end
    if (reset) begin
      _T_3890_60 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_60 <= _T_4800;
      end
    end
    if (reset) begin
      _T_3890_61 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_61 <= _T_4802;
      end
    end
    if (reset) begin
      _T_3890_62 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_62 <= _T_4804;
      end
    end
    if (reset) begin
      _T_3890_63 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_3890_63 <= _T_4806;
      end
    end
    if (reset) begin
      _T_4161_0 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_0 <= _T_4878;
      end
    end
    if (reset) begin
      _T_4161_1 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_1 <= _T_4879;
      end
    end
    if (reset) begin
      _T_4161_2 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_2 <= _T_4880;
      end
    end
    if (reset) begin
      _T_4161_3 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_3 <= _T_4881;
      end
    end
    if (reset) begin
      _T_4161_4 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_4 <= _T_4882;
      end
    end
    if (reset) begin
      _T_4161_5 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_5 <= _T_4883;
      end
    end
    if (reset) begin
      _T_4161_6 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_6 <= _T_4884;
      end
    end
    if (reset) begin
      _T_4161_7 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_7 <= _T_4885;
      end
    end
    if (reset) begin
      _T_4161_8 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_8 <= _T_4886;
      end
    end
    if (reset) begin
      _T_4161_9 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_9 <= _T_4887;
      end
    end
    if (reset) begin
      _T_4161_10 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_10 <= _T_4888;
      end
    end
    if (reset) begin
      _T_4161_11 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_11 <= _T_4889;
      end
    end
    if (reset) begin
      _T_4161_12 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_12 <= _T_4890;
      end
    end
    if (reset) begin
      _T_4161_13 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_13 <= _T_4891;
      end
    end
    if (reset) begin
      _T_4161_14 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_14 <= _T_4892;
      end
    end
    if (reset) begin
      _T_4161_15 <= 1'h0;
    end else begin
      if (_T_4877) begin
        _T_4161_15 <= _T_4893;
      end
    end
    if (reset) begin
      _T_4288_0 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_0 <= _T_4917;
      end
    end
    if (reset) begin
      _T_4288_1 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_1 <= _T_4918;
      end
    end
    if (reset) begin
      _T_4288_2 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_2 <= _T_4919;
      end
    end
    if (reset) begin
      _T_4288_3 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_3 <= _T_4920;
      end
    end
    if (reset) begin
      _T_4288_4 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_4 <= _T_4921;
      end
    end
    if (reset) begin
      _T_4288_5 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_5 <= _T_4922;
      end
    end
    if (reset) begin
      _T_4288_6 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_6 <= _T_4923;
      end
    end
    if (reset) begin
      _T_4288_7 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_7 <= _T_4924;
      end
    end
    if (reset) begin
      _T_4288_8 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_8 <= _T_4925;
      end
    end
    if (reset) begin
      _T_4288_9 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_9 <= _T_4926;
      end
    end
    if (reset) begin
      _T_4288_10 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_10 <= _T_4927;
      end
    end
    if (reset) begin
      _T_4288_11 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_11 <= _T_4928;
      end
    end
    if (reset) begin
      _T_4288_12 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_12 <= _T_4929;
      end
    end
    if (reset) begin
      _T_4288_13 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_13 <= _T_4930;
      end
    end
    if (reset) begin
      _T_4288_14 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_14 <= _T_4931;
      end
    end
    if (reset) begin
      _T_4288_15 <= 1'h0;
    end else begin
      if (_T_4916) begin
        _T_4288_15 <= _T_4932;
      end
    end
    if (_T_4482) begin
      _T_4344_0 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_0;
    end
    if (_T_4484) begin
      _T_4344_1 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_1;
    end
    if (_T_4486) begin
      _T_4344_2 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_2;
    end
    if (_T_4488) begin
      _T_4344_3 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_3;
    end
    if (_T_4490) begin
      _T_4344_4 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_4;
    end
    if (_T_4492) begin
      _T_4344_5 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_5;
    end
    if (_T_4494) begin
      _T_4344_6 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_6;
    end
    if (_T_4496) begin
      _T_4344_7 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_7;
    end
    if (_T_4498) begin
      _T_4344_8 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_8;
    end
    if (_T_4500) begin
      _T_4344_9 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_9;
    end
    if (_T_4502) begin
      _T_4344_10 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_10;
    end
    if (_T_4504) begin
      _T_4344_11 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_11;
    end
    if (_T_4506) begin
      _T_4344_12 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_12;
    end
    if (_T_4508) begin
      _T_4344_13 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_13;
    end
    if (_T_4510) begin
      _T_4344_14 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_14;
    end
    if (_T_4512) begin
      _T_4344_15 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_15;
    end
    if (_T_4514) begin
      _T_4344_16 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_16;
    end
    if (_T_4516) begin
      _T_4344_17 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_17;
    end
    if (_T_4518) begin
      _T_4344_18 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_18;
    end
    if (_T_4520) begin
      _T_4344_19 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_19;
    end
    if (_T_4522) begin
      _T_4344_20 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_20;
    end
    if (_T_4524) begin
      _T_4344_21 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_21;
    end
    if (_T_4526) begin
      _T_4344_22 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_22;
    end
    if (_T_4528) begin
      _T_4344_23 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_23;
    end
    if (_T_4530) begin
      _T_4344_24 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_24;
    end
    if (_T_4532) begin
      _T_4344_25 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_25;
    end
    if (_T_4534) begin
      _T_4344_26 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_26;
    end
    if (_T_4536) begin
      _T_4344_27 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_27;
    end
    if (_T_4538) begin
      _T_4344_28 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_28;
    end
    if (_T_4540) begin
      _T_4344_29 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_29;
    end
    if (_T_4542) begin
      _T_4344_30 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_30;
    end
    if (_T_4544) begin
      _T_4344_31 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_31;
    end
    if (_T_4546) begin
      _T_4344_32 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_32;
    end
    if (_T_4548) begin
      _T_4344_33 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_33;
    end
    if (_T_4550) begin
      _T_4344_34 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_34;
    end
    if (_T_4552) begin
      _T_4344_35 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_35;
    end
    if (_T_4554) begin
      _T_4344_36 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_36;
    end
    if (_T_4556) begin
      _T_4344_37 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_37;
    end
    if (_T_4558) begin
      _T_4344_38 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_38;
    end
    if (_T_4560) begin
      _T_4344_39 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_39;
    end
    if (_T_4562) begin
      _T_4344_40 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_40;
    end
    if (_T_4564) begin
      _T_4344_41 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_41;
    end
    if (_T_4566) begin
      _T_4344_42 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_42;
    end
    if (_T_4568) begin
      _T_4344_43 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_43;
    end
    if (_T_4570) begin
      _T_4344_44 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_44;
    end
    if (_T_4572) begin
      _T_4344_45 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_45;
    end
    if (_T_4574) begin
      _T_4344_46 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_46;
    end
    if (_T_4576) begin
      _T_4344_47 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_47;
    end
    if (_T_4578) begin
      _T_4344_48 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_48;
    end
    if (_T_4580) begin
      _T_4344_49 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_49;
    end
    if (_T_4582) begin
      _T_4344_50 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_50;
    end
    if (_T_4584) begin
      _T_4344_51 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_51;
    end
    if (_T_4586) begin
      _T_4344_52 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_52;
    end
    if (_T_4588) begin
      _T_4344_53 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_53;
    end
    if (_T_4590) begin
      _T_4344_54 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_54;
    end
    if (_T_4592) begin
      _T_4344_55 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_55;
    end
    if (_T_4594) begin
      _T_4344_56 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_56;
    end
    if (_T_4596) begin
      _T_4344_57 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_57;
    end
    if (_T_4598) begin
      _T_4344_58 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_58;
    end
    if (_T_4600) begin
      _T_4344_59 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_59;
    end
    if (_T_4602) begin
      _T_4344_60 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_60;
    end
    if (_T_4604) begin
      _T_4344_61 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_61;
    end
    if (_T_4606) begin
      _T_4344_62 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_62;
    end
    if (_T_4608) begin
      _T_4344_63 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_63;
    end
    if (_T_4680) begin
      _T_4414_0 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_0;
    end
    if (_T_4682) begin
      _T_4414_1 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_1;
    end
    if (_T_4684) begin
      _T_4414_2 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_2;
    end
    if (_T_4686) begin
      _T_4414_3 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_3;
    end
    if (_T_4688) begin
      _T_4414_4 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_4;
    end
    if (_T_4690) begin
      _T_4414_5 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_5;
    end
    if (_T_4692) begin
      _T_4414_6 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_6;
    end
    if (_T_4694) begin
      _T_4414_7 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_7;
    end
    if (_T_4696) begin
      _T_4414_8 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_8;
    end
    if (_T_4698) begin
      _T_4414_9 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_9;
    end
    if (_T_4700) begin
      _T_4414_10 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_10;
    end
    if (_T_4702) begin
      _T_4414_11 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_11;
    end
    if (_T_4704) begin
      _T_4414_12 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_12;
    end
    if (_T_4706) begin
      _T_4414_13 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_13;
    end
    if (_T_4708) begin
      _T_4414_14 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_14;
    end
    if (_T_4710) begin
      _T_4414_15 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_15;
    end
    if (_T_4712) begin
      _T_4414_16 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_16;
    end
    if (_T_4714) begin
      _T_4414_17 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_17;
    end
    if (_T_4716) begin
      _T_4414_18 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_18;
    end
    if (_T_4718) begin
      _T_4414_19 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_19;
    end
    if (_T_4720) begin
      _T_4414_20 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_20;
    end
    if (_T_4722) begin
      _T_4414_21 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_21;
    end
    if (_T_4724) begin
      _T_4414_22 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_22;
    end
    if (_T_4726) begin
      _T_4414_23 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_23;
    end
    if (_T_4728) begin
      _T_4414_24 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_24;
    end
    if (_T_4730) begin
      _T_4414_25 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_25;
    end
    if (_T_4732) begin
      _T_4414_26 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_26;
    end
    if (_T_4734) begin
      _T_4414_27 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_27;
    end
    if (_T_4736) begin
      _T_4414_28 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_28;
    end
    if (_T_4738) begin
      _T_4414_29 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_29;
    end
    if (_T_4740) begin
      _T_4414_30 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_30;
    end
    if (_T_4742) begin
      _T_4414_31 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_31;
    end
    if (_T_4744) begin
      _T_4414_32 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_32;
    end
    if (_T_4746) begin
      _T_4414_33 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_33;
    end
    if (_T_4748) begin
      _T_4414_34 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_34;
    end
    if (_T_4750) begin
      _T_4414_35 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_35;
    end
    if (_T_4752) begin
      _T_4414_36 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_36;
    end
    if (_T_4754) begin
      _T_4414_37 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_37;
    end
    if (_T_4756) begin
      _T_4414_38 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_38;
    end
    if (_T_4758) begin
      _T_4414_39 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_39;
    end
    if (_T_4760) begin
      _T_4414_40 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_40;
    end
    if (_T_4762) begin
      _T_4414_41 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_41;
    end
    if (_T_4764) begin
      _T_4414_42 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_42;
    end
    if (_T_4766) begin
      _T_4414_43 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_43;
    end
    if (_T_4768) begin
      _T_4414_44 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_44;
    end
    if (_T_4770) begin
      _T_4414_45 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_45;
    end
    if (_T_4772) begin
      _T_4414_46 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_46;
    end
    if (_T_4774) begin
      _T_4414_47 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_47;
    end
    if (_T_4776) begin
      _T_4414_48 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_48;
    end
    if (_T_4778) begin
      _T_4414_49 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_49;
    end
    if (_T_4780) begin
      _T_4414_50 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_50;
    end
    if (_T_4782) begin
      _T_4414_51 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_51;
    end
    if (_T_4784) begin
      _T_4414_52 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_52;
    end
    if (_T_4786) begin
      _T_4414_53 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_53;
    end
    if (_T_4788) begin
      _T_4414_54 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_54;
    end
    if (_T_4790) begin
      _T_4414_55 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_55;
    end
    if (_T_4792) begin
      _T_4414_56 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_56;
    end
    if (_T_4794) begin
      _T_4414_57 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_57;
    end
    if (_T_4796) begin
      _T_4414_58 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_58;
    end
    if (_T_4798) begin
      _T_4414_59 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_59;
    end
    if (_T_4800) begin
      _T_4414_60 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_60;
    end
    if (_T_4802) begin
      _T_4414_61 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_61;
    end
    if (_T_4804) begin
      _T_4414_62 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_62;
    end
    if (_T_4806) begin
      _T_4414_63 <= NV_NVDLA_CSC_WL_dec_io_output_bits_data_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_798 <= 15'h0;
    end else begin
      if (_T_847) begin
        if (io_sc2cdma_wt_pending_req) begin
          _T_798 <= 15'h0;
        end else begin
          if (!(_T_810)) begin
            if (_T_808) begin
              _T_798 <= _T_805;
            end else begin
              _T_798 <= _T_800;
            end
          end
        end
      end
    end
  end
endmodule
