module NV_NVDLA_CDMA_single_reg( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_reg_rd_data, // @[:@6.4]
  input  [11:0] io_reg_offset, // @[:@6.4]
  input  [31:0] io_reg_wr_data, // @[:@6.4]
  input         io_reg_wr_en, // @[:@6.4]
  output        io_producer, // @[:@6.4]
  output [3:0]  io_arb_wmb, // @[:@6.4]
  input         io_flush_done, // @[:@6.4]
  input         io_consumer, // @[:@6.4]
  input  [1:0]  io_status_0, // @[:@6.4]
  input  [1:0]  io_status_1 // @[:@6.4]
);
  wire [31:0] _GEN_3; // @[NV_NVDLA_CDMA_single_reg.scala 48:54:@8.4]
  wire  _T_30; // @[NV_NVDLA_CDMA_single_reg.scala 48:54:@8.4]
  wire  nvdla_cdma_s_arbiter_0_wren; // @[NV_NVDLA_CDMA_single_reg.scala 48:76:@9.4]
  wire  _T_34; // @[NV_NVDLA_CDMA_single_reg.scala 50:54:@12.4]
  wire  nvdla_cdma_s_pointer_0_wren; // @[NV_NVDLA_CDMA_single_reg.scala 50:76:@13.4]
  wire [31:0] _T_43; // @[Cat.scala 30:58:@18.4]
  wire [31:0] _T_46; // @[Cat.scala 30:58:@19.4]
  wire [31:0] _T_52; // @[Cat.scala 30:58:@22.4]
  wire [31:0] _T_58; // @[Cat.scala 30:58:@25.4]
  wire  _T_59; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_60; // @[Mux.scala 46:16:@27.4]
  wire  _T_61; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_62; // @[Mux.scala 46:16:@29.4]
  wire  _T_63; // @[Mux.scala 46:19:@30.4]
  wire [31:0] _T_64; // @[Mux.scala 46:16:@31.4]
  wire  _T_65; // @[Mux.scala 46:19:@32.4]
  wire [3:0] _T_71; // @[NV_NVDLA_CDMA_single_reg.scala 68:43:@41.4]
  reg [3:0] _T_74; // @[Reg.scala 19:20:@42.4]
  reg [31:0] _RAND_0;
  wire [3:0] _GEN_1; // @[Reg.scala 20:19:@43.4]
  wire  _T_75; // @[NV_NVDLA_CDMA_single_reg.scala 69:44:@47.4]
  reg  _T_78; // @[Reg.scala 19:20:@48.4]
  reg [31:0] _RAND_1;
  wire  _GEN_2; // @[Reg.scala 20:19:@49.4]
  assign _GEN_3 = {{20'd0}, io_reg_offset}; // @[NV_NVDLA_CDMA_single_reg.scala 48:54:@8.4]
  assign _T_30 = _GEN_3 == 32'h8; // @[NV_NVDLA_CDMA_single_reg.scala 48:54:@8.4]
  assign nvdla_cdma_s_arbiter_0_wren = _T_30 & io_reg_wr_en; // @[NV_NVDLA_CDMA_single_reg.scala 48:76:@9.4]
  assign _T_34 = _GEN_3 == 32'h4; // @[NV_NVDLA_CDMA_single_reg.scala 50:54:@12.4]
  assign nvdla_cdma_s_pointer_0_wren = _T_34 & io_reg_wr_en; // @[NV_NVDLA_CDMA_single_reg.scala 50:76:@13.4]
  assign _T_43 = {12'h0,io_arb_wmb,15'h0,io_producer}; // @[Cat.scala 30:58:@18.4]
  assign _T_46 = {31'h0,io_flush_done}; // @[Cat.scala 30:58:@19.4]
  assign _T_52 = {15'h0,io_consumer,15'h0,io_producer}; // @[Cat.scala 30:58:@22.4]
  assign _T_58 = {14'h0,io_status_1,14'h0,io_status_0}; // @[Cat.scala 30:58:@25.4]
  assign _T_59 = 32'h0 == _GEN_3; // @[Mux.scala 46:19:@26.4]
  assign _T_60 = _T_59 ? _T_58 : 32'h0; // @[Mux.scala 46:16:@27.4]
  assign _T_61 = 32'h4 == _GEN_3; // @[Mux.scala 46:19:@28.4]
  assign _T_62 = _T_61 ? _T_52 : _T_60; // @[Mux.scala 46:16:@29.4]
  assign _T_63 = 32'hc == _GEN_3; // @[Mux.scala 46:19:@30.4]
  assign _T_64 = _T_63 ? _T_46 : _T_62; // @[Mux.scala 46:16:@31.4]
  assign _T_65 = 32'h8 == _GEN_3; // @[Mux.scala 46:19:@32.4]
  assign _T_71 = io_reg_wr_data[19:16]; // @[NV_NVDLA_CDMA_single_reg.scala 68:43:@41.4]
  assign _GEN_1 = nvdla_cdma_s_arbiter_0_wren ? _T_71 : _T_74; // @[Reg.scala 20:19:@43.4]
  assign _T_75 = io_reg_wr_data[0]; // @[NV_NVDLA_CDMA_single_reg.scala 69:44:@47.4]
  assign _GEN_2 = nvdla_cdma_s_pointer_0_wren ? _T_75 : _T_78; // @[Reg.scala 20:19:@49.4]
  assign io_reg_rd_data = _T_65 ? _T_43 : _T_64; // @[NV_NVDLA_CDMA_single_reg.scala 54:20:@34.4]
  assign io_producer = _T_78; // @[NV_NVDLA_CDMA_single_reg.scala 69:17:@52.4]
  assign io_arb_wmb = _T_74; // @[NV_NVDLA_CDMA_single_reg.scala 68:16:@46.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_74 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_78 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_74 <= 4'h3;
    end else begin
      if (nvdla_cdma_s_arbiter_0_wren) begin
        _T_74 <= _T_71;
      end
    end
    if (reset) begin
      _T_78 <= 1'h0;
    end else begin
      if (nvdla_cdma_s_pointer_0_wren) begin
        _T_78 <= _T_75;
      end
    end
  end
endmodule
module NV_NVDLA_CDMA_dual_reg( // @[:@54.2]
  input         reset, // @[:@56.4]
  input         io_nvdla_core_clk, // @[:@57.4]
  output [31:0] io_reg_rd_data, // @[:@57.4]
  input  [11:0] io_reg_offset, // @[:@57.4]
  input  [31:0] io_reg_wr_data, // @[:@57.4]
  input         io_reg_wr_en, // @[:@57.4]
  output [4:0]  io_field_data_bank, // @[:@57.4]
  output [4:0]  io_field_weight_bank, // @[:@57.4]
  output [4:0]  io_field_batches, // @[:@57.4]
  output [31:0] io_field_batch_stride, // @[:@57.4]
  output [2:0]  io_field_conv_x_stride, // @[:@57.4]
  output [2:0]  io_field_conv_y_stride, // @[:@57.4]
  output        io_field_cvt_en, // @[:@57.4]
  output [5:0]  io_field_cvt_truncate, // @[:@57.4]
  output [15:0] io_field_cvt_offset, // @[:@57.4]
  output [15:0] io_field_cvt_scale, // @[:@57.4]
  output [31:0] io_field_cya, // @[:@57.4]
  output [31:0] io_field_datain_addr_high_0, // @[:@57.4]
  output [31:0] io_field_datain_addr_high_1, // @[:@57.4]
  output [31:0] io_field_datain_addr_low_0, // @[:@57.4]
  output [31:0] io_field_datain_addr_low_1, // @[:@57.4]
  output        io_field_line_packed, // @[:@57.4]
  output        io_field_surf_packed, // @[:@57.4]
  output        io_field_datain_ram_type, // @[:@57.4]
  output        io_field_datain_format, // @[:@57.4]
  output [5:0]  io_field_pixel_format, // @[:@57.4]
  output        io_field_pixel_mapping, // @[:@57.4]
  output        io_field_pixel_sign_override, // @[:@57.4]
  output [12:0] io_field_datain_height, // @[:@57.4]
  output [12:0] io_field_datain_width, // @[:@57.4]
  output [12:0] io_field_datain_channel, // @[:@57.4]
  output [12:0] io_field_datain_height_ext, // @[:@57.4]
  output [12:0] io_field_datain_width_ext, // @[:@57.4]
  output [13:0] io_field_entries, // @[:@57.4]
  output [11:0] io_field_grains, // @[:@57.4]
  output [31:0] io_field_line_stride, // @[:@57.4]
  output [31:0] io_field_uv_line_stride, // @[:@57.4]
  output        io_field_mean_format, // @[:@57.4]
  output [15:0] io_field_mean_gu, // @[:@57.4]
  output [15:0] io_field_mean_ry, // @[:@57.4]
  output [15:0] io_field_mean_ax, // @[:@57.4]
  output [15:0] io_field_mean_bv, // @[:@57.4]
  output        io_field_conv_mode, // @[:@57.4]
  output        io_field_data_reuse, // @[:@57.4]
  output [1:0]  io_field_in_precision, // @[:@57.4]
  output [1:0]  io_field_proc_precision, // @[:@57.4]
  output        io_field_skip_data_rls, // @[:@57.4]
  output        io_field_skip_weight_rls, // @[:@57.4]
  output        io_field_weight_reuse, // @[:@57.4]
  output        io_field_nan_to_zero, // @[:@57.4]
  output        io_field_dma_en, // @[:@57.4]
  output [4:0]  io_field_pixel_x_offset, // @[:@57.4]
  output [2:0]  io_field_pixel_y_offset, // @[:@57.4]
  output [9:0]  io_field_rsv_per_line, // @[:@57.4]
  output [9:0]  io_field_rsv_per_uv_line, // @[:@57.4]
  output [2:0]  io_field_rsv_height, // @[:@57.4]
  output [4:0]  io_field_rsv_y_index, // @[:@57.4]
  output [31:0] io_field_surf_stride, // @[:@57.4]
  output [31:0] io_field_weight_addr_high, // @[:@57.4]
  output [31:0] io_field_weight_addr_low, // @[:@57.4]
  output [31:0] io_field_weight_bytes, // @[:@57.4]
  output        io_field_weight_format, // @[:@57.4]
  output        io_field_weight_ram_type, // @[:@57.4]
  output [17:0] io_field_byte_per_kernel, // @[:@57.4]
  output [12:0] io_field_weight_kernel, // @[:@57.4]
  output [31:0] io_field_wgs_addr_high, // @[:@57.4]
  output [31:0] io_field_wgs_addr_low, // @[:@57.4]
  output [31:0] io_field_wmb_addr_high, // @[:@57.4]
  output [31:0] io_field_wmb_addr_low, // @[:@57.4]
  output [27:0] io_field_wmb_bytes, // @[:@57.4]
  output [5:0]  io_field_pad_bottom, // @[:@57.4]
  output [4:0]  io_field_pad_left, // @[:@57.4]
  output [5:0]  io_field_pad_right, // @[:@57.4]
  output [4:0]  io_field_pad_top, // @[:@57.4]
  output [15:0] io_field_pad_value, // @[:@57.4]
  output        io_op_en_trigger, // @[:@57.4]
  input  [31:0] io_inf_data_num, // @[:@57.4]
  input  [31:0] io_inf_weight_num, // @[:@57.4]
  input  [31:0] io_nan_data_num, // @[:@57.4]
  input  [31:0] io_nan_weight_num, // @[:@57.4]
  input         io_op_en, // @[:@57.4]
  input  [31:0] io_dat_rd_latency, // @[:@57.4]
  input  [31:0] io_dat_rd_stall, // @[:@57.4]
  input  [31:0] io_wt_rd_latency, // @[:@57.4]
  input  [31:0] io_wt_rd_stall // @[:@57.4]
);
  wire [31:0] _GEN_69; // @[NV_NVDLA_CDMA_dual_reg.scala 54:51:@59.4]
  wire  _T_174; // @[NV_NVDLA_CDMA_dual_reg.scala 54:51:@59.4]
  wire  _T_175; // @[NV_NVDLA_CDMA_dual_reg.scala 54:75:@60.4]
  wire  _T_177; // @[NV_NVDLA_CDMA_dual_reg.scala 55:59:@61.4]
  wire  _T_178; // @[NV_NVDLA_CDMA_dual_reg.scala 55:83:@62.4]
  wire  _T_180; // @[NV_NVDLA_CDMA_dual_reg.scala 56:59:@63.4]
  wire  _T_181; // @[NV_NVDLA_CDMA_dual_reg.scala 56:83:@64.4]
  wire  _T_183; // @[NV_NVDLA_CDMA_dual_reg.scala 57:58:@65.4]
  wire  _T_184; // @[NV_NVDLA_CDMA_dual_reg.scala 57:82:@66.4]
  wire  _T_186; // @[NV_NVDLA_CDMA_dual_reg.scala 58:54:@67.4]
  wire  _T_187; // @[NV_NVDLA_CDMA_dual_reg.scala 58:78:@68.4]
  wire  _T_189; // @[NV_NVDLA_CDMA_dual_reg.scala 59:57:@69.4]
  wire  _T_190; // @[NV_NVDLA_CDMA_dual_reg.scala 59:81:@70.4]
  wire  _T_192; // @[NV_NVDLA_CDMA_dual_reg.scala 60:56:@71.4]
  wire  _T_193; // @[NV_NVDLA_CDMA_dual_reg.scala 60:80:@72.4]
  wire  _T_195; // @[NV_NVDLA_CDMA_dual_reg.scala 61:50:@73.4]
  wire  _T_196; // @[NV_NVDLA_CDMA_dual_reg.scala 61:74:@74.4]
  wire  _T_198; // @[NV_NVDLA_CDMA_dual_reg.scala 62:63:@75.4]
  wire  _T_199; // @[NV_NVDLA_CDMA_dual_reg.scala 62:87:@76.4]
  wire  _T_201; // @[NV_NVDLA_CDMA_dual_reg.scala 63:63:@77.4]
  wire  _T_202; // @[NV_NVDLA_CDMA_dual_reg.scala 63:87:@78.4]
  wire  _T_204; // @[NV_NVDLA_CDMA_dual_reg.scala 64:62:@79.4]
  wire  _T_205; // @[NV_NVDLA_CDMA_dual_reg.scala 64:86:@80.4]
  wire  _T_207; // @[NV_NVDLA_CDMA_dual_reg.scala 65:62:@81.4]
  wire  _T_208; // @[NV_NVDLA_CDMA_dual_reg.scala 65:86:@82.4]
  wire  _T_210; // @[NV_NVDLA_CDMA_dual_reg.scala 66:55:@83.4]
  wire  _T_211; // @[NV_NVDLA_CDMA_dual_reg.scala 66:79:@84.4]
  wire  _T_213; // @[NV_NVDLA_CDMA_dual_reg.scala 67:60:@85.4]
  wire  _T_214; // @[NV_NVDLA_CDMA_dual_reg.scala 67:84:@86.4]
  wire  _T_216; // @[NV_NVDLA_CDMA_dual_reg.scala 68:60:@87.4]
  wire  _T_217; // @[NV_NVDLA_CDMA_dual_reg.scala 68:84:@88.4]
  wire  _T_219; // @[NV_NVDLA_CDMA_dual_reg.scala 69:60:@89.4]
  wire  _T_220; // @[NV_NVDLA_CDMA_dual_reg.scala 69:84:@90.4]
  wire  _T_222; // @[NV_NVDLA_CDMA_dual_reg.scala 70:60:@91.4]
  wire  _T_223; // @[NV_NVDLA_CDMA_dual_reg.scala 70:84:@92.4]
  wire  _T_225; // @[NV_NVDLA_CDMA_dual_reg.scala 71:64:@93.4]
  wire  _T_226; // @[NV_NVDLA_CDMA_dual_reg.scala 71:88:@94.4]
  wire  _T_228; // @[NV_NVDLA_CDMA_dual_reg.scala 72:62:@95.4]
  wire  _T_229; // @[NV_NVDLA_CDMA_dual_reg.scala 72:86:@96.4]
  wire  _T_231; // @[NV_NVDLA_CDMA_dual_reg.scala 73:58:@97.4]
  wire  _T_232; // @[NV_NVDLA_CDMA_dual_reg.scala 73:82:@98.4]
  wire  _T_240; // @[NV_NVDLA_CDMA_dual_reg.scala 76:58:@103.4]
  wire  _T_241; // @[NV_NVDLA_CDMA_dual_reg.scala 76:82:@104.4]
  wire  _T_243; // @[NV_NVDLA_CDMA_dual_reg.scala 77:61:@105.4]
  wire  _T_244; // @[NV_NVDLA_CDMA_dual_reg.scala 77:85:@106.4]
  wire  _T_246; // @[NV_NVDLA_CDMA_dual_reg.scala 78:58:@107.4]
  wire  _T_247; // @[NV_NVDLA_CDMA_dual_reg.scala 78:82:@108.4]
  wire  _T_249; // @[NV_NVDLA_CDMA_dual_reg.scala 79:60:@109.4]
  wire  _T_250; // @[NV_NVDLA_CDMA_dual_reg.scala 79:84:@110.4]
  wire  _T_252; // @[NV_NVDLA_CDMA_dual_reg.scala 80:60:@111.4]
  wire  _T_253; // @[NV_NVDLA_CDMA_dual_reg.scala 80:84:@112.4]
  wire  _T_255; // @[NV_NVDLA_CDMA_dual_reg.scala 81:55:@113.4]
  wire  _T_256; // @[NV_NVDLA_CDMA_dual_reg.scala 81:79:@114.4]
  wire  _T_258; // @[NV_NVDLA_CDMA_dual_reg.scala 82:64:@115.4]
  wire  _T_259; // @[NV_NVDLA_CDMA_dual_reg.scala 82:88:@116.4]
  wire  _T_267; // @[NV_NVDLA_CDMA_dual_reg.scala 85:56:@121.4]
  wire  _T_276; // @[NV_NVDLA_CDMA_dual_reg.scala 88:58:@127.4]
  wire  _T_277; // @[NV_NVDLA_CDMA_dual_reg.scala 88:82:@128.4]
  wire  _T_285; // @[NV_NVDLA_CDMA_dual_reg.scala 91:59:@133.4]
  wire  _T_286; // @[NV_NVDLA_CDMA_dual_reg.scala 91:83:@134.4]
  wire  _T_288; // @[NV_NVDLA_CDMA_dual_reg.scala 92:61:@135.4]
  wire  _T_289; // @[NV_NVDLA_CDMA_dual_reg.scala 92:85:@136.4]
  wire  _T_291; // @[NV_NVDLA_CDMA_dual_reg.scala 93:61:@137.4]
  wire  _T_292; // @[NV_NVDLA_CDMA_dual_reg.scala 93:85:@138.4]
  wire  _T_294; // @[NV_NVDLA_CDMA_dual_reg.scala 94:58:@139.4]
  wire  _T_295; // @[NV_NVDLA_CDMA_dual_reg.scala 94:82:@140.4]
  wire  _T_297; // @[NV_NVDLA_CDMA_dual_reg.scala 95:63:@141.4]
  wire  _T_298; // @[NV_NVDLA_CDMA_dual_reg.scala 95:87:@142.4]
  wire  _T_300; // @[NV_NVDLA_CDMA_dual_reg.scala 96:62:@143.4]
  wire  _T_301; // @[NV_NVDLA_CDMA_dual_reg.scala 96:86:@144.4]
  wire  _T_303; // @[NV_NVDLA_CDMA_dual_reg.scala 97:59:@145.4]
  wire  _T_304; // @[NV_NVDLA_CDMA_dual_reg.scala 97:83:@146.4]
  wire  _T_306; // @[NV_NVDLA_CDMA_dual_reg.scala 98:60:@147.4]
  wire  _T_307; // @[NV_NVDLA_CDMA_dual_reg.scala 98:84:@148.4]
  wire  _T_309; // @[NV_NVDLA_CDMA_dual_reg.scala 99:62:@149.4]
  wire  _T_310; // @[NV_NVDLA_CDMA_dual_reg.scala 99:86:@150.4]
  wire  _T_312; // @[NV_NVDLA_CDMA_dual_reg.scala 100:60:@151.4]
  wire  _T_313; // @[NV_NVDLA_CDMA_dual_reg.scala 100:84:@152.4]
  wire  _T_315; // @[NV_NVDLA_CDMA_dual_reg.scala 101:60:@153.4]
  wire  _T_316; // @[NV_NVDLA_CDMA_dual_reg.scala 101:84:@154.4]
  wire  _T_318; // @[NV_NVDLA_CDMA_dual_reg.scala 102:60:@155.4]
  wire  _T_319; // @[NV_NVDLA_CDMA_dual_reg.scala 102:84:@156.4]
  wire  _T_321; // @[NV_NVDLA_CDMA_dual_reg.scala 103:59:@157.4]
  wire  _T_322; // @[NV_NVDLA_CDMA_dual_reg.scala 103:83:@158.4]
  wire  _T_324; // @[NV_NVDLA_CDMA_dual_reg.scala 104:60:@159.4]
  wire  _T_325; // @[NV_NVDLA_CDMA_dual_reg.scala 104:84:@160.4]
  wire  _T_327; // @[NV_NVDLA_CDMA_dual_reg.scala 105:59:@161.4]
  wire  _T_328; // @[NV_NVDLA_CDMA_dual_reg.scala 105:83:@162.4]
  wire  _T_330; // @[NV_NVDLA_CDMA_dual_reg.scala 106:56:@163.4]
  wire  _T_331; // @[NV_NVDLA_CDMA_dual_reg.scala 106:80:@164.4]
  wire  _T_333; // @[NV_NVDLA_CDMA_dual_reg.scala 107:59:@165.4]
  wire  _T_334; // @[NV_NVDLA_CDMA_dual_reg.scala 107:83:@166.4]
  wire  _T_336; // @[NV_NVDLA_CDMA_dual_reg.scala 108:65:@167.4]
  wire  _T_337; // @[NV_NVDLA_CDMA_dual_reg.scala 108:89:@168.4]
  wire [31:0] _T_344; // @[Cat.scala 30:58:@172.4]
  wire [31:0] _T_347; // @[Cat.scala 30:58:@173.4]
  wire [31:0] _T_354; // @[Cat.scala 30:58:@176.4]
  wire [31:0] _T_360; // @[Cat.scala 30:58:@179.4]
  wire [31:0] _T_363; // @[Cat.scala 30:58:@180.4]
  wire [31:0] _T_366; // @[Cat.scala 30:58:@181.4]
  wire [31:0] _T_377; // @[Cat.scala 30:58:@184.4]
  wire [31:0] _T_380; // @[Cat.scala 30:58:@185.4]
  wire [31:0] _T_392; // @[Cat.scala 30:58:@192.4]
  wire [31:0] _T_398; // @[Cat.scala 30:58:@195.4]
  wire [31:0] _T_401; // @[Cat.scala 30:58:@196.4]
  wire [31:0] _T_407; // @[Cat.scala 30:58:@199.4]
  wire [31:0] _T_410; // @[Cat.scala 30:58:@200.4]
  wire [31:0] _T_413; // @[Cat.scala 30:58:@201.4]
  wire [31:0] _T_420; // @[Cat.scala 30:58:@202.4]
  wire [31:0] _T_422; // @[Cat.scala 30:58:@203.4]
  wire [31:0] _T_424; // @[Cat.scala 30:58:@204.4]
  wire [16:0] _T_438; // @[Cat.scala 30:58:@210.4]
  wire [31:0] _T_445; // @[Cat.scala 30:58:@217.4]
  wire [31:0] _T_448; // @[Cat.scala 30:58:@218.4]
  wire [31:0] _T_453; // @[Cat.scala 30:58:@219.4]
  wire [31:0] _T_458; // @[Cat.scala 30:58:@220.4]
  wire [31:0] _T_466; // @[Cat.scala 30:58:@223.4]
  wire [31:0] _T_472; // @[Cat.scala 30:58:@226.4]
  wire [31:0] _T_478; // @[Cat.scala 30:58:@229.4]
  wire [31:0] _T_485; // @[Cat.scala 30:58:@230.4]
  wire [31:0] _T_488; // @[Cat.scala 30:58:@231.4]
  wire [31:0] _T_491; // @[Cat.scala 30:58:@232.4]
  wire [31:0] _T_494; // @[Cat.scala 30:58:@233.4]
  wire [31:0] _T_501; // @[Cat.scala 30:58:@234.4]
  wire [31:0] _T_513; // @[Cat.scala 30:58:@241.4]
  wire [31:0] _T_516; // @[Cat.scala 30:58:@242.4]
  wire  _T_517; // @[Mux.scala 46:19:@243.4]
  wire [31:0] _T_518; // @[Mux.scala 46:16:@244.4]
  wire  _T_519; // @[Mux.scala 46:19:@245.4]
  wire [31:0] _T_520; // @[Mux.scala 46:16:@246.4]
  wire  _T_521; // @[Mux.scala 46:19:@247.4]
  wire [31:0] _T_522; // @[Mux.scala 46:16:@248.4]
  wire  _T_523; // @[Mux.scala 46:19:@249.4]
  wire [31:0] _T_524; // @[Mux.scala 46:16:@250.4]
  wire  _T_525; // @[Mux.scala 46:19:@251.4]
  wire [31:0] _T_526; // @[Mux.scala 46:16:@252.4]
  wire  _T_527; // @[Mux.scala 46:19:@253.4]
  wire [31:0] _T_528; // @[Mux.scala 46:16:@254.4]
  wire  _T_529; // @[Mux.scala 46:19:@255.4]
  wire [31:0] _T_530; // @[Mux.scala 46:16:@256.4]
  wire  _T_531; // @[Mux.scala 46:19:@257.4]
  wire [31:0] _T_532; // @[Mux.scala 46:16:@258.4]
  wire  _T_533; // @[Mux.scala 46:19:@259.4]
  wire [31:0] _T_534; // @[Mux.scala 46:16:@260.4]
  wire  _T_535; // @[Mux.scala 46:19:@261.4]
  wire [31:0] _T_536; // @[Mux.scala 46:16:@262.4]
  wire  _T_537; // @[Mux.scala 46:19:@263.4]
  wire [31:0] _T_538; // @[Mux.scala 46:16:@264.4]
  wire  _T_539; // @[Mux.scala 46:19:@265.4]
  wire [31:0] _T_540; // @[Mux.scala 46:16:@266.4]
  wire  _T_541; // @[Mux.scala 46:19:@267.4]
  wire [31:0] _T_542; // @[Mux.scala 46:16:@268.4]
  wire  _T_543; // @[Mux.scala 46:19:@269.4]
  wire [31:0] _T_544; // @[Mux.scala 46:16:@270.4]
  wire  _T_545; // @[Mux.scala 46:19:@271.4]
  wire [31:0] _T_546; // @[Mux.scala 46:16:@272.4]
  wire  _T_547; // @[Mux.scala 46:19:@273.4]
  wire [31:0] _T_548; // @[Mux.scala 46:16:@274.4]
  wire  _T_549; // @[Mux.scala 46:19:@275.4]
  wire [31:0] _T_550; // @[Mux.scala 46:16:@276.4]
  wire  _T_551; // @[Mux.scala 46:19:@277.4]
  wire [31:0] _T_552; // @[Mux.scala 46:16:@278.4]
  wire  _T_553; // @[Mux.scala 46:19:@279.4]
  wire [31:0] _T_554; // @[Mux.scala 46:16:@280.4]
  wire  _T_555; // @[Mux.scala 46:19:@281.4]
  wire [31:0] _T_556; // @[Mux.scala 46:16:@282.4]
  wire  _T_557; // @[Mux.scala 46:19:@283.4]
  wire [31:0] _T_558; // @[Mux.scala 46:16:@284.4]
  wire  _T_559; // @[Mux.scala 46:19:@285.4]
  wire [31:0] _T_560; // @[Mux.scala 46:16:@286.4]
  wire  _T_561; // @[Mux.scala 46:19:@287.4]
  wire [31:0] _T_562; // @[Mux.scala 46:16:@288.4]
  wire  _T_563; // @[Mux.scala 46:19:@289.4]
  wire [31:0] _T_564; // @[Mux.scala 46:16:@290.4]
  wire  _T_565; // @[Mux.scala 46:19:@291.4]
  wire [31:0] _T_566; // @[Mux.scala 46:16:@292.4]
  wire  _T_567; // @[Mux.scala 46:19:@293.4]
  wire [31:0] _T_568; // @[Mux.scala 46:16:@294.4]
  wire  _T_569; // @[Mux.scala 46:19:@295.4]
  wire [31:0] _T_570; // @[Mux.scala 46:16:@296.4]
  wire  _T_571; // @[Mux.scala 46:19:@297.4]
  wire [31:0] _T_572; // @[Mux.scala 46:16:@298.4]
  wire  _T_573; // @[Mux.scala 46:19:@299.4]
  wire [31:0] _T_574; // @[Mux.scala 46:16:@300.4]
  wire  _T_575; // @[Mux.scala 46:19:@301.4]
  wire [31:0] _T_576; // @[Mux.scala 46:16:@302.4]
  wire  _T_577; // @[Mux.scala 46:19:@303.4]
  wire [31:0] _T_578; // @[Mux.scala 46:16:@304.4]
  wire  _T_579; // @[Mux.scala 46:19:@305.4]
  wire [31:0] _T_580; // @[Mux.scala 46:16:@306.4]
  wire  _T_581; // @[Mux.scala 46:19:@307.4]
  wire [31:0] _T_582; // @[Mux.scala 46:16:@308.4]
  wire  _T_583; // @[Mux.scala 46:19:@309.4]
  wire [31:0] _T_584; // @[Mux.scala 46:16:@310.4]
  wire  _T_585; // @[Mux.scala 46:19:@311.4]
  wire [31:0] _T_586; // @[Mux.scala 46:16:@312.4]
  wire  _T_587; // @[Mux.scala 46:19:@313.4]
  wire [31:0] _T_588; // @[Mux.scala 46:16:@314.4]
  wire  _T_589; // @[Mux.scala 46:19:@315.4]
  wire [31:0] _T_590; // @[Mux.scala 46:16:@316.4]
  wire  _T_591; // @[Mux.scala 46:19:@317.4]
  wire [31:0] _T_592; // @[Mux.scala 46:16:@318.4]
  wire  _T_593; // @[Mux.scala 46:19:@319.4]
  wire [31:0] _T_594; // @[Mux.scala 46:16:@320.4]
  wire  _T_595; // @[Mux.scala 46:19:@321.4]
  wire [31:0] _T_596; // @[Mux.scala 46:16:@322.4]
  wire  _T_597; // @[Mux.scala 46:19:@323.4]
  wire [31:0] _T_598; // @[Mux.scala 46:16:@324.4]
  wire  _T_599; // @[Mux.scala 46:19:@325.4]
  wire [31:0] _T_600; // @[Mux.scala 46:16:@326.4]
  wire  _T_601; // @[Mux.scala 46:19:@327.4]
  wire [31:0] _T_602; // @[Mux.scala 46:16:@328.4]
  wire  _T_603; // @[Mux.scala 46:19:@329.4]
  wire [31:0] _T_604; // @[Mux.scala 46:16:@330.4]
  wire  _T_605; // @[Mux.scala 46:19:@331.4]
  wire [31:0] _T_606; // @[Mux.scala 46:16:@332.4]
  wire  _T_607; // @[Mux.scala 46:19:@333.4]
  wire [31:0] _T_608; // @[Mux.scala 46:16:@334.4]
  wire  _T_609; // @[Mux.scala 46:19:@335.4]
  wire [31:0] _T_610; // @[Mux.scala 46:16:@336.4]
  wire  _T_611; // @[Mux.scala 46:19:@337.4]
  wire [31:0] _T_612; // @[Mux.scala 46:16:@338.4]
  wire  _T_613; // @[Mux.scala 46:19:@339.4]
  wire [31:0] _T_614; // @[Mux.scala 46:16:@340.4]
  wire  _T_615; // @[Mux.scala 46:19:@341.4]
  wire [31:0] _T_616; // @[Mux.scala 46:16:@342.4]
  wire  _T_617; // @[Mux.scala 46:19:@343.4]
  wire [31:0] _T_618; // @[Mux.scala 46:16:@344.4]
  wire  _T_619; // @[Mux.scala 46:19:@345.4]
  wire [31:0] _T_620; // @[Mux.scala 46:16:@346.4]
  wire  _T_621; // @[Mux.scala 46:19:@347.4]
  wire [31:0] _T_622; // @[Mux.scala 46:16:@348.4]
  wire  _T_623; // @[Mux.scala 46:19:@349.4]
  wire [31:0] _T_624; // @[Mux.scala 46:16:@350.4]
  wire  _T_625; // @[Mux.scala 46:19:@351.4]
  wire [4:0] _T_627; // @[NV_NVDLA_CDMA_dual_reg.scala 232:51:@354.4]
  reg [4:0] _T_630; // @[Reg.scala 19:20:@355.4]
  reg [31:0] _RAND_0;
  wire [4:0] _GEN_0; // @[Reg.scala 20:19:@356.4]
  wire [4:0] _T_631; // @[NV_NVDLA_CDMA_dual_reg.scala 234:53:@360.4]
  reg [4:0] _T_634; // @[Reg.scala 19:20:@361.4]
  reg [31:0] _RAND_1;
  wire [4:0] _GEN_1; // @[Reg.scala 20:19:@362.4]
  reg [4:0] _T_638; // @[Reg.scala 19:20:@367.4]
  reg [31:0] _RAND_2;
  wire [4:0] _GEN_2; // @[Reg.scala 20:19:@368.4]
  reg [31:0] _T_642; // @[Reg.scala 19:20:@373.4]
  reg [31:0] _RAND_3;
  wire [31:0] _GEN_3; // @[Reg.scala 20:19:@374.4]
  wire [2:0] _T_643; // @[NV_NVDLA_CDMA_dual_reg.scala 240:55:@378.4]
  reg [2:0] _T_646; // @[Reg.scala 19:20:@379.4]
  reg [31:0] _RAND_4;
  wire [2:0] _GEN_4; // @[Reg.scala 20:19:@380.4]
  wire [2:0] _T_647; // @[NV_NVDLA_CDMA_dual_reg.scala 242:55:@384.4]
  reg [2:0] _T_650; // @[Reg.scala 19:20:@385.4]
  reg [31:0] _RAND_5;
  wire [2:0] _GEN_5; // @[Reg.scala 20:19:@386.4]
  wire  _T_651; // @[NV_NVDLA_CDMA_dual_reg.scala 244:48:@390.4]
  reg  _T_654; // @[Reg.scala 19:20:@391.4]
  reg [31:0] _RAND_6;
  wire  _GEN_6; // @[Reg.scala 20:19:@392.4]
  wire [5:0] _T_655; // @[NV_NVDLA_CDMA_dual_reg.scala 246:54:@396.4]
  reg [5:0] _T_658; // @[Reg.scala 19:20:@397.4]
  reg [31:0] _RAND_7;
  wire [5:0] _GEN_7; // @[Reg.scala 20:19:@398.4]
  wire [15:0] _T_659; // @[NV_NVDLA_CDMA_dual_reg.scala 248:52:@402.4]
  reg [15:0] _T_662; // @[Reg.scala 19:20:@403.4]
  reg [31:0] _RAND_8;
  wire [15:0] _GEN_8; // @[Reg.scala 20:19:@404.4]
  reg [15:0] _T_666; // @[Reg.scala 19:20:@409.4]
  reg [31:0] _RAND_9;
  wire [15:0] _GEN_9; // @[Reg.scala 20:19:@410.4]
  reg [31:0] _T_670; // @[Reg.scala 19:20:@415.4]
  reg [31:0] _RAND_10;
  wire [31:0] _GEN_10; // @[Reg.scala 20:19:@416.4]
  reg [31:0] _T_674; // @[Reg.scala 19:20:@421.4]
  reg [31:0] _RAND_11;
  wire [31:0] _GEN_11; // @[Reg.scala 20:19:@422.4]
  reg [31:0] _T_678; // @[Reg.scala 19:20:@427.4]
  reg [31:0] _RAND_12;
  wire [31:0] _GEN_12; // @[Reg.scala 20:19:@428.4]
  reg [31:0] _T_682; // @[Reg.scala 19:20:@433.4]
  reg [31:0] _RAND_13;
  wire [31:0] _GEN_13; // @[Reg.scala 20:19:@434.4]
  reg [31:0] _T_686; // @[Reg.scala 19:20:@439.4]
  reg [31:0] _RAND_14;
  wire [31:0] _GEN_14; // @[Reg.scala 20:19:@440.4]
  reg  _T_690; // @[Reg.scala 19:20:@445.4]
  reg [31:0] _RAND_15;
  wire  _GEN_15; // @[Reg.scala 20:19:@446.4]
  wire  _T_691; // @[NV_NVDLA_CDMA_dual_reg.scala 264:53:@450.4]
  reg  _T_694; // @[Reg.scala 19:20:@451.4]
  reg [31:0] _RAND_16;
  wire  _GEN_16; // @[Reg.scala 20:19:@452.4]
  reg  _T_698; // @[Reg.scala 19:20:@457.4]
  reg [31:0] _RAND_17;
  wire  _GEN_17; // @[Reg.scala 20:19:@458.4]
  reg  _T_702; // @[Reg.scala 19:20:@463.4]
  reg [31:0] _RAND_18;
  wire  _GEN_18; // @[Reg.scala 20:19:@464.4]
  wire [5:0] _T_703; // @[NV_NVDLA_CDMA_dual_reg.scala 270:54:@468.4]
  reg [5:0] _T_706; // @[Reg.scala 19:20:@469.4]
  reg [31:0] _RAND_19;
  wire [5:0] _GEN_19; // @[Reg.scala 20:19:@470.4]
  reg  _T_710; // @[Reg.scala 19:20:@475.4]
  reg [31:0] _RAND_20;
  wire  _GEN_20; // @[Reg.scala 20:19:@476.4]
  wire  _T_711; // @[NV_NVDLA_CDMA_dual_reg.scala 274:61:@480.4]
  reg  _T_714; // @[Reg.scala 19:20:@481.4]
  reg [31:0] _RAND_21;
  wire  _GEN_21; // @[Reg.scala 20:19:@482.4]
  wire [12:0] _T_715; // @[NV_NVDLA_CDMA_dual_reg.scala 276:55:@486.4]
  reg [12:0] _T_718; // @[Reg.scala 19:20:@487.4]
  reg [31:0] _RAND_22;
  wire [12:0] _GEN_22; // @[Reg.scala 20:19:@488.4]
  wire [12:0] _T_719; // @[NV_NVDLA_CDMA_dual_reg.scala 278:54:@492.4]
  reg [12:0] _T_722; // @[Reg.scala 19:20:@493.4]
  reg [31:0] _RAND_23;
  wire [12:0] _GEN_23; // @[Reg.scala 20:19:@494.4]
  reg [12:0] _T_726; // @[Reg.scala 19:20:@499.4]
  reg [31:0] _RAND_24;
  wire [12:0] _GEN_24; // @[Reg.scala 20:19:@500.4]
  reg [12:0] _T_730; // @[Reg.scala 19:20:@505.4]
  reg [31:0] _RAND_25;
  wire [12:0] _GEN_25; // @[Reg.scala 20:19:@506.4]
  reg [12:0] _T_734; // @[Reg.scala 19:20:@511.4]
  reg [31:0] _RAND_26;
  wire [12:0] _GEN_26; // @[Reg.scala 20:19:@512.4]
  wire [13:0] _T_735; // @[NV_NVDLA_CDMA_dual_reg.scala 286:49:@516.4]
  reg [13:0] _T_738; // @[Reg.scala 19:20:@517.4]
  reg [31:0] _RAND_27;
  wire [13:0] _GEN_27; // @[Reg.scala 20:19:@518.4]
  wire [11:0] _T_739; // @[NV_NVDLA_CDMA_dual_reg.scala 288:48:@522.4]
  reg [11:0] _T_742; // @[Reg.scala 19:20:@523.4]
  reg [31:0] _RAND_28;
  wire [11:0] _GEN_28; // @[Reg.scala 20:19:@524.4]
  reg [31:0] _T_746; // @[Reg.scala 19:20:@529.4]
  reg [31:0] _RAND_29;
  wire [31:0] _GEN_29; // @[Reg.scala 20:19:@530.4]
  reg [31:0] _T_750; // @[Reg.scala 19:20:@535.4]
  reg [31:0] _RAND_30;
  wire [31:0] _GEN_30; // @[Reg.scala 20:19:@536.4]
  reg  _T_754; // @[Reg.scala 19:20:@541.4]
  reg [31:0] _RAND_31;
  wire  _GEN_31; // @[Reg.scala 20:19:@542.4]
  wire [15:0] _T_755; // @[NV_NVDLA_CDMA_dual_reg.scala 296:49:@546.4]
  reg [15:0] _T_758; // @[Reg.scala 19:20:@547.4]
  reg [31:0] _RAND_32;
  wire [15:0] _GEN_32; // @[Reg.scala 20:19:@548.4]
  reg [15:0] _T_762; // @[Reg.scala 19:20:@553.4]
  reg [31:0] _RAND_33;
  wire [15:0] _GEN_33; // @[Reg.scala 20:19:@554.4]
  reg [15:0] _T_766; // @[Reg.scala 19:20:@559.4]
  reg [31:0] _RAND_34;
  wire [15:0] _GEN_34; // @[Reg.scala 20:19:@560.4]
  reg [15:0] _T_770; // @[Reg.scala 19:20:@565.4]
  reg [31:0] _RAND_35;
  wire [15:0] _GEN_35; // @[Reg.scala 20:19:@566.4]
  reg  _T_774; // @[Reg.scala 19:20:@571.4]
  reg [31:0] _RAND_36;
  wire  _GEN_36; // @[Reg.scala 20:19:@572.4]
  reg  _T_778; // @[Reg.scala 19:20:@577.4]
  reg [31:0] _RAND_37;
  wire  _GEN_37; // @[Reg.scala 20:19:@578.4]
  wire [1:0] _T_779; // @[NV_NVDLA_CDMA_dual_reg.scala 308:54:@582.4]
  reg [1:0] _T_782; // @[Reg.scala 19:20:@583.4]
  reg [31:0] _RAND_38;
  wire [1:0] _GEN_38; // @[Reg.scala 20:19:@584.4]
  wire [1:0] _T_783; // @[NV_NVDLA_CDMA_dual_reg.scala 310:56:@588.4]
  reg [1:0] _T_786; // @[Reg.scala 19:20:@589.4]
  reg [31:0] _RAND_39;
  wire [1:0] _GEN_39; // @[Reg.scala 20:19:@590.4]
  wire  _T_787; // @[NV_NVDLA_CDMA_dual_reg.scala 312:55:@594.4]
  reg  _T_790; // @[Reg.scala 19:20:@595.4]
  reg [31:0] _RAND_40;
  wire  _GEN_40; // @[Reg.scala 20:19:@596.4]
  wire  _T_791; // @[NV_NVDLA_CDMA_dual_reg.scala 314:57:@600.4]
  reg  _T_794; // @[Reg.scala 19:20:@601.4]
  reg [31:0] _RAND_41;
  wire  _GEN_41; // @[Reg.scala 20:19:@602.4]
  reg  _T_798; // @[Reg.scala 19:20:@607.4]
  reg [31:0] _RAND_42;
  wire  _GEN_42; // @[Reg.scala 20:19:@608.4]
  reg  _T_802; // @[Reg.scala 19:20:@613.4]
  reg [31:0] _RAND_43;
  wire  _GEN_43; // @[Reg.scala 20:19:@614.4]
  reg  _T_806; // @[Reg.scala 19:20:@619.4]
  reg [31:0] _RAND_44;
  wire  _GEN_44; // @[Reg.scala 20:19:@620.4]
  reg [4:0] _T_810; // @[Reg.scala 19:20:@625.4]
  reg [31:0] _RAND_45;
  wire [4:0] _GEN_45; // @[Reg.scala 20:19:@626.4]
  reg [2:0] _T_814; // @[Reg.scala 19:20:@631.4]
  reg [31:0] _RAND_46;
  wire [2:0] _GEN_46; // @[Reg.scala 20:19:@632.4]
  wire [9:0] _T_815; // @[NV_NVDLA_CDMA_dual_reg.scala 326:54:@636.4]
  reg [9:0] _T_818; // @[Reg.scala 19:20:@637.4]
  reg [31:0] _RAND_47;
  wire [9:0] _GEN_47; // @[Reg.scala 20:19:@638.4]
  wire [9:0] _T_819; // @[NV_NVDLA_CDMA_dual_reg.scala 328:57:@642.4]
  reg [9:0] _T_822; // @[Reg.scala 19:20:@643.4]
  reg [31:0] _RAND_48;
  wire [9:0] _GEN_48; // @[Reg.scala 20:19:@644.4]
  reg [2:0] _T_826; // @[Reg.scala 19:20:@649.4]
  reg [31:0] _RAND_49;
  wire [2:0] _GEN_49; // @[Reg.scala 20:19:@650.4]
  reg [4:0] _T_830; // @[Reg.scala 19:20:@655.4]
  reg [31:0] _RAND_50;
  wire [4:0] _GEN_50; // @[Reg.scala 20:19:@656.4]
  reg [31:0] _T_834; // @[Reg.scala 19:20:@661.4]
  reg [31:0] _RAND_51;
  wire [31:0] _GEN_51; // @[Reg.scala 20:19:@662.4]
  reg [31:0] _T_838; // @[Reg.scala 19:20:@667.4]
  reg [31:0] _RAND_52;
  wire [31:0] _GEN_52; // @[Reg.scala 20:19:@668.4]
  reg [31:0] _T_842; // @[Reg.scala 19:20:@673.4]
  reg [31:0] _RAND_53;
  wire [31:0] _GEN_53; // @[Reg.scala 20:19:@674.4]
  reg [31:0] _T_846; // @[Reg.scala 19:20:@679.4]
  reg [31:0] _RAND_54;
  wire [31:0] _GEN_54; // @[Reg.scala 20:19:@680.4]
  reg  _T_850; // @[Reg.scala 19:20:@685.4]
  reg [31:0] _RAND_55;
  wire  _GEN_55; // @[Reg.scala 20:19:@686.4]
  reg  _T_854; // @[Reg.scala 19:20:@691.4]
  reg [31:0] _RAND_56;
  wire  _GEN_56; // @[Reg.scala 20:19:@692.4]
  wire [17:0] _T_855; // @[NV_NVDLA_CDMA_dual_reg.scala 346:57:@696.4]
  reg [17:0] _T_858; // @[Reg.scala 19:20:@697.4]
  reg [31:0] _RAND_57;
  wire [17:0] _GEN_57; // @[Reg.scala 20:19:@698.4]
  reg [12:0] _T_862; // @[Reg.scala 19:20:@703.4]
  reg [31:0] _RAND_58;
  wire [12:0] _GEN_58; // @[Reg.scala 20:19:@704.4]
  reg [31:0] _T_866; // @[Reg.scala 19:20:@709.4]
  reg [31:0] _RAND_59;
  wire [31:0] _GEN_59; // @[Reg.scala 20:19:@710.4]
  reg [31:0] _T_870; // @[Reg.scala 19:20:@715.4]
  reg [31:0] _RAND_60;
  wire [31:0] _GEN_60; // @[Reg.scala 20:19:@716.4]
  reg [31:0] _T_874; // @[Reg.scala 19:20:@721.4]
  reg [31:0] _RAND_61;
  wire [31:0] _GEN_61; // @[Reg.scala 20:19:@722.4]
  reg [31:0] _T_878; // @[Reg.scala 19:20:@727.4]
  reg [31:0] _RAND_62;
  wire [31:0] _GEN_62; // @[Reg.scala 20:19:@728.4]
  wire [27:0] _T_879; // @[NV_NVDLA_CDMA_dual_reg.scala 358:51:@732.4]
  reg [27:0] _T_882; // @[Reg.scala 19:20:@733.4]
  reg [31:0] _RAND_63;
  wire [27:0] _GEN_63; // @[Reg.scala 20:19:@734.4]
  wire [5:0] _T_883; // @[NV_NVDLA_CDMA_dual_reg.scala 360:52:@738.4]
  reg [5:0] _T_886; // @[Reg.scala 19:20:@739.4]
  reg [31:0] _RAND_64;
  wire [5:0] _GEN_64; // @[Reg.scala 20:19:@740.4]
  reg [4:0] _T_890; // @[Reg.scala 19:20:@745.4]
  reg [31:0] _RAND_65;
  wire [4:0] _GEN_65; // @[Reg.scala 20:19:@746.4]
  reg [5:0] _T_894; // @[Reg.scala 19:20:@751.4]
  reg [31:0] _RAND_66;
  wire [5:0] _GEN_66; // @[Reg.scala 20:19:@752.4]
  reg [4:0] _T_898; // @[Reg.scala 19:20:@757.4]
  reg [31:0] _RAND_67;
  wire [4:0] _GEN_67; // @[Reg.scala 20:19:@758.4]
  reg [15:0] _T_902; // @[Reg.scala 19:20:@763.4]
  reg [31:0] _RAND_68;
  wire [15:0] _GEN_68; // @[Reg.scala 20:19:@764.4]
  assign _GEN_69 = {{20'd0}, io_reg_offset}; // @[NV_NVDLA_CDMA_dual_reg.scala 54:51:@59.4]
  assign _T_174 = _GEN_69 == 32'hbc; // @[NV_NVDLA_CDMA_dual_reg.scala 54:51:@59.4]
  assign _T_175 = _T_174 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 54:75:@60.4]
  assign _T_177 = _GEN_69 == 32'h58; // @[NV_NVDLA_CDMA_dual_reg.scala 55:59:@61.4]
  assign _T_178 = _T_177 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 55:83:@62.4]
  assign _T_180 = _GEN_69 == 32'h5c; // @[NV_NVDLA_CDMA_dual_reg.scala 56:59:@63.4]
  assign _T_181 = _T_180 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 56:83:@64.4]
  assign _T_183 = _GEN_69 == 32'hb0; // @[NV_NVDLA_CDMA_dual_reg.scala 57:58:@65.4]
  assign _T_184 = _T_183 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 57:82:@66.4]
  assign _T_186 = _GEN_69 == 32'ha4; // @[NV_NVDLA_CDMA_dual_reg.scala 58:54:@67.4]
  assign _T_187 = _T_186 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 58:78:@68.4]
  assign _T_189 = _GEN_69 == 32'ha8; // @[NV_NVDLA_CDMA_dual_reg.scala 59:57:@69.4]
  assign _T_190 = _T_189 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 59:81:@70.4]
  assign _T_192 = _GEN_69 == 32'hac; // @[NV_NVDLA_CDMA_dual_reg.scala 60:56:@71.4]
  assign _T_193 = _T_192 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 60:80:@72.4]
  assign _T_195 = _GEN_69 == 32'he8; // @[NV_NVDLA_CDMA_dual_reg.scala 61:50:@73.4]
  assign _T_196 = _T_195 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 61:74:@74.4]
  assign _T_198 = _GEN_69 == 32'h30; // @[NV_NVDLA_CDMA_dual_reg.scala 62:63:@75.4]
  assign _T_199 = _T_198 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 62:87:@76.4]
  assign _T_201 = _GEN_69 == 32'h38; // @[NV_NVDLA_CDMA_dual_reg.scala 63:63:@77.4]
  assign _T_202 = _T_201 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 63:87:@78.4]
  assign _T_204 = _GEN_69 == 32'h34; // @[NV_NVDLA_CDMA_dual_reg.scala 64:62:@79.4]
  assign _T_205 = _T_204 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 64:86:@80.4]
  assign _T_207 = _GEN_69 == 32'h3c; // @[NV_NVDLA_CDMA_dual_reg.scala 65:62:@81.4]
  assign _T_208 = _T_207 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 65:86:@82.4]
  assign _T_210 = _GEN_69 == 32'h4c; // @[NV_NVDLA_CDMA_dual_reg.scala 66:55:@83.4]
  assign _T_211 = _T_210 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 66:79:@84.4]
  assign _T_213 = _GEN_69 == 32'h2c; // @[NV_NVDLA_CDMA_dual_reg.scala 67:60:@85.4]
  assign _T_214 = _T_213 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 67:84:@86.4]
  assign _T_216 = _GEN_69 == 32'h18; // @[NV_NVDLA_CDMA_dual_reg.scala 68:60:@87.4]
  assign _T_217 = _T_216 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 68:84:@88.4]
  assign _T_219 = _GEN_69 == 32'h1c; // @[NV_NVDLA_CDMA_dual_reg.scala 69:60:@89.4]
  assign _T_220 = _T_219 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 69:84:@90.4]
  assign _T_222 = _GEN_69 == 32'h20; // @[NV_NVDLA_CDMA_dual_reg.scala 70:60:@91.4]
  assign _T_223 = _T_222 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 70:84:@92.4]
  assign _T_225 = _GEN_69 == 32'h24; // @[NV_NVDLA_CDMA_dual_reg.scala 71:64:@93.4]
  assign _T_226 = _T_225 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 71:88:@94.4]
  assign _T_228 = _GEN_69 == 32'h60; // @[NV_NVDLA_CDMA_dual_reg.scala 72:62:@95.4]
  assign _T_229 = _T_228 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 72:86:@96.4]
  assign _T_231 = _GEN_69 == 32'h64; // @[NV_NVDLA_CDMA_dual_reg.scala 73:58:@97.4]
  assign _T_232 = _T_231 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 73:82:@98.4]
  assign _T_240 = _GEN_69 == 32'h40; // @[NV_NVDLA_CDMA_dual_reg.scala 76:58:@103.4]
  assign _T_241 = _T_240 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 76:82:@104.4]
  assign _T_243 = _GEN_69 == 32'h44; // @[NV_NVDLA_CDMA_dual_reg.scala 77:61:@105.4]
  assign _T_244 = _T_243 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 77:85:@106.4]
  assign _T_246 = _GEN_69 == 32'h98; // @[NV_NVDLA_CDMA_dual_reg.scala 78:58:@107.4]
  assign _T_247 = _T_246 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 78:82:@108.4]
  assign _T_249 = _GEN_69 == 32'h9c; // @[NV_NVDLA_CDMA_dual_reg.scala 79:60:@109.4]
  assign _T_250 = _T_249 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 79:84:@110.4]
  assign _T_252 = _GEN_69 == 32'ha0; // @[NV_NVDLA_CDMA_dual_reg.scala 80:60:@111.4]
  assign _T_253 = _T_252 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 80:84:@112.4]
  assign _T_255 = _GEN_69 == 32'h14; // @[NV_NVDLA_CDMA_dual_reg.scala 81:55:@113.4]
  assign _T_256 = _T_255 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 81:79:@114.4]
  assign _T_258 = _GEN_69 == 32'hc0; // @[NV_NVDLA_CDMA_dual_reg.scala 82:64:@115.4]
  assign _T_259 = _T_258 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 82:88:@116.4]
  assign _T_267 = _GEN_69 == 32'h10; // @[NV_NVDLA_CDMA_dual_reg.scala 85:56:@121.4]
  assign _T_276 = _GEN_69 == 32'hd4; // @[NV_NVDLA_CDMA_dual_reg.scala 88:58:@127.4]
  assign _T_277 = _T_276 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 88:82:@128.4]
  assign _T_285 = _GEN_69 == 32'h28; // @[NV_NVDLA_CDMA_dual_reg.scala 91:59:@133.4]
  assign _T_286 = _T_285 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 91:83:@134.4]
  assign _T_288 = _GEN_69 == 32'h50; // @[NV_NVDLA_CDMA_dual_reg.scala 92:61:@135.4]
  assign _T_289 = _T_288 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 92:85:@136.4]
  assign _T_291 = _GEN_69 == 32'h54; // @[NV_NVDLA_CDMA_dual_reg.scala 93:61:@137.4]
  assign _T_292 = _T_291 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 93:85:@138.4]
  assign _T_294 = _GEN_69 == 32'h48; // @[NV_NVDLA_CDMA_dual_reg.scala 94:58:@139.4]
  assign _T_295 = _T_294 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 94:82:@140.4]
  assign _T_297 = _GEN_69 == 32'h78; // @[NV_NVDLA_CDMA_dual_reg.scala 95:63:@141.4]
  assign _T_298 = _T_297 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 95:87:@142.4]
  assign _T_300 = _GEN_69 == 32'h7c; // @[NV_NVDLA_CDMA_dual_reg.scala 96:62:@143.4]
  assign _T_301 = _T_300 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 96:86:@144.4]
  assign _T_303 = _GEN_69 == 32'h80; // @[NV_NVDLA_CDMA_dual_reg.scala 97:59:@145.4]
  assign _T_304 = _T_303 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 97:83:@146.4]
  assign _T_306 = _GEN_69 == 32'h68; // @[NV_NVDLA_CDMA_dual_reg.scala 98:60:@147.4]
  assign _T_307 = _T_306 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 98:84:@148.4]
  assign _T_309 = _GEN_69 == 32'h74; // @[NV_NVDLA_CDMA_dual_reg.scala 99:62:@149.4]
  assign _T_310 = _T_309 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 99:86:@150.4]
  assign _T_312 = _GEN_69 == 32'h6c; // @[NV_NVDLA_CDMA_dual_reg.scala 100:60:@151.4]
  assign _T_313 = _T_312 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 100:84:@152.4]
  assign _T_315 = _GEN_69 == 32'h70; // @[NV_NVDLA_CDMA_dual_reg.scala 101:60:@153.4]
  assign _T_316 = _T_315 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 101:84:@154.4]
  assign _T_318 = _GEN_69 == 32'h84; // @[NV_NVDLA_CDMA_dual_reg.scala 102:60:@155.4]
  assign _T_319 = _T_318 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 102:84:@156.4]
  assign _T_321 = _GEN_69 == 32'h88; // @[NV_NVDLA_CDMA_dual_reg.scala 103:59:@157.4]
  assign _T_322 = _T_321 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 103:83:@158.4]
  assign _T_324 = _GEN_69 == 32'h8c; // @[NV_NVDLA_CDMA_dual_reg.scala 104:60:@159.4]
  assign _T_325 = _T_324 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 104:84:@160.4]
  assign _T_327 = _GEN_69 == 32'h90; // @[NV_NVDLA_CDMA_dual_reg.scala 105:59:@161.4]
  assign _T_328 = _T_327 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 105:83:@162.4]
  assign _T_330 = _GEN_69 == 32'h94; // @[NV_NVDLA_CDMA_dual_reg.scala 106:56:@163.4]
  assign _T_331 = _T_330 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 106:80:@164.4]
  assign _T_333 = _GEN_69 == 32'hb4; // @[NV_NVDLA_CDMA_dual_reg.scala 107:59:@165.4]
  assign _T_334 = _T_333 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 107:83:@166.4]
  assign _T_336 = _GEN_69 == 32'hb8; // @[NV_NVDLA_CDMA_dual_reg.scala 108:65:@167.4]
  assign _T_337 = _T_336 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 108:89:@168.4]
  assign _T_344 = {11'h0,io_field_weight_bank,11'h0,io_field_data_bank}; // @[Cat.scala 30:58:@172.4]
  assign _T_347 = {27'h0,io_field_batches}; // @[Cat.scala 30:58:@173.4]
  assign _T_354 = {13'h0,io_field_conv_y_stride,13'h0,io_field_conv_x_stride}; // @[Cat.scala 30:58:@176.4]
  assign _T_360 = {22'h0,io_field_cvt_truncate,3'h0,io_field_cvt_en}; // @[Cat.scala 30:58:@179.4]
  assign _T_363 = {16'h0,io_field_cvt_offset}; // @[Cat.scala 30:58:@180.4]
  assign _T_366 = {16'h0,io_field_cvt_scale}; // @[Cat.scala 30:58:@181.4]
  assign _T_377 = {15'h0,io_field_surf_packed,15'h0,io_field_line_packed}; // @[Cat.scala 30:58:@184.4]
  assign _T_380 = {31'h0,io_field_datain_ram_type}; // @[Cat.scala 30:58:@185.4]
  assign _T_392 = {11'h0,io_field_pixel_sign_override,3'h0,io_field_pixel_mapping,2'h0,io_field_pixel_format,7'h0,io_field_datain_format}; // @[Cat.scala 30:58:@192.4]
  assign _T_398 = {3'h0,io_field_datain_height,3'h0,io_field_datain_width}; // @[Cat.scala 30:58:@195.4]
  assign _T_401 = {19'h0,io_field_datain_channel}; // @[Cat.scala 30:58:@196.4]
  assign _T_407 = {3'h0,io_field_datain_height_ext,3'h0,io_field_datain_width_ext}; // @[Cat.scala 30:58:@199.4]
  assign _T_410 = {18'h0,io_field_entries}; // @[Cat.scala 30:58:@200.4]
  assign _T_413 = {20'h0,io_field_grains}; // @[Cat.scala 30:58:@201.4]
  assign _T_420 = {31'h0,io_field_mean_format}; // @[Cat.scala 30:58:@202.4]
  assign _T_422 = {io_field_mean_gu,io_field_mean_ry}; // @[Cat.scala 30:58:@203.4]
  assign _T_424 = {io_field_mean_ax,io_field_mean_bv}; // @[Cat.scala 30:58:@204.4]
  assign _T_438 = {io_field_data_reuse,2'h0,io_field_proc_precision,2'h0,io_field_in_precision,7'h0,io_field_conv_mode}; // @[Cat.scala 30:58:@210.4]
  assign _T_445 = {3'h0,io_field_skip_weight_rls,3'h0,io_field_skip_data_rls,3'h0,io_field_weight_reuse,3'h0,_T_438}; // @[Cat.scala 30:58:@217.4]
  assign _T_448 = {31'h0,io_field_nan_to_zero}; // @[Cat.scala 30:58:@218.4]
  assign _T_453 = {31'h0,io_op_en}; // @[Cat.scala 30:58:@219.4]
  assign _T_458 = {31'h0,io_field_dma_en}; // @[Cat.scala 30:58:@220.4]
  assign _T_466 = {13'h0,io_field_pixel_y_offset,11'h0,io_field_pixel_x_offset}; // @[Cat.scala 30:58:@223.4]
  assign _T_472 = {6'h0,io_field_rsv_per_uv_line,6'h0,io_field_rsv_per_line}; // @[Cat.scala 30:58:@226.4]
  assign _T_478 = {11'h0,io_field_rsv_y_index,13'h0,io_field_rsv_height}; // @[Cat.scala 30:58:@229.4]
  assign _T_485 = {31'h0,io_field_weight_format}; // @[Cat.scala 30:58:@230.4]
  assign _T_488 = {31'h0,io_field_weight_ram_type}; // @[Cat.scala 30:58:@231.4]
  assign _T_491 = {14'h0,io_field_byte_per_kernel}; // @[Cat.scala 30:58:@232.4]
  assign _T_494 = {19'h0,io_field_weight_kernel}; // @[Cat.scala 30:58:@233.4]
  assign _T_501 = {4'h0,io_field_wmb_bytes}; // @[Cat.scala 30:58:@234.4]
  assign _T_513 = {2'h0,io_field_pad_bottom,3'h0,io_field_pad_top,2'h0,io_field_pad_right,3'h0,io_field_pad_left}; // @[Cat.scala 30:58:@241.4]
  assign _T_516 = {16'h0,io_field_pad_value}; // @[Cat.scala 30:58:@242.4]
  assign _T_517 = 32'hb8 == _GEN_69; // @[Mux.scala 46:19:@243.4]
  assign _T_518 = _T_517 ? _T_516 : 32'h0; // @[Mux.scala 46:16:@244.4]
  assign _T_519 = 32'hb4 == _GEN_69; // @[Mux.scala 46:19:@245.4]
  assign _T_520 = _T_519 ? _T_513 : _T_518; // @[Mux.scala 46:16:@246.4]
  assign _T_521 = 32'h94 == _GEN_69; // @[Mux.scala 46:19:@247.4]
  assign _T_522 = _T_521 ? _T_501 : _T_520; // @[Mux.scala 46:16:@248.4]
  assign _T_523 = 32'h90 == _GEN_69; // @[Mux.scala 46:19:@249.4]
  assign _T_524 = _T_523 ? io_field_wmb_addr_low : _T_522; // @[Mux.scala 46:16:@250.4]
  assign _T_525 = 32'h8c == _GEN_69; // @[Mux.scala 46:19:@251.4]
  assign _T_526 = _T_525 ? io_field_wmb_addr_high : _T_524; // @[Mux.scala 46:16:@252.4]
  assign _T_527 = 32'h88 == _GEN_69; // @[Mux.scala 46:19:@253.4]
  assign _T_528 = _T_527 ? io_field_wgs_addr_low : _T_526; // @[Mux.scala 46:16:@254.4]
  assign _T_529 = 32'h84 == _GEN_69; // @[Mux.scala 46:19:@255.4]
  assign _T_530 = _T_529 ? io_field_wgs_addr_high : _T_528; // @[Mux.scala 46:16:@256.4]
  assign _T_531 = 32'h70 == _GEN_69; // @[Mux.scala 46:19:@257.4]
  assign _T_532 = _T_531 ? _T_494 : _T_530; // @[Mux.scala 46:16:@258.4]
  assign _T_533 = 32'h6c == _GEN_69; // @[Mux.scala 46:19:@259.4]
  assign _T_534 = _T_533 ? _T_491 : _T_532; // @[Mux.scala 46:16:@260.4]
  assign _T_535 = 32'h74 == _GEN_69; // @[Mux.scala 46:19:@261.4]
  assign _T_536 = _T_535 ? _T_488 : _T_534; // @[Mux.scala 46:16:@262.4]
  assign _T_537 = 32'h68 == _GEN_69; // @[Mux.scala 46:19:@263.4]
  assign _T_538 = _T_537 ? _T_485 : _T_536; // @[Mux.scala 46:16:@264.4]
  assign _T_539 = 32'h80 == _GEN_69; // @[Mux.scala 46:19:@265.4]
  assign _T_540 = _T_539 ? io_field_weight_bytes : _T_538; // @[Mux.scala 46:16:@266.4]
  assign _T_541 = 32'h7c == _GEN_69; // @[Mux.scala 46:19:@267.4]
  assign _T_542 = _T_541 ? io_field_weight_addr_low : _T_540; // @[Mux.scala 46:16:@268.4]
  assign _T_543 = 32'h78 == _GEN_69; // @[Mux.scala 46:19:@269.4]
  assign _T_544 = _T_543 ? io_field_weight_addr_high : _T_542; // @[Mux.scala 46:16:@270.4]
  assign _T_545 = 32'h48 == _GEN_69; // @[Mux.scala 46:19:@271.4]
  assign _T_546 = _T_545 ? io_field_surf_stride : _T_544; // @[Mux.scala 46:16:@272.4]
  assign _T_547 = 32'h54 == _GEN_69; // @[Mux.scala 46:19:@273.4]
  assign _T_548 = _T_547 ? _T_478 : _T_546; // @[Mux.scala 46:16:@274.4]
  assign _T_549 = 32'h50 == _GEN_69; // @[Mux.scala 46:19:@275.4]
  assign _T_550 = _T_549 ? _T_472 : _T_548; // @[Mux.scala 46:16:@276.4]
  assign _T_551 = 32'h28 == _GEN_69; // @[Mux.scala 46:19:@277.4]
  assign _T_552 = _T_551 ? _T_466 : _T_550; // @[Mux.scala 46:16:@278.4]
  assign _T_553 = 32'hdc == _GEN_69; // @[Mux.scala 46:19:@279.4]
  assign _T_554 = _T_553 ? io_wt_rd_stall : _T_552; // @[Mux.scala 46:16:@280.4]
  assign _T_555 = 32'he4 == _GEN_69; // @[Mux.scala 46:19:@281.4]
  assign _T_556 = _T_555 ? io_wt_rd_latency : _T_554; // @[Mux.scala 46:16:@282.4]
  assign _T_557 = 32'hd4 == _GEN_69; // @[Mux.scala 46:19:@283.4]
  assign _T_558 = _T_557 ? _T_458 : _T_556; // @[Mux.scala 46:16:@284.4]
  assign _T_559 = 32'hd8 == _GEN_69; // @[Mux.scala 46:19:@285.4]
  assign _T_560 = _T_559 ? io_dat_rd_stall : _T_558; // @[Mux.scala 46:16:@286.4]
  assign _T_561 = 32'he0 == _GEN_69; // @[Mux.scala 46:19:@287.4]
  assign _T_562 = _T_561 ? io_dat_rd_latency : _T_560; // @[Mux.scala 46:16:@288.4]
  assign _T_563 = 32'h10 == _GEN_69; // @[Mux.scala 46:19:@289.4]
  assign _T_564 = _T_563 ? _T_453 : _T_562; // @[Mux.scala 46:16:@290.4]
  assign _T_565 = 32'hc8 == _GEN_69; // @[Mux.scala 46:19:@291.4]
  assign _T_566 = _T_565 ? io_nan_weight_num : _T_564; // @[Mux.scala 46:16:@292.4]
  assign _T_567 = 32'hc4 == _GEN_69; // @[Mux.scala 46:19:@293.4]
  assign _T_568 = _T_567 ? io_nan_data_num : _T_566; // @[Mux.scala 46:16:@294.4]
  assign _T_569 = 32'hc0 == _GEN_69; // @[Mux.scala 46:19:@295.4]
  assign _T_570 = _T_569 ? _T_448 : _T_568; // @[Mux.scala 46:16:@296.4]
  assign _T_571 = 32'h14 == _GEN_69; // @[Mux.scala 46:19:@297.4]
  assign _T_572 = _T_571 ? _T_445 : _T_570; // @[Mux.scala 46:16:@298.4]
  assign _T_573 = 32'ha0 == _GEN_69; // @[Mux.scala 46:19:@299.4]
  assign _T_574 = _T_573 ? _T_424 : _T_572; // @[Mux.scala 46:16:@300.4]
  assign _T_575 = 32'h9c == _GEN_69; // @[Mux.scala 46:19:@301.4]
  assign _T_576 = _T_575 ? _T_422 : _T_574; // @[Mux.scala 46:16:@302.4]
  assign _T_577 = 32'h98 == _GEN_69; // @[Mux.scala 46:19:@303.4]
  assign _T_578 = _T_577 ? _T_420 : _T_576; // @[Mux.scala 46:16:@304.4]
  assign _T_579 = 32'h44 == _GEN_69; // @[Mux.scala 46:19:@305.4]
  assign _T_580 = _T_579 ? io_field_uv_line_stride : _T_578; // @[Mux.scala 46:16:@306.4]
  assign _T_581 = 32'h40 == _GEN_69; // @[Mux.scala 46:19:@307.4]
  assign _T_582 = _T_581 ? io_field_line_stride : _T_580; // @[Mux.scala 46:16:@308.4]
  assign _T_583 = 32'hd0 == _GEN_69; // @[Mux.scala 46:19:@309.4]
  assign _T_584 = _T_583 ? io_inf_weight_num : _T_582; // @[Mux.scala 46:16:@310.4]
  assign _T_585 = 32'hcc == _GEN_69; // @[Mux.scala 46:19:@311.4]
  assign _T_586 = _T_585 ? io_inf_data_num : _T_584; // @[Mux.scala 46:16:@312.4]
  assign _T_587 = 32'h64 == _GEN_69; // @[Mux.scala 46:19:@313.4]
  assign _T_588 = _T_587 ? _T_413 : _T_586; // @[Mux.scala 46:16:@314.4]
  assign _T_589 = 32'h60 == _GEN_69; // @[Mux.scala 46:19:@315.4]
  assign _T_590 = _T_589 ? _T_410 : _T_588; // @[Mux.scala 46:16:@316.4]
  assign _T_591 = 32'h24 == _GEN_69; // @[Mux.scala 46:19:@317.4]
  assign _T_592 = _T_591 ? _T_407 : _T_590; // @[Mux.scala 46:16:@318.4]
  assign _T_593 = 32'h20 == _GEN_69; // @[Mux.scala 46:19:@319.4]
  assign _T_594 = _T_593 ? _T_401 : _T_592; // @[Mux.scala 46:16:@320.4]
  assign _T_595 = 32'h1c == _GEN_69; // @[Mux.scala 46:19:@321.4]
  assign _T_596 = _T_595 ? _T_398 : _T_594; // @[Mux.scala 46:16:@322.4]
  assign _T_597 = 32'h18 == _GEN_69; // @[Mux.scala 46:19:@323.4]
  assign _T_598 = _T_597 ? _T_392 : _T_596; // @[Mux.scala 46:16:@324.4]
  assign _T_599 = 32'h2c == _GEN_69; // @[Mux.scala 46:19:@325.4]
  assign _T_600 = _T_599 ? _T_380 : _T_598; // @[Mux.scala 46:16:@326.4]
  assign _T_601 = 32'h4c == _GEN_69; // @[Mux.scala 46:19:@327.4]
  assign _T_602 = _T_601 ? _T_377 : _T_600; // @[Mux.scala 46:16:@328.4]
  assign _T_603 = 32'h3c == _GEN_69; // @[Mux.scala 46:19:@329.4]
  assign _T_604 = _T_603 ? io_field_datain_addr_low_1 : _T_602; // @[Mux.scala 46:16:@330.4]
  assign _T_605 = 32'h34 == _GEN_69; // @[Mux.scala 46:19:@331.4]
  assign _T_606 = _T_605 ? io_field_datain_addr_low_0 : _T_604; // @[Mux.scala 46:16:@332.4]
  assign _T_607 = 32'h38 == _GEN_69; // @[Mux.scala 46:19:@333.4]
  assign _T_608 = _T_607 ? io_field_datain_addr_high_1 : _T_606; // @[Mux.scala 46:16:@334.4]
  assign _T_609 = 32'h30 == _GEN_69; // @[Mux.scala 46:19:@335.4]
  assign _T_610 = _T_609 ? io_field_datain_addr_high_0 : _T_608; // @[Mux.scala 46:16:@336.4]
  assign _T_611 = 32'he8 == _GEN_69; // @[Mux.scala 46:19:@337.4]
  assign _T_612 = _T_611 ? io_field_cya : _T_610; // @[Mux.scala 46:16:@338.4]
  assign _T_613 = 32'hac == _GEN_69; // @[Mux.scala 46:19:@339.4]
  assign _T_614 = _T_613 ? _T_366 : _T_612; // @[Mux.scala 46:16:@340.4]
  assign _T_615 = 32'ha8 == _GEN_69; // @[Mux.scala 46:19:@341.4]
  assign _T_616 = _T_615 ? _T_363 : _T_614; // @[Mux.scala 46:16:@342.4]
  assign _T_617 = 32'ha4 == _GEN_69; // @[Mux.scala 46:19:@343.4]
  assign _T_618 = _T_617 ? _T_360 : _T_616; // @[Mux.scala 46:16:@344.4]
  assign _T_619 = 32'hb0 == _GEN_69; // @[Mux.scala 46:19:@345.4]
  assign _T_620 = _T_619 ? _T_354 : _T_618; // @[Mux.scala 46:16:@346.4]
  assign _T_621 = 32'h5c == _GEN_69; // @[Mux.scala 46:19:@347.4]
  assign _T_622 = _T_621 ? io_field_batch_stride : _T_620; // @[Mux.scala 46:16:@348.4]
  assign _T_623 = 32'h58 == _GEN_69; // @[Mux.scala 46:19:@349.4]
  assign _T_624 = _T_623 ? _T_347 : _T_622; // @[Mux.scala 46:16:@350.4]
  assign _T_625 = 32'hbc == _GEN_69; // @[Mux.scala 46:19:@351.4]
  assign _T_627 = io_reg_wr_data[4:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 232:51:@354.4]
  assign _GEN_0 = _T_175 ? _T_627 : _T_630; // @[Reg.scala 20:19:@356.4]
  assign _T_631 = io_reg_wr_data[20:16]; // @[NV_NVDLA_CDMA_dual_reg.scala 234:53:@360.4]
  assign _GEN_1 = _T_175 ? _T_631 : _T_634; // @[Reg.scala 20:19:@362.4]
  assign _GEN_2 = _T_178 ? _T_627 : _T_638; // @[Reg.scala 20:19:@368.4]
  assign _GEN_3 = _T_181 ? io_reg_wr_data : _T_642; // @[Reg.scala 20:19:@374.4]
  assign _T_643 = io_reg_wr_data[2:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 240:55:@378.4]
  assign _GEN_4 = _T_184 ? _T_643 : _T_646; // @[Reg.scala 20:19:@380.4]
  assign _T_647 = io_reg_wr_data[18:16]; // @[NV_NVDLA_CDMA_dual_reg.scala 242:55:@384.4]
  assign _GEN_5 = _T_184 ? _T_647 : _T_650; // @[Reg.scala 20:19:@386.4]
  assign _T_651 = io_reg_wr_data[0]; // @[NV_NVDLA_CDMA_dual_reg.scala 244:48:@390.4]
  assign _GEN_6 = _T_187 ? _T_651 : _T_654; // @[Reg.scala 20:19:@392.4]
  assign _T_655 = io_reg_wr_data[9:4]; // @[NV_NVDLA_CDMA_dual_reg.scala 246:54:@396.4]
  assign _GEN_7 = _T_187 ? _T_655 : _T_658; // @[Reg.scala 20:19:@398.4]
  assign _T_659 = io_reg_wr_data[15:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 248:52:@402.4]
  assign _GEN_8 = _T_190 ? _T_659 : _T_662; // @[Reg.scala 20:19:@404.4]
  assign _GEN_9 = _T_193 ? _T_659 : _T_666; // @[Reg.scala 20:19:@410.4]
  assign _GEN_10 = _T_196 ? io_reg_wr_data : _T_670; // @[Reg.scala 20:19:@416.4]
  assign _GEN_11 = _T_199 ? io_reg_wr_data : _T_674; // @[Reg.scala 20:19:@422.4]
  assign _GEN_12 = _T_202 ? io_reg_wr_data : _T_678; // @[Reg.scala 20:19:@428.4]
  assign _GEN_13 = _T_205 ? io_reg_wr_data : _T_682; // @[Reg.scala 20:19:@434.4]
  assign _GEN_14 = _T_208 ? io_reg_wr_data : _T_686; // @[Reg.scala 20:19:@440.4]
  assign _GEN_15 = _T_211 ? _T_651 : _T_690; // @[Reg.scala 20:19:@446.4]
  assign _T_691 = io_reg_wr_data[16]; // @[NV_NVDLA_CDMA_dual_reg.scala 264:53:@450.4]
  assign _GEN_16 = _T_211 ? _T_691 : _T_694; // @[Reg.scala 20:19:@452.4]
  assign _GEN_17 = _T_214 ? _T_651 : _T_698; // @[Reg.scala 20:19:@458.4]
  assign _GEN_18 = _T_217 ? _T_651 : _T_702; // @[Reg.scala 20:19:@464.4]
  assign _T_703 = io_reg_wr_data[13:8]; // @[NV_NVDLA_CDMA_dual_reg.scala 270:54:@468.4]
  assign _GEN_19 = _T_217 ? _T_703 : _T_706; // @[Reg.scala 20:19:@470.4]
  assign _GEN_20 = _T_217 ? _T_691 : _T_710; // @[Reg.scala 20:19:@476.4]
  assign _T_711 = io_reg_wr_data[20]; // @[NV_NVDLA_CDMA_dual_reg.scala 274:61:@480.4]
  assign _GEN_21 = _T_217 ? _T_711 : _T_714; // @[Reg.scala 20:19:@482.4]
  assign _T_715 = io_reg_wr_data[28:16]; // @[NV_NVDLA_CDMA_dual_reg.scala 276:55:@486.4]
  assign _GEN_22 = _T_220 ? _T_715 : _T_718; // @[Reg.scala 20:19:@488.4]
  assign _T_719 = io_reg_wr_data[12:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 278:54:@492.4]
  assign _GEN_23 = _T_220 ? _T_719 : _T_722; // @[Reg.scala 20:19:@494.4]
  assign _GEN_24 = _T_223 ? _T_719 : _T_726; // @[Reg.scala 20:19:@500.4]
  assign _GEN_25 = _T_226 ? _T_715 : _T_730; // @[Reg.scala 20:19:@506.4]
  assign _GEN_26 = _T_226 ? _T_719 : _T_734; // @[Reg.scala 20:19:@512.4]
  assign _T_735 = io_reg_wr_data[13:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 286:49:@516.4]
  assign _GEN_27 = _T_229 ? _T_735 : _T_738; // @[Reg.scala 20:19:@518.4]
  assign _T_739 = io_reg_wr_data[11:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 288:48:@522.4]
  assign _GEN_28 = _T_232 ? _T_739 : _T_742; // @[Reg.scala 20:19:@524.4]
  assign _GEN_29 = _T_241 ? io_reg_wr_data : _T_746; // @[Reg.scala 20:19:@530.4]
  assign _GEN_30 = _T_244 ? io_reg_wr_data : _T_750; // @[Reg.scala 20:19:@536.4]
  assign _GEN_31 = _T_247 ? _T_651 : _T_754; // @[Reg.scala 20:19:@542.4]
  assign _T_755 = io_reg_wr_data[31:16]; // @[NV_NVDLA_CDMA_dual_reg.scala 296:49:@546.4]
  assign _GEN_32 = _T_250 ? _T_755 : _T_758; // @[Reg.scala 20:19:@548.4]
  assign _GEN_33 = _T_250 ? _T_659 : _T_762; // @[Reg.scala 20:19:@554.4]
  assign _GEN_34 = _T_253 ? _T_755 : _T_766; // @[Reg.scala 20:19:@560.4]
  assign _GEN_35 = _T_253 ? _T_659 : _T_770; // @[Reg.scala 20:19:@566.4]
  assign _GEN_36 = _T_256 ? _T_651 : _T_774; // @[Reg.scala 20:19:@572.4]
  assign _GEN_37 = _T_256 ? _T_691 : _T_778; // @[Reg.scala 20:19:@578.4]
  assign _T_779 = io_reg_wr_data[9:8]; // @[NV_NVDLA_CDMA_dual_reg.scala 308:54:@582.4]
  assign _GEN_38 = _T_256 ? _T_779 : _T_782; // @[Reg.scala 20:19:@584.4]
  assign _T_783 = io_reg_wr_data[13:12]; // @[NV_NVDLA_CDMA_dual_reg.scala 310:56:@588.4]
  assign _GEN_39 = _T_256 ? _T_783 : _T_786; // @[Reg.scala 20:19:@590.4]
  assign _T_787 = io_reg_wr_data[24]; // @[NV_NVDLA_CDMA_dual_reg.scala 312:55:@594.4]
  assign _GEN_40 = _T_256 ? _T_787 : _T_790; // @[Reg.scala 20:19:@596.4]
  assign _T_791 = io_reg_wr_data[28]; // @[NV_NVDLA_CDMA_dual_reg.scala 314:57:@600.4]
  assign _GEN_41 = _T_256 ? _T_791 : _T_794; // @[Reg.scala 20:19:@602.4]
  assign _GEN_42 = _T_256 ? _T_711 : _T_798; // @[Reg.scala 20:19:@608.4]
  assign _GEN_43 = _T_259 ? _T_651 : _T_802; // @[Reg.scala 20:19:@614.4]
  assign _GEN_44 = _T_277 ? _T_651 : _T_806; // @[Reg.scala 20:19:@620.4]
  assign _GEN_45 = _T_286 ? _T_627 : _T_810; // @[Reg.scala 20:19:@626.4]
  assign _GEN_46 = _T_286 ? _T_647 : _T_814; // @[Reg.scala 20:19:@632.4]
  assign _T_815 = io_reg_wr_data[9:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 326:54:@636.4]
  assign _GEN_47 = _T_289 ? _T_815 : _T_818; // @[Reg.scala 20:19:@638.4]
  assign _T_819 = io_reg_wr_data[25:16]; // @[NV_NVDLA_CDMA_dual_reg.scala 328:57:@642.4]
  assign _GEN_48 = _T_289 ? _T_819 : _T_822; // @[Reg.scala 20:19:@644.4]
  assign _GEN_49 = _T_292 ? _T_643 : _T_826; // @[Reg.scala 20:19:@650.4]
  assign _GEN_50 = _T_292 ? _T_631 : _T_830; // @[Reg.scala 20:19:@656.4]
  assign _GEN_51 = _T_295 ? io_reg_wr_data : _T_834; // @[Reg.scala 20:19:@662.4]
  assign _GEN_52 = _T_298 ? io_reg_wr_data : _T_838; // @[Reg.scala 20:19:@668.4]
  assign _GEN_53 = _T_301 ? io_reg_wr_data : _T_842; // @[Reg.scala 20:19:@674.4]
  assign _GEN_54 = _T_304 ? io_reg_wr_data : _T_846; // @[Reg.scala 20:19:@680.4]
  assign _GEN_55 = _T_307 ? _T_651 : _T_850; // @[Reg.scala 20:19:@686.4]
  assign _GEN_56 = _T_310 ? _T_651 : _T_854; // @[Reg.scala 20:19:@692.4]
  assign _T_855 = io_reg_wr_data[17:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 346:57:@696.4]
  assign _GEN_57 = _T_313 ? _T_855 : _T_858; // @[Reg.scala 20:19:@698.4]
  assign _GEN_58 = _T_316 ? _T_719 : _T_862; // @[Reg.scala 20:19:@704.4]
  assign _GEN_59 = _T_319 ? io_reg_wr_data : _T_866; // @[Reg.scala 20:19:@710.4]
  assign _GEN_60 = _T_322 ? io_reg_wr_data : _T_870; // @[Reg.scala 20:19:@716.4]
  assign _GEN_61 = _T_325 ? io_reg_wr_data : _T_874; // @[Reg.scala 20:19:@722.4]
  assign _GEN_62 = _T_328 ? io_reg_wr_data : _T_878; // @[Reg.scala 20:19:@728.4]
  assign _T_879 = io_reg_wr_data[27:0]; // @[NV_NVDLA_CDMA_dual_reg.scala 358:51:@732.4]
  assign _GEN_63 = _T_331 ? _T_879 : _T_882; // @[Reg.scala 20:19:@734.4]
  assign _T_883 = io_reg_wr_data[29:24]; // @[NV_NVDLA_CDMA_dual_reg.scala 360:52:@738.4]
  assign _GEN_64 = _T_334 ? _T_883 : _T_886; // @[Reg.scala 20:19:@740.4]
  assign _GEN_65 = _T_334 ? _T_627 : _T_890; // @[Reg.scala 20:19:@746.4]
  assign _GEN_66 = _T_334 ? _T_703 : _T_894; // @[Reg.scala 20:19:@752.4]
  assign _GEN_67 = _T_334 ? _T_631 : _T_898; // @[Reg.scala 20:19:@758.4]
  assign _GEN_68 = _T_337 ? _T_659 : _T_902; // @[Reg.scala 20:19:@764.4]
  assign io_reg_rd_data = _T_625 ? _T_344 : _T_624; // @[NV_NVDLA_CDMA_dual_reg.scala 114:20:@353.4]
  assign io_field_data_bank = _T_630; // @[NV_NVDLA_CDMA_dual_reg.scala 232:24:@359.4]
  assign io_field_weight_bank = _T_634; // @[NV_NVDLA_CDMA_dual_reg.scala 234:26:@365.4]
  assign io_field_batches = _T_638; // @[NV_NVDLA_CDMA_dual_reg.scala 236:22:@371.4]
  assign io_field_batch_stride = _T_642; // @[NV_NVDLA_CDMA_dual_reg.scala 238:27:@377.4]
  assign io_field_conv_x_stride = _T_646; // @[NV_NVDLA_CDMA_dual_reg.scala 240:28:@383.4]
  assign io_field_conv_y_stride = _T_650; // @[NV_NVDLA_CDMA_dual_reg.scala 242:28:@389.4]
  assign io_field_cvt_en = _T_654; // @[NV_NVDLA_CDMA_dual_reg.scala 244:21:@395.4]
  assign io_field_cvt_truncate = _T_658; // @[NV_NVDLA_CDMA_dual_reg.scala 246:27:@401.4]
  assign io_field_cvt_offset = _T_662; // @[NV_NVDLA_CDMA_dual_reg.scala 248:25:@407.4]
  assign io_field_cvt_scale = _T_666; // @[NV_NVDLA_CDMA_dual_reg.scala 250:24:@413.4]
  assign io_field_cya = _T_670; // @[NV_NVDLA_CDMA_dual_reg.scala 252:18:@419.4]
  assign io_field_datain_addr_high_0 = _T_674; // @[NV_NVDLA_CDMA_dual_reg.scala 254:33:@425.4]
  assign io_field_datain_addr_high_1 = _T_678; // @[NV_NVDLA_CDMA_dual_reg.scala 256:33:@431.4]
  assign io_field_datain_addr_low_0 = _T_682; // @[NV_NVDLA_CDMA_dual_reg.scala 258:32:@437.4]
  assign io_field_datain_addr_low_1 = _T_686; // @[NV_NVDLA_CDMA_dual_reg.scala 260:32:@443.4]
  assign io_field_line_packed = _T_690; // @[NV_NVDLA_CDMA_dual_reg.scala 262:26:@449.4]
  assign io_field_surf_packed = _T_694; // @[NV_NVDLA_CDMA_dual_reg.scala 264:26:@455.4]
  assign io_field_datain_ram_type = _T_698; // @[NV_NVDLA_CDMA_dual_reg.scala 266:30:@461.4]
  assign io_field_datain_format = _T_702; // @[NV_NVDLA_CDMA_dual_reg.scala 268:28:@467.4]
  assign io_field_pixel_format = _T_706; // @[NV_NVDLA_CDMA_dual_reg.scala 270:27:@473.4]
  assign io_field_pixel_mapping = _T_710; // @[NV_NVDLA_CDMA_dual_reg.scala 272:28:@479.4]
  assign io_field_pixel_sign_override = _T_714; // @[NV_NVDLA_CDMA_dual_reg.scala 274:34:@485.4]
  assign io_field_datain_height = _T_718; // @[NV_NVDLA_CDMA_dual_reg.scala 276:28:@491.4]
  assign io_field_datain_width = _T_722; // @[NV_NVDLA_CDMA_dual_reg.scala 278:27:@497.4]
  assign io_field_datain_channel = _T_726; // @[NV_NVDLA_CDMA_dual_reg.scala 280:29:@503.4]
  assign io_field_datain_height_ext = _T_730; // @[NV_NVDLA_CDMA_dual_reg.scala 282:32:@509.4]
  assign io_field_datain_width_ext = _T_734; // @[NV_NVDLA_CDMA_dual_reg.scala 284:31:@515.4]
  assign io_field_entries = _T_738; // @[NV_NVDLA_CDMA_dual_reg.scala 286:22:@521.4]
  assign io_field_grains = _T_742; // @[NV_NVDLA_CDMA_dual_reg.scala 288:21:@527.4]
  assign io_field_line_stride = _T_746; // @[NV_NVDLA_CDMA_dual_reg.scala 290:26:@533.4]
  assign io_field_uv_line_stride = _T_750; // @[NV_NVDLA_CDMA_dual_reg.scala 292:29:@539.4]
  assign io_field_mean_format = _T_754; // @[NV_NVDLA_CDMA_dual_reg.scala 294:26:@545.4]
  assign io_field_mean_gu = _T_758; // @[NV_NVDLA_CDMA_dual_reg.scala 296:22:@551.4]
  assign io_field_mean_ry = _T_762; // @[NV_NVDLA_CDMA_dual_reg.scala 298:22:@557.4]
  assign io_field_mean_ax = _T_766; // @[NV_NVDLA_CDMA_dual_reg.scala 300:22:@563.4]
  assign io_field_mean_bv = _T_770; // @[NV_NVDLA_CDMA_dual_reg.scala 302:22:@569.4]
  assign io_field_conv_mode = _T_774; // @[NV_NVDLA_CDMA_dual_reg.scala 304:24:@575.4]
  assign io_field_data_reuse = _T_778; // @[NV_NVDLA_CDMA_dual_reg.scala 306:25:@581.4]
  assign io_field_in_precision = _T_782; // @[NV_NVDLA_CDMA_dual_reg.scala 308:27:@587.4]
  assign io_field_proc_precision = _T_786; // @[NV_NVDLA_CDMA_dual_reg.scala 310:29:@593.4]
  assign io_field_skip_data_rls = _T_790; // @[NV_NVDLA_CDMA_dual_reg.scala 312:28:@599.4]
  assign io_field_skip_weight_rls = _T_794; // @[NV_NVDLA_CDMA_dual_reg.scala 314:30:@605.4]
  assign io_field_weight_reuse = _T_798; // @[NV_NVDLA_CDMA_dual_reg.scala 316:27:@611.4]
  assign io_field_nan_to_zero = _T_802; // @[NV_NVDLA_CDMA_dual_reg.scala 318:26:@617.4]
  assign io_field_dma_en = _T_806; // @[NV_NVDLA_CDMA_dual_reg.scala 320:21:@623.4]
  assign io_field_pixel_x_offset = _T_810; // @[NV_NVDLA_CDMA_dual_reg.scala 322:29:@629.4]
  assign io_field_pixel_y_offset = _T_814; // @[NV_NVDLA_CDMA_dual_reg.scala 324:29:@635.4]
  assign io_field_rsv_per_line = _T_818; // @[NV_NVDLA_CDMA_dual_reg.scala 326:27:@641.4]
  assign io_field_rsv_per_uv_line = _T_822; // @[NV_NVDLA_CDMA_dual_reg.scala 328:30:@647.4]
  assign io_field_rsv_height = _T_826; // @[NV_NVDLA_CDMA_dual_reg.scala 330:25:@653.4]
  assign io_field_rsv_y_index = _T_830; // @[NV_NVDLA_CDMA_dual_reg.scala 332:26:@659.4]
  assign io_field_surf_stride = _T_834; // @[NV_NVDLA_CDMA_dual_reg.scala 334:26:@665.4]
  assign io_field_weight_addr_high = _T_838; // @[NV_NVDLA_CDMA_dual_reg.scala 336:31:@671.4]
  assign io_field_weight_addr_low = _T_842; // @[NV_NVDLA_CDMA_dual_reg.scala 338:30:@677.4]
  assign io_field_weight_bytes = _T_846; // @[NV_NVDLA_CDMA_dual_reg.scala 340:27:@683.4]
  assign io_field_weight_format = _T_850; // @[NV_NVDLA_CDMA_dual_reg.scala 342:28:@689.4]
  assign io_field_weight_ram_type = _T_854; // @[NV_NVDLA_CDMA_dual_reg.scala 344:30:@695.4]
  assign io_field_byte_per_kernel = _T_858; // @[NV_NVDLA_CDMA_dual_reg.scala 346:30:@701.4]
  assign io_field_weight_kernel = _T_862; // @[NV_NVDLA_CDMA_dual_reg.scala 348:28:@707.4]
  assign io_field_wgs_addr_high = _T_866; // @[NV_NVDLA_CDMA_dual_reg.scala 350:28:@713.4]
  assign io_field_wgs_addr_low = _T_870; // @[NV_NVDLA_CDMA_dual_reg.scala 352:27:@719.4]
  assign io_field_wmb_addr_high = _T_874; // @[NV_NVDLA_CDMA_dual_reg.scala 354:28:@725.4]
  assign io_field_wmb_addr_low = _T_878; // @[NV_NVDLA_CDMA_dual_reg.scala 356:27:@731.4]
  assign io_field_wmb_bytes = _T_882; // @[NV_NVDLA_CDMA_dual_reg.scala 358:24:@737.4]
  assign io_field_pad_bottom = _T_886; // @[NV_NVDLA_CDMA_dual_reg.scala 360:25:@743.4]
  assign io_field_pad_left = _T_890; // @[NV_NVDLA_CDMA_dual_reg.scala 362:23:@749.4]
  assign io_field_pad_right = _T_894; // @[NV_NVDLA_CDMA_dual_reg.scala 364:24:@755.4]
  assign io_field_pad_top = _T_898; // @[NV_NVDLA_CDMA_dual_reg.scala 366:22:@761.4]
  assign io_field_pad_value = _T_902; // @[NV_NVDLA_CDMA_dual_reg.scala 368:24:@767.4]
  assign io_op_en_trigger = _T_267 & io_reg_wr_en; // @[NV_NVDLA_CDMA_dual_reg.scala 110:22:@169.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_630 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_634 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_638 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_642 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_646 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_650 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_654 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_658 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_662 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_666 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_670 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_674 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_678 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_682 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_686 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_690 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_694 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_698 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_702 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_706 = _RAND_19[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_710 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_714 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_718 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_722 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_726 = _RAND_24[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_730 = _RAND_25[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_734 = _RAND_26[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_738 = _RAND_27[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_742 = _RAND_28[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_746 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_750 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_754 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_758 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_762 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_766 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_770 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_774 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_778 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_782 = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_786 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_790 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_794 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_798 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_802 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_806 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_810 = _RAND_45[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_814 = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_818 = _RAND_47[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_822 = _RAND_48[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_826 = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_830 = _RAND_50[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_834 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_838 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_842 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_846 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_850 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_854 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_858 = _RAND_57[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_862 = _RAND_58[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_866 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_870 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_874 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_878 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_882 = _RAND_63[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_886 = _RAND_64[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_890 = _RAND_65[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_894 = _RAND_66[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_898 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_902 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_630 <= 5'h0;
    end else begin
      if (_T_175) begin
        _T_630 <= _T_627;
      end
    end
    if (reset) begin
      _T_634 <= 5'h0;
    end else begin
      if (_T_175) begin
        _T_634 <= _T_631;
      end
    end
    if (reset) begin
      _T_638 <= 5'h0;
    end else begin
      if (_T_178) begin
        _T_638 <= _T_627;
      end
    end
    if (reset) begin
      _T_642 <= 32'h0;
    end else begin
      if (_T_181) begin
        _T_642 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_646 <= 3'h0;
    end else begin
      if (_T_184) begin
        _T_646 <= _T_643;
      end
    end
    if (reset) begin
      _T_650 <= 3'h0;
    end else begin
      if (_T_184) begin
        _T_650 <= _T_647;
      end
    end
    if (reset) begin
      _T_654 <= 1'h0;
    end else begin
      if (_T_187) begin
        _T_654 <= _T_651;
      end
    end
    if (reset) begin
      _T_658 <= 6'h0;
    end else begin
      if (_T_187) begin
        _T_658 <= _T_655;
      end
    end
    if (reset) begin
      _T_662 <= 16'h0;
    end else begin
      if (_T_190) begin
        _T_662 <= _T_659;
      end
    end
    if (reset) begin
      _T_666 <= 16'h0;
    end else begin
      if (_T_193) begin
        _T_666 <= _T_659;
      end
    end
    if (reset) begin
      _T_670 <= 32'h0;
    end else begin
      if (_T_196) begin
        _T_670 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_674 <= 32'h0;
    end else begin
      if (_T_199) begin
        _T_674 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_678 <= 32'h0;
    end else begin
      if (_T_202) begin
        _T_678 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_682 <= 32'h0;
    end else begin
      if (_T_205) begin
        _T_682 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_686 <= 32'h0;
    end else begin
      if (_T_208) begin
        _T_686 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_690 <= 1'h0;
    end else begin
      if (_T_211) begin
        _T_690 <= _T_651;
      end
    end
    if (reset) begin
      _T_694 <= 1'h0;
    end else begin
      if (_T_211) begin
        _T_694 <= _T_691;
      end
    end
    if (reset) begin
      _T_698 <= 1'h0;
    end else begin
      if (_T_214) begin
        _T_698 <= _T_651;
      end
    end
    if (reset) begin
      _T_702 <= 1'h0;
    end else begin
      if (_T_217) begin
        _T_702 <= _T_651;
      end
    end
    if (reset) begin
      _T_706 <= 6'hc;
    end else begin
      if (_T_217) begin
        _T_706 <= _T_703;
      end
    end
    if (reset) begin
      _T_710 <= 1'h0;
    end else begin
      if (_T_217) begin
        _T_710 <= _T_691;
      end
    end
    if (reset) begin
      _T_714 <= 1'h0;
    end else begin
      if (_T_217) begin
        _T_714 <= _T_711;
      end
    end
    if (reset) begin
      _T_718 <= 13'h0;
    end else begin
      if (_T_220) begin
        _T_718 <= _T_715;
      end
    end
    if (reset) begin
      _T_722 <= 13'h0;
    end else begin
      if (_T_220) begin
        _T_722 <= _T_719;
      end
    end
    if (reset) begin
      _T_726 <= 13'h0;
    end else begin
      if (_T_223) begin
        _T_726 <= _T_719;
      end
    end
    if (reset) begin
      _T_730 <= 13'h0;
    end else begin
      if (_T_226) begin
        _T_730 <= _T_715;
      end
    end
    if (reset) begin
      _T_734 <= 13'h0;
    end else begin
      if (_T_226) begin
        _T_734 <= _T_719;
      end
    end
    if (reset) begin
      _T_738 <= 14'h0;
    end else begin
      if (_T_229) begin
        _T_738 <= _T_735;
      end
    end
    if (reset) begin
      _T_742 <= 12'h0;
    end else begin
      if (_T_232) begin
        _T_742 <= _T_739;
      end
    end
    if (reset) begin
      _T_746 <= 32'h0;
    end else begin
      if (_T_241) begin
        _T_746 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_750 <= 32'h0;
    end else begin
      if (_T_244) begin
        _T_750 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_754 <= 1'h0;
    end else begin
      if (_T_247) begin
        _T_754 <= _T_651;
      end
    end
    if (reset) begin
      _T_758 <= 16'h0;
    end else begin
      if (_T_250) begin
        _T_758 <= _T_755;
      end
    end
    if (reset) begin
      _T_762 <= 16'h0;
    end else begin
      if (_T_250) begin
        _T_762 <= _T_659;
      end
    end
    if (reset) begin
      _T_766 <= 16'h0;
    end else begin
      if (_T_253) begin
        _T_766 <= _T_755;
      end
    end
    if (reset) begin
      _T_770 <= 16'h0;
    end else begin
      if (_T_253) begin
        _T_770 <= _T_659;
      end
    end
    if (reset) begin
      _T_774 <= 1'h0;
    end else begin
      if (_T_256) begin
        _T_774 <= _T_651;
      end
    end
    if (reset) begin
      _T_778 <= 1'h0;
    end else begin
      if (_T_256) begin
        _T_778 <= _T_691;
      end
    end
    if (reset) begin
      _T_782 <= 2'h1;
    end else begin
      if (_T_256) begin
        _T_782 <= _T_779;
      end
    end
    if (reset) begin
      _T_786 <= 2'h1;
    end else begin
      if (_T_256) begin
        _T_786 <= _T_783;
      end
    end
    if (reset) begin
      _T_790 <= 1'h0;
    end else begin
      if (_T_256) begin
        _T_790 <= _T_787;
      end
    end
    if (reset) begin
      _T_794 <= 1'h0;
    end else begin
      if (_T_256) begin
        _T_794 <= _T_791;
      end
    end
    if (reset) begin
      _T_798 <= 1'h0;
    end else begin
      if (_T_256) begin
        _T_798 <= _T_711;
      end
    end
    if (reset) begin
      _T_802 <= 1'h0;
    end else begin
      if (_T_259) begin
        _T_802 <= _T_651;
      end
    end
    if (reset) begin
      _T_806 <= 1'h0;
    end else begin
      if (_T_277) begin
        _T_806 <= _T_651;
      end
    end
    if (reset) begin
      _T_810 <= 5'h0;
    end else begin
      if (_T_286) begin
        _T_810 <= _T_627;
      end
    end
    if (reset) begin
      _T_814 <= 3'h0;
    end else begin
      if (_T_286) begin
        _T_814 <= _T_647;
      end
    end
    if (reset) begin
      _T_818 <= 10'h0;
    end else begin
      if (_T_289) begin
        _T_818 <= _T_815;
      end
    end
    if (reset) begin
      _T_822 <= 10'h0;
    end else begin
      if (_T_289) begin
        _T_822 <= _T_819;
      end
    end
    if (reset) begin
      _T_826 <= 3'h0;
    end else begin
      if (_T_292) begin
        _T_826 <= _T_643;
      end
    end
    if (reset) begin
      _T_830 <= 5'h0;
    end else begin
      if (_T_292) begin
        _T_830 <= _T_631;
      end
    end
    if (reset) begin
      _T_834 <= 32'h0;
    end else begin
      if (_T_295) begin
        _T_834 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_838 <= 32'h0;
    end else begin
      if (_T_298) begin
        _T_838 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_842 <= 32'h0;
    end else begin
      if (_T_301) begin
        _T_842 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_846 <= 32'h0;
    end else begin
      if (_T_304) begin
        _T_846 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_850 <= 1'h0;
    end else begin
      if (_T_307) begin
        _T_850 <= _T_651;
      end
    end
    if (reset) begin
      _T_854 <= 1'h0;
    end else begin
      if (_T_310) begin
        _T_854 <= _T_651;
      end
    end
    if (reset) begin
      _T_858 <= 18'h0;
    end else begin
      if (_T_313) begin
        _T_858 <= _T_855;
      end
    end
    if (reset) begin
      _T_862 <= 13'h0;
    end else begin
      if (_T_316) begin
        _T_862 <= _T_719;
      end
    end
    if (reset) begin
      _T_866 <= 32'h0;
    end else begin
      if (_T_319) begin
        _T_866 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_870 <= 32'h0;
    end else begin
      if (_T_322) begin
        _T_870 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_874 <= 32'h0;
    end else begin
      if (_T_325) begin
        _T_874 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_878 <= 32'h0;
    end else begin
      if (_T_328) begin
        _T_878 <= io_reg_wr_data;
      end
    end
    if (reset) begin
      _T_882 <= 28'h0;
    end else begin
      if (_T_331) begin
        _T_882 <= _T_879;
      end
    end
    if (reset) begin
      _T_886 <= 6'h0;
    end else begin
      if (_T_334) begin
        _T_886 <= _T_883;
      end
    end
    if (reset) begin
      _T_890 <= 5'h0;
    end else begin
      if (_T_334) begin
        _T_890 <= _T_627;
      end
    end
    if (reset) begin
      _T_894 <= 6'h0;
    end else begin
      if (_T_334) begin
        _T_894 <= _T_703;
      end
    end
    if (reset) begin
      _T_898 <= 5'h0;
    end else begin
      if (_T_334) begin
        _T_898 <= _T_631;
      end
    end
    if (reset) begin
      _T_902 <= 16'h0;
    end else begin
      if (_T_337) begin
        _T_902 <= _T_659;
      end
    end
  end
endmodule
module NV_NVDLA_CSB_LOGIC( // @[:@1484.2]
  input         reset, // @[:@1486.4]
  input         io_clk, // @[:@1487.4]
  input         io_csb2dp_req_valid, // @[:@1487.4]
  input  [62:0] io_csb2dp_req_bits, // @[:@1487.4]
  output        io_csb2dp_resp_valid, // @[:@1487.4]
  output [33:0] io_csb2dp_resp_bits, // @[:@1487.4]
  input  [31:0] io_reg_rd_data, // @[:@1487.4]
  output [11:0] io_reg_offset, // @[:@1487.4]
  output [31:0] io_reg_wr_data, // @[:@1487.4]
  output        io_reg_wr_en // @[:@1487.4]
);
  reg  _T_43; // @[NV_NVDLA_CSB_LOGIC.scala 45:27:@1489.4]
  reg [31:0] _RAND_0;
  reg [62:0] _T_46; // @[NV_NVDLA_CSB_LOGIC.scala 46:25:@1490.4]
  reg [63:0] _RAND_1;
  wire [62:0] _GEN_0; // @[NV_NVDLA_CSB_LOGIC.scala 49:30:@1492.4]
  wire [21:0] _T_47; // @[NV_NVDLA_CSB_LOGIC.scala 54:26:@1495.4]
  wire  _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 56:27:@1497.4]
  wire  _T_50; // @[NV_NVDLA_CSB_LOGIC.scala 57:29:@1498.4]
  wire [23:0] _T_56; // @[Cat.scala 30:58:@1503.4]
  wire  _T_58; // @[NV_NVDLA_CSB_LOGIC.scala 68:32:@1508.4]
  wire  _T_59; // @[NV_NVDLA_CSB_LOGIC.scala 68:30:@1509.4]
  wire [33:0] _T_63; // @[Cat.scala 30:58:@1511.4]
  reg [33:0] _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 83:37:@1514.4]
  reg [63:0] _RAND_2;
  reg  _T_74; // @[NV_NVDLA_CSB_LOGIC.scala 84:40:@1515.4]
  reg [31:0] _RAND_3;
  wire  _T_75; // @[NV_NVDLA_CSB_LOGIC.scala 89:28:@1520.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSB_LOGIC.scala 89:42:@1521.6]
  wire [33:0] _GEN_2; // @[NV_NVDLA_CSB_LOGIC.scala 86:20:@1516.4]
  wire  _T_77; // @[NV_NVDLA_CSB_LOGIC.scala 92:59:@1525.4]
  assign _GEN_0 = io_csb2dp_req_valid ? io_csb2dp_req_bits : _T_46; // @[NV_NVDLA_CSB_LOGIC.scala 49:30:@1492.4]
  assign _T_47 = _T_46[21:0]; // @[NV_NVDLA_CSB_LOGIC.scala 54:26:@1495.4]
  assign _T_49 = _T_46[54]; // @[NV_NVDLA_CSB_LOGIC.scala 56:27:@1497.4]
  assign _T_50 = _T_46[55]; // @[NV_NVDLA_CSB_LOGIC.scala 57:29:@1498.4]
  assign _T_56 = {_T_47,2'h0}; // @[Cat.scala 30:58:@1503.4]
  assign _T_58 = ~ _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 68:32:@1508.4]
  assign _T_59 = _T_43 & _T_58; // @[NV_NVDLA_CSB_LOGIC.scala 68:30:@1509.4]
  assign _T_63 = {2'h0,io_reg_rd_data}; // @[Cat.scala 30:58:@1511.4]
  assign _T_75 = io_reg_wr_en & _T_50; // @[NV_NVDLA_CSB_LOGIC.scala 89:28:@1520.6]
  assign _GEN_1 = _T_75 ? 34'h200000000 : _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 89:42:@1521.6]
  assign _GEN_2 = _T_59 ? _T_63 : _GEN_1; // @[NV_NVDLA_CSB_LOGIC.scala 86:20:@1516.4]
  assign _T_77 = _T_75 | _T_59; // @[NV_NVDLA_CSB_LOGIC.scala 92:59:@1525.4]
  assign io_csb2dp_resp_valid = _T_74; // @[NV_NVDLA_CSB_LOGIC.scala 95:26:@1528.4]
  assign io_csb2dp_resp_bits = _T_71; // @[NV_NVDLA_CSB_LOGIC.scala 94:25:@1527.4]
  assign io_reg_offset = _T_56[11:0]; // @[NV_NVDLA_CSB_LOGIC.scala 65:19:@1504.4]
  assign io_reg_wr_data = _T_46[53:22]; // @[NV_NVDLA_CSB_LOGIC.scala 66:20:@1505.4]
  assign io_reg_wr_en = _T_43 & _T_49; // @[NV_NVDLA_CSB_LOGIC.scala 67:18:@1507.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_43 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_46 = _RAND_1[62:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_71 = _RAND_2[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_74 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      _T_43 <= io_csb2dp_req_valid;
    end
    if (reset) begin
      _T_46 <= 63'h0;
    end else begin
      if (io_csb2dp_req_valid) begin
        _T_46 <= io_csb2dp_req_bits;
      end
    end
    if (reset) begin
      _T_71 <= 34'h0;
    end else begin
      if (_T_59) begin
        _T_71 <= _T_63;
      end else begin
        if (_T_75) begin
          _T_71 <= 34'h200000000;
        end
      end
    end
    if (reset) begin
      _T_74 <= 1'h0;
    end else begin
      _T_74 <= _T_77;
    end
  end
endmodule
module NV_NVDLA_CDMA_regfile( // @[:@1530.2]
  input         reset, // @[:@1532.4]
  input         io_nvdla_core_clk, // @[:@1533.4]
  input         io_csb2cdma_req_valid, // @[:@1533.4]
  input  [62:0] io_csb2cdma_req_bits, // @[:@1533.4]
  output        io_csb2cdma_resp_valid, // @[:@1533.4]
  output [33:0] io_csb2cdma_resp_bits, // @[:@1533.4]
  input         io_dp2reg_done, // @[:@1533.4]
  input  [31:0] io_dp2reg_dc_rd_latency, // @[:@1533.4]
  input  [31:0] io_dp2reg_dc_rd_stall, // @[:@1533.4]
  input  [31:0] io_dp2reg_img_rd_latency, // @[:@1533.4]
  input  [31:0] io_dp2reg_img_rd_stall, // @[:@1533.4]
  input         io_dp2reg_dat_flush_done, // @[:@1533.4]
  input         io_dp2reg_wt_flush_done, // @[:@1533.4]
  input  [31:0] io_dp2reg_wt_rd_stall, // @[:@1533.4]
  output        io_dp2reg_consumer, // @[:@1533.4]
  output [4:0]  io_reg2dp_field_data_bank, // @[:@1533.4]
  output [4:0]  io_reg2dp_field_weight_bank, // @[:@1533.4]
  output [4:0]  io_reg2dp_field_batches, // @[:@1533.4]
  output [31:0] io_reg2dp_field_batch_stride, // @[:@1533.4]
  output        io_reg2dp_field_cvt_en, // @[:@1533.4]
  output [5:0]  io_reg2dp_field_cvt_truncate, // @[:@1533.4]
  output [15:0] io_reg2dp_field_cvt_offset, // @[:@1533.4]
  output [15:0] io_reg2dp_field_cvt_scale, // @[:@1533.4]
  output [31:0] io_reg2dp_field_datain_addr_high_0, // @[:@1533.4]
  output [31:0] io_reg2dp_field_datain_addr_high_1, // @[:@1533.4]
  output [31:0] io_reg2dp_field_datain_addr_low_0, // @[:@1533.4]
  output [31:0] io_reg2dp_field_datain_addr_low_1, // @[:@1533.4]
  output        io_reg2dp_field_line_packed, // @[:@1533.4]
  output        io_reg2dp_field_surf_packed, // @[:@1533.4]
  output        io_reg2dp_field_datain_ram_type, // @[:@1533.4]
  output        io_reg2dp_field_datain_format, // @[:@1533.4]
  output [5:0]  io_reg2dp_field_pixel_format, // @[:@1533.4]
  output        io_reg2dp_field_pixel_sign_override, // @[:@1533.4]
  output [12:0] io_reg2dp_field_datain_height, // @[:@1533.4]
  output [12:0] io_reg2dp_field_datain_width, // @[:@1533.4]
  output [12:0] io_reg2dp_field_datain_channel, // @[:@1533.4]
  output [13:0] io_reg2dp_field_entries, // @[:@1533.4]
  output [11:0] io_reg2dp_field_grains, // @[:@1533.4]
  output [31:0] io_reg2dp_field_line_stride, // @[:@1533.4]
  output [31:0] io_reg2dp_field_uv_line_stride, // @[:@1533.4]
  output        io_reg2dp_field_mean_format, // @[:@1533.4]
  output [15:0] io_reg2dp_field_mean_gu, // @[:@1533.4]
  output [15:0] io_reg2dp_field_mean_ry, // @[:@1533.4]
  output [15:0] io_reg2dp_field_mean_ax, // @[:@1533.4]
  output [15:0] io_reg2dp_field_mean_bv, // @[:@1533.4]
  output        io_reg2dp_field_conv_mode, // @[:@1533.4]
  output        io_reg2dp_field_data_reuse, // @[:@1533.4]
  output [1:0]  io_reg2dp_field_proc_precision, // @[:@1533.4]
  output        io_reg2dp_field_skip_data_rls, // @[:@1533.4]
  output        io_reg2dp_field_skip_weight_rls, // @[:@1533.4]
  output        io_reg2dp_field_weight_reuse, // @[:@1533.4]
  output        io_reg2dp_field_dma_en, // @[:@1533.4]
  output [4:0]  io_reg2dp_field_pixel_x_offset, // @[:@1533.4]
  output [31:0] io_reg2dp_field_surf_stride, // @[:@1533.4]
  output [31:0] io_reg2dp_field_weight_addr_high, // @[:@1533.4]
  output [31:0] io_reg2dp_field_weight_addr_low, // @[:@1533.4]
  output [31:0] io_reg2dp_field_weight_bytes, // @[:@1533.4]
  output        io_reg2dp_field_weight_ram_type, // @[:@1533.4]
  output [17:0] io_reg2dp_field_byte_per_kernel, // @[:@1533.4]
  output [12:0] io_reg2dp_field_weight_kernel, // @[:@1533.4]
  output [4:0]  io_reg2dp_field_pad_left, // @[:@1533.4]
  output [5:0]  io_reg2dp_field_pad_right, // @[:@1533.4]
  output [15:0] io_reg2dp_field_pad_value, // @[:@1533.4]
  output        io_reg2dp_op_en // @[:@1533.4]
);
  wire  NV_NVDLA_CDMA_single_reg_clock; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_single_reg_reset; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [31:0] NV_NVDLA_CDMA_single_reg_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [11:0] NV_NVDLA_CDMA_single_reg_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [31:0] NV_NVDLA_CDMA_single_reg_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_single_reg_io_reg_wr_en; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_single_reg_io_producer; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [3:0] NV_NVDLA_CDMA_single_reg_io_arb_wmb; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_single_reg_io_flush_done; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_single_reg_io_consumer; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [1:0] NV_NVDLA_CDMA_single_reg_io_status_0; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire [1:0] NV_NVDLA_CDMA_single_reg_io_status_1; // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
  wire  NV_NVDLA_CDMA_dual_reg_reset; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [11:0] NV_NVDLA_CDMA_dual_reg_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_reg_wr_en; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_data_bank; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_weight_bank; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_batches; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_batch_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_io_field_conv_x_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_io_field_conv_y_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_cvt_en; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_io_field_cvt_truncate; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_cvt_offset; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_cvt_scale; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_cya; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_0; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_1; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_0; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_1; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_line_packed; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_surf_packed; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_datain_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_datain_format; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_io_field_pixel_format; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_pixel_mapping; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_pixel_sign_override; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_height; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_width; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_channel; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_height_ext; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_datain_width_ext; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [13:0] NV_NVDLA_CDMA_dual_reg_io_field_entries; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [11:0] NV_NVDLA_CDMA_dual_reg_io_field_grains; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_uv_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_mean_format; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_mean_gu; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_mean_ry; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_mean_ax; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_mean_bv; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_conv_mode; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_data_reuse; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [1:0] NV_NVDLA_CDMA_dual_reg_io_field_in_precision; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [1:0] NV_NVDLA_CDMA_dual_reg_io_field_proc_precision; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_skip_data_rls; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_skip_weight_rls; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_weight_reuse; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_nan_to_zero; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_dma_en; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_pixel_x_offset; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_io_field_pixel_y_offset; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [9:0] NV_NVDLA_CDMA_dual_reg_io_field_rsv_per_line; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [9:0] NV_NVDLA_CDMA_dual_reg_io_field_rsv_per_uv_line; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_io_field_rsv_height; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_rsv_y_index; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_surf_stride; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_weight_bytes; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_weight_format; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_field_weight_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [17:0] NV_NVDLA_CDMA_dual_reg_io_field_byte_per_kernel; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_io_field_weight_kernel; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_wgs_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_wgs_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_wmb_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_field_wmb_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [27:0] NV_NVDLA_CDMA_dual_reg_io_field_wmb_bytes; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_io_field_pad_bottom; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_pad_left; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_io_field_pad_right; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_io_field_pad_top; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_io_field_pad_value; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_op_en_trigger; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_inf_data_num; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_inf_weight_num; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_nan_data_num; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_nan_weight_num; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_io_op_en; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_dat_rd_latency; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_dat_rd_stall; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_wt_rd_latency; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_io_wt_rd_stall; // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_reset; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [11:0] NV_NVDLA_CDMA_dual_reg_1_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_en; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_data_bank; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bank; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_batches; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_batch_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_1_io_field_conv_x_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_1_io_field_conv_y_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_en; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_truncate; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_offset; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_scale; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_cya; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_0; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_1; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_0; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_1; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_line_packed; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_surf_packed; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_datain_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_datain_format; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_format; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_mapping; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_sign_override; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_height; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_width; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_channel; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_height_ext; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_datain_width_ext; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [13:0] NV_NVDLA_CDMA_dual_reg_1_io_field_entries; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [11:0] NV_NVDLA_CDMA_dual_reg_1_io_field_grains; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_uv_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_mean_format; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_mean_gu; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ry; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ax; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_mean_bv; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_conv_mode; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_data_reuse; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [1:0] NV_NVDLA_CDMA_dual_reg_1_io_field_in_precision; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [1:0] NV_NVDLA_CDMA_dual_reg_1_io_field_proc_precision; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_skip_data_rls; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_skip_weight_rls; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_weight_reuse; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_nan_to_zero; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_dma_en; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_x_offset; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_y_offset; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [9:0] NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_per_line; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [9:0] NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_per_uv_line; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [2:0] NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_height; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_y_index; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_surf_stride; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bytes; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_weight_format; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_field_weight_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [17:0] NV_NVDLA_CDMA_dual_reg_1_io_field_byte_per_kernel; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [12:0] NV_NVDLA_CDMA_dual_reg_1_io_field_weight_kernel; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_wgs_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_wgs_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [27:0] NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_bytes; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pad_bottom; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pad_left; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [5:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pad_right; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [4:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pad_top; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [15:0] NV_NVDLA_CDMA_dual_reg_1_io_field_pad_value; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_op_en_trigger; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_inf_data_num; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_inf_weight_num; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_nan_data_num; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_nan_weight_num; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CDMA_dual_reg_1_io_op_en; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_latency; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_stall; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_latency; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire [31:0] NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_stall; // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
  wire  NV_NVDLA_CSB_LOGIC_reset; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire  NV_NVDLA_CSB_LOGIC_io_clk; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire  NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire [62:0] NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire  NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire [33:0] NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire [31:0] NV_NVDLA_CSB_LOGIC_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire [11:0] NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire [31:0] NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  wire  NV_NVDLA_CSB_LOGIC_io_reg_wr_en; // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
  reg  _T_203; // @[NV_NVDLA_CDMA_regfile.scala 69:38:@1535.4]
  reg [31:0] _RAND_0;
  reg  _T_206; // @[NV_NVDLA_CDMA_regfile.scala 70:36:@1536.4]
  reg [31:0] _RAND_1;
  reg  _T_221; // @[NV_NVDLA_CDMA_regfile.scala 94:34:@1556.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_224; // @[NV_NVDLA_CDMA_regfile.scala 95:41:@1557.4]
  reg [31:0] _RAND_3;
  reg [31:0] _T_227; // @[NV_NVDLA_CDMA_regfile.scala 96:43:@1558.4]
  reg [31:0] _RAND_4;
  reg [31:0] _T_230; // @[NV_NVDLA_CDMA_regfile.scala 97:41:@1559.4]
  reg [31:0] _RAND_5;
  reg [31:0] _T_233; // @[NV_NVDLA_CDMA_regfile.scala 98:43:@1560.4]
  reg [31:0] _RAND_6;
  reg [31:0] _T_236; // @[NV_NVDLA_CDMA_regfile.scala 99:43:@1561.4]
  reg [31:0] _RAND_7;
  reg [31:0] _T_239; // @[NV_NVDLA_CDMA_regfile.scala 100:41:@1562.4]
  reg [31:0] _RAND_8;
  reg [31:0] _T_242; // @[NV_NVDLA_CDMA_regfile.scala 101:42:@1563.4]
  reg [31:0] _RAND_9;
  reg [31:0] _T_245; // @[NV_NVDLA_CDMA_regfile.scala 102:40:@1564.4]
  reg [31:0] _RAND_10;
  reg  _T_250; // @[NV_NVDLA_CDMA_regfile.scala 123:34:@1582.4]
  reg [31:0] _RAND_11;
  reg [31:0] _T_253; // @[NV_NVDLA_CDMA_regfile.scala 124:41:@1583.4]
  reg [31:0] _RAND_12;
  reg [31:0] _T_256; // @[NV_NVDLA_CDMA_regfile.scala 125:43:@1584.4]
  reg [31:0] _RAND_13;
  reg [31:0] _T_259; // @[NV_NVDLA_CDMA_regfile.scala 126:41:@1585.4]
  reg [31:0] _RAND_14;
  reg [31:0] _T_262; // @[NV_NVDLA_CDMA_regfile.scala 127:43:@1586.4]
  reg [31:0] _RAND_15;
  reg [31:0] _T_265; // @[NV_NVDLA_CDMA_regfile.scala 128:43:@1587.4]
  reg [31:0] _RAND_16;
  reg [31:0] _T_268; // @[NV_NVDLA_CDMA_regfile.scala 129:41:@1588.4]
  reg [31:0] _RAND_17;
  reg [31:0] _T_271; // @[NV_NVDLA_CDMA_regfile.scala 130:42:@1589.4]
  reg [31:0] _RAND_18;
  reg [31:0] _T_274; // @[NV_NVDLA_CDMA_regfile.scala 131:40:@1590.4]
  reg [31:0] _RAND_19;
  wire  _T_275; // @[NV_NVDLA_CDMA_regfile.scala 156:33:@1607.4]
  wire  _GEN_0; // @[NV_NVDLA_CDMA_regfile.scala 158:25:@1608.4]
  wire  _T_277; // @[NV_NVDLA_CDMA_regfile.scala 169:44:@1612.4]
  wire [1:0] _T_283; // @[NV_NVDLA_CDMA_regfile.scala 170:27:@1614.4]
  wire [1:0] _T_284; // @[NV_NVDLA_CDMA_regfile.scala 169:27:@1615.4]
  wire  _T_286; // @[NV_NVDLA_CDMA_regfile.scala 173:44:@1617.4]
  wire  _T_289; // @[NV_NVDLA_CDMA_regfile.scala 174:48:@1618.4]
  wire [1:0] _T_292; // @[NV_NVDLA_CDMA_regfile.scala 174:27:@1619.4]
  wire [1:0] _T_293; // @[NV_NVDLA_CDMA_regfile.scala 173:27:@1620.4]
  reg [2:0] _T_296; // @[NV_NVDLA_CDMA_regfile.scala 182:35:@1622.4]
  reg [31:0] _RAND_20;
  wire  _T_297; // @[NV_NVDLA_CDMA_regfile.scala 183:33:@1623.4]
  wire  _T_298; // @[NV_NVDLA_CDMA_regfile.scala 183:50:@1624.4]
  wire [31:0] _T_210; // @[NV_NVDLA_CDMA_regfile.scala 72:27:@1538.4 NV_NVDLA_CDMA_regfile.scala 229:17:@1705.4]
  wire  _T_299; // @[NV_NVDLA_CDMA_regfile.scala 183:88:@1625.4]
  wire  _T_302; // @[NV_NVDLA_CDMA_regfile.scala 184:48:@1627.4]
  wire  _T_304; // @[NV_NVDLA_CDMA_regfile.scala 184:32:@1628.4]
  wire  _T_305; // @[NV_NVDLA_CDMA_regfile.scala 183:32:@1629.4]
  wire  _T_306; // @[NV_NVDLA_CDMA_regfile.scala 188:34:@1631.4]
  wire  _T_307; // @[NV_NVDLA_CDMA_regfile.scala 188:51:@1632.4]
  wire  _T_311; // @[NV_NVDLA_CDMA_regfile.scala 189:49:@1635.4]
  wire  _T_313; // @[NV_NVDLA_CDMA_regfile.scala 189:33:@1636.4]
  wire  _T_314; // @[NV_NVDLA_CDMA_regfile.scala 188:33:@1637.4]
  wire  _T_315; // @[NV_NVDLA_CDMA_regfile.scala 193:31:@1639.4]
  wire [1:0] _T_317; // @[NV_NVDLA_CDMA_regfile.scala 194:89:@1640.4]
  wire [2:0] _T_318; // @[Cat.scala 30:58:@1641.4]
  wire [2:0] _T_319; // @[NV_NVDLA_CDMA_regfile.scala 194:33:@1642.4]
  wire [11:0] _T_208; // @[NV_NVDLA_CDMA_regfile.scala 71:26:@1537.4 NV_NVDLA_CDMA_regfile.scala 227:16:@1703.4]
  wire [31:0] _GEN_20; // @[NV_NVDLA_CDMA_regfile.scala 207:41:@1663.4]
  wire  _T_336; // @[NV_NVDLA_CDMA_regfile.scala 207:41:@1663.4]
  wire  _T_342; // @[NV_NVDLA_CDMA_regfile.scala 208:39:@1666.4]
  wire  _T_344; // @[NV_NVDLA_CDMA_regfile.scala 208:83:@1667.4]
  wire  _T_345; // @[NV_NVDLA_CDMA_regfile.scala 208:64:@1668.4]
  wire  _T_350; // @[NV_NVDLA_CDMA_regfile.scala 209:83:@1671.4]
  wire  _T_351; // @[NV_NVDLA_CDMA_regfile.scala 209:64:@1672.4]
  wire  _T_333; // @[NV_NVDLA_CDMA_regfile.scala 206:25:@1661.4 NV_NVDLA_CDMA_regfile.scala 228:15:@1704.4]
  wire  _T_353; // @[NV_NVDLA_CDMA_regfile.scala 212:31:@1675.4]
  wire  _T_357; // @[NV_NVDLA_CDMA_regfile.scala 213:31:@1679.4]
  wire [31:0] _T_364; // @[Bitwise.scala 72:12:@1684.4]
  wire [31:0] _T_365; // @[NV_NVDLA_CDMA_regfile.scala 215:43:@1685.4]
  wire [31:0] _T_369; // @[Bitwise.scala 72:12:@1687.4]
  wire [31:0] _T_370; // @[NV_NVDLA_CDMA_regfile.scala 216:44:@1688.4]
  wire [31:0] _T_371; // @[NV_NVDLA_CDMA_regfile.scala 215:59:@1689.4]
  wire [31:0] _T_375; // @[Bitwise.scala 72:12:@1691.4]
  wire [31:0] _T_376; // @[NV_NVDLA_CDMA_regfile.scala 217:43:@1692.4]
  wire  _T_448; // @[NV_NVDLA_CDMA_regfile.scala 251:50:@1777.4]
  wire  _T_449; // @[NV_NVDLA_CDMA_regfile.scala 256:43:@1779.4]
  wire  _T_450; // @[NV_NVDLA_CDMA_regfile.scala 256:41:@1780.4]
  wire  _T_452; // @[NV_NVDLA_CDMA_regfile.scala 257:42:@1782.4]
  wire  _T_453; // @[NV_NVDLA_CDMA_regfile.scala 258:41:@1783.4]
  wire  _T_454; // @[NV_NVDLA_CDMA_regfile.scala 260:43:@1784.4]
  wire  _T_455; // @[NV_NVDLA_CDMA_regfile.scala 260:41:@1785.4]
  wire  _T_457; // @[NV_NVDLA_CDMA_regfile.scala 261:42:@1787.4]
  wire  _T_458; // @[NV_NVDLA_CDMA_regfile.scala 262:41:@1788.4]
  wire [31:0] _T_460; // @[NV_NVDLA_CDMA_regfile.scala 269:41:@1789.4]
  wire [31:0] _T_461; // @[NV_NVDLA_CDMA_regfile.scala 268:41:@1790.4]
  wire [31:0] _T_463; // @[NV_NVDLA_CDMA_regfile.scala 272:41:@1791.4]
  wire [31:0] _T_464; // @[NV_NVDLA_CDMA_regfile.scala 271:41:@1792.4]
  wire [31:0] _T_466; // @[NV_NVDLA_CDMA_regfile.scala 275:41:@1793.4]
  wire [31:0] _T_467; // @[NV_NVDLA_CDMA_regfile.scala 274:39:@1794.4]
  wire [31:0] _T_469; // @[NV_NVDLA_CDMA_regfile.scala 278:41:@1795.4]
  wire [31:0] _T_470; // @[NV_NVDLA_CDMA_regfile.scala 277:39:@1796.4]
  wire [31:0] _GEN_4; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  wire [31:0] _GEN_5; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  wire [31:0] _GEN_6; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  wire [31:0] _GEN_7; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  wire [31:0] _T_472; // @[NV_NVDLA_CDMA_regfile.scala 290:41:@1803.4]
  wire [31:0] _T_473; // @[NV_NVDLA_CDMA_regfile.scala 289:41:@1804.4]
  wire [31:0] _T_475; // @[NV_NVDLA_CDMA_regfile.scala 293:41:@1805.4]
  wire [31:0] _T_476; // @[NV_NVDLA_CDMA_regfile.scala 292:41:@1806.4]
  wire [31:0] _T_478; // @[NV_NVDLA_CDMA_regfile.scala 296:41:@1807.4]
  wire [31:0] _T_479; // @[NV_NVDLA_CDMA_regfile.scala 295:39:@1808.4]
  wire [31:0] _T_481; // @[NV_NVDLA_CDMA_regfile.scala 299:41:@1809.4]
  wire [31:0] _T_482; // @[NV_NVDLA_CDMA_regfile.scala 298:39:@1810.4]
  wire [31:0] _GEN_8; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  wire [31:0] _GEN_9; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  wire [31:0] _GEN_10; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  wire [31:0] _GEN_11; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  wire [31:0] _T_484; // @[NV_NVDLA_CDMA_regfile.scala 314:41:@1817.4]
  wire [31:0] _T_485; // @[NV_NVDLA_CDMA_regfile.scala 313:38:@1818.4]
  wire [31:0] _T_487; // @[NV_NVDLA_CDMA_regfile.scala 317:41:@1819.4]
  wire [31:0] _T_488; // @[NV_NVDLA_CDMA_regfile.scala 316:40:@1820.4]
  wire [31:0] _T_490; // @[NV_NVDLA_CDMA_regfile.scala 319:102:@1822.4]
  wire [31:0] _T_492; // @[NV_NVDLA_CDMA_regfile.scala 320:41:@1823.4]
  wire [31:0] _T_493; // @[NV_NVDLA_CDMA_regfile.scala 319:39:@1824.4]
  wire [31:0] _T_495; // @[NV_NVDLA_CDMA_regfile.scala 322:108:@1826.4]
  wire [31:0] _T_497; // @[NV_NVDLA_CDMA_regfile.scala 323:41:@1827.4]
  wire [31:0] _T_498; // @[NV_NVDLA_CDMA_regfile.scala 322:41:@1828.4]
  wire [31:0] _GEN_12; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  wire [31:0] _GEN_13; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  wire [31:0] _GEN_14; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  wire [31:0] _GEN_15; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  wire [31:0] _T_500; // @[NV_NVDLA_CDMA_regfile.scala 334:41:@1835.4]
  wire [31:0] _T_501; // @[NV_NVDLA_CDMA_regfile.scala 333:38:@1836.4]
  wire [31:0] _T_503; // @[NV_NVDLA_CDMA_regfile.scala 337:41:@1837.4]
  wire [31:0] _T_504; // @[NV_NVDLA_CDMA_regfile.scala 336:40:@1838.4]
  wire [31:0] _T_508; // @[NV_NVDLA_CDMA_regfile.scala 340:41:@1841.4]
  wire [31:0] _T_509; // @[NV_NVDLA_CDMA_regfile.scala 339:39:@1842.4]
  wire [31:0] _T_513; // @[NV_NVDLA_CDMA_regfile.scala 343:41:@1845.4]
  wire [31:0] _T_514; // @[NV_NVDLA_CDMA_regfile.scala 342:41:@1846.4]
  wire [31:0] _GEN_16; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  wire [31:0] _GEN_17; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  wire [31:0] _GEN_18; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  wire [31:0] _GEN_19; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  wire  _T_214; // @[NV_NVDLA_CDMA_regfile.scala 74:31:@1540.4 NV_NVDLA_CDMA_regfile.scala 169:21:@1616.4]
  wire  _T_216; // @[NV_NVDLA_CDMA_regfile.scala 75:31:@1541.4 NV_NVDLA_CDMA_regfile.scala 173:21:@1621.4]
  NV_NVDLA_CDMA_single_reg NV_NVDLA_CDMA_single_reg ( // @[NV_NVDLA_CDMA_regfile.scala 77:30:@1542.4]
    .clock(NV_NVDLA_CDMA_single_reg_clock),
    .reset(NV_NVDLA_CDMA_single_reg_reset),
    .io_reg_rd_data(NV_NVDLA_CDMA_single_reg_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CDMA_single_reg_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CDMA_single_reg_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CDMA_single_reg_io_reg_wr_en),
    .io_producer(NV_NVDLA_CDMA_single_reg_io_producer),
    .io_arb_wmb(NV_NVDLA_CDMA_single_reg_io_arb_wmb),
    .io_flush_done(NV_NVDLA_CDMA_single_reg_io_flush_done),
    .io_consumer(NV_NVDLA_CDMA_single_reg_io_consumer),
    .io_status_0(NV_NVDLA_CDMA_single_reg_io_status_0),
    .io_status_1(NV_NVDLA_CDMA_single_reg_io_status_1)
  );
  NV_NVDLA_CDMA_dual_reg NV_NVDLA_CDMA_dual_reg ( // @[NV_NVDLA_CDMA_regfile.scala 104:31:@1565.4]
    .reset(NV_NVDLA_CDMA_dual_reg_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_dual_reg_io_nvdla_core_clk),
    .io_reg_rd_data(NV_NVDLA_CDMA_dual_reg_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CDMA_dual_reg_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CDMA_dual_reg_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CDMA_dual_reg_io_reg_wr_en),
    .io_field_data_bank(NV_NVDLA_CDMA_dual_reg_io_field_data_bank),
    .io_field_weight_bank(NV_NVDLA_CDMA_dual_reg_io_field_weight_bank),
    .io_field_batches(NV_NVDLA_CDMA_dual_reg_io_field_batches),
    .io_field_batch_stride(NV_NVDLA_CDMA_dual_reg_io_field_batch_stride),
    .io_field_conv_x_stride(NV_NVDLA_CDMA_dual_reg_io_field_conv_x_stride),
    .io_field_conv_y_stride(NV_NVDLA_CDMA_dual_reg_io_field_conv_y_stride),
    .io_field_cvt_en(NV_NVDLA_CDMA_dual_reg_io_field_cvt_en),
    .io_field_cvt_truncate(NV_NVDLA_CDMA_dual_reg_io_field_cvt_truncate),
    .io_field_cvt_offset(NV_NVDLA_CDMA_dual_reg_io_field_cvt_offset),
    .io_field_cvt_scale(NV_NVDLA_CDMA_dual_reg_io_field_cvt_scale),
    .io_field_cya(NV_NVDLA_CDMA_dual_reg_io_field_cya),
    .io_field_datain_addr_high_0(NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_0),
    .io_field_datain_addr_high_1(NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_1),
    .io_field_datain_addr_low_0(NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_0),
    .io_field_datain_addr_low_1(NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_1),
    .io_field_line_packed(NV_NVDLA_CDMA_dual_reg_io_field_line_packed),
    .io_field_surf_packed(NV_NVDLA_CDMA_dual_reg_io_field_surf_packed),
    .io_field_datain_ram_type(NV_NVDLA_CDMA_dual_reg_io_field_datain_ram_type),
    .io_field_datain_format(NV_NVDLA_CDMA_dual_reg_io_field_datain_format),
    .io_field_pixel_format(NV_NVDLA_CDMA_dual_reg_io_field_pixel_format),
    .io_field_pixel_mapping(NV_NVDLA_CDMA_dual_reg_io_field_pixel_mapping),
    .io_field_pixel_sign_override(NV_NVDLA_CDMA_dual_reg_io_field_pixel_sign_override),
    .io_field_datain_height(NV_NVDLA_CDMA_dual_reg_io_field_datain_height),
    .io_field_datain_width(NV_NVDLA_CDMA_dual_reg_io_field_datain_width),
    .io_field_datain_channel(NV_NVDLA_CDMA_dual_reg_io_field_datain_channel),
    .io_field_datain_height_ext(NV_NVDLA_CDMA_dual_reg_io_field_datain_height_ext),
    .io_field_datain_width_ext(NV_NVDLA_CDMA_dual_reg_io_field_datain_width_ext),
    .io_field_entries(NV_NVDLA_CDMA_dual_reg_io_field_entries),
    .io_field_grains(NV_NVDLA_CDMA_dual_reg_io_field_grains),
    .io_field_line_stride(NV_NVDLA_CDMA_dual_reg_io_field_line_stride),
    .io_field_uv_line_stride(NV_NVDLA_CDMA_dual_reg_io_field_uv_line_stride),
    .io_field_mean_format(NV_NVDLA_CDMA_dual_reg_io_field_mean_format),
    .io_field_mean_gu(NV_NVDLA_CDMA_dual_reg_io_field_mean_gu),
    .io_field_mean_ry(NV_NVDLA_CDMA_dual_reg_io_field_mean_ry),
    .io_field_mean_ax(NV_NVDLA_CDMA_dual_reg_io_field_mean_ax),
    .io_field_mean_bv(NV_NVDLA_CDMA_dual_reg_io_field_mean_bv),
    .io_field_conv_mode(NV_NVDLA_CDMA_dual_reg_io_field_conv_mode),
    .io_field_data_reuse(NV_NVDLA_CDMA_dual_reg_io_field_data_reuse),
    .io_field_in_precision(NV_NVDLA_CDMA_dual_reg_io_field_in_precision),
    .io_field_proc_precision(NV_NVDLA_CDMA_dual_reg_io_field_proc_precision),
    .io_field_skip_data_rls(NV_NVDLA_CDMA_dual_reg_io_field_skip_data_rls),
    .io_field_skip_weight_rls(NV_NVDLA_CDMA_dual_reg_io_field_skip_weight_rls),
    .io_field_weight_reuse(NV_NVDLA_CDMA_dual_reg_io_field_weight_reuse),
    .io_field_nan_to_zero(NV_NVDLA_CDMA_dual_reg_io_field_nan_to_zero),
    .io_field_dma_en(NV_NVDLA_CDMA_dual_reg_io_field_dma_en),
    .io_field_pixel_x_offset(NV_NVDLA_CDMA_dual_reg_io_field_pixel_x_offset),
    .io_field_pixel_y_offset(NV_NVDLA_CDMA_dual_reg_io_field_pixel_y_offset),
    .io_field_rsv_per_line(NV_NVDLA_CDMA_dual_reg_io_field_rsv_per_line),
    .io_field_rsv_per_uv_line(NV_NVDLA_CDMA_dual_reg_io_field_rsv_per_uv_line),
    .io_field_rsv_height(NV_NVDLA_CDMA_dual_reg_io_field_rsv_height),
    .io_field_rsv_y_index(NV_NVDLA_CDMA_dual_reg_io_field_rsv_y_index),
    .io_field_surf_stride(NV_NVDLA_CDMA_dual_reg_io_field_surf_stride),
    .io_field_weight_addr_high(NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_high),
    .io_field_weight_addr_low(NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_low),
    .io_field_weight_bytes(NV_NVDLA_CDMA_dual_reg_io_field_weight_bytes),
    .io_field_weight_format(NV_NVDLA_CDMA_dual_reg_io_field_weight_format),
    .io_field_weight_ram_type(NV_NVDLA_CDMA_dual_reg_io_field_weight_ram_type),
    .io_field_byte_per_kernel(NV_NVDLA_CDMA_dual_reg_io_field_byte_per_kernel),
    .io_field_weight_kernel(NV_NVDLA_CDMA_dual_reg_io_field_weight_kernel),
    .io_field_wgs_addr_high(NV_NVDLA_CDMA_dual_reg_io_field_wgs_addr_high),
    .io_field_wgs_addr_low(NV_NVDLA_CDMA_dual_reg_io_field_wgs_addr_low),
    .io_field_wmb_addr_high(NV_NVDLA_CDMA_dual_reg_io_field_wmb_addr_high),
    .io_field_wmb_addr_low(NV_NVDLA_CDMA_dual_reg_io_field_wmb_addr_low),
    .io_field_wmb_bytes(NV_NVDLA_CDMA_dual_reg_io_field_wmb_bytes),
    .io_field_pad_bottom(NV_NVDLA_CDMA_dual_reg_io_field_pad_bottom),
    .io_field_pad_left(NV_NVDLA_CDMA_dual_reg_io_field_pad_left),
    .io_field_pad_right(NV_NVDLA_CDMA_dual_reg_io_field_pad_right),
    .io_field_pad_top(NV_NVDLA_CDMA_dual_reg_io_field_pad_top),
    .io_field_pad_value(NV_NVDLA_CDMA_dual_reg_io_field_pad_value),
    .io_op_en_trigger(NV_NVDLA_CDMA_dual_reg_io_op_en_trigger),
    .io_inf_data_num(NV_NVDLA_CDMA_dual_reg_io_inf_data_num),
    .io_inf_weight_num(NV_NVDLA_CDMA_dual_reg_io_inf_weight_num),
    .io_nan_data_num(NV_NVDLA_CDMA_dual_reg_io_nan_data_num),
    .io_nan_weight_num(NV_NVDLA_CDMA_dual_reg_io_nan_weight_num),
    .io_op_en(NV_NVDLA_CDMA_dual_reg_io_op_en),
    .io_dat_rd_latency(NV_NVDLA_CDMA_dual_reg_io_dat_rd_latency),
    .io_dat_rd_stall(NV_NVDLA_CDMA_dual_reg_io_dat_rd_stall),
    .io_wt_rd_latency(NV_NVDLA_CDMA_dual_reg_io_wt_rd_latency),
    .io_wt_rd_stall(NV_NVDLA_CDMA_dual_reg_io_wt_rd_stall)
  );
  NV_NVDLA_CDMA_dual_reg NV_NVDLA_CDMA_dual_reg_1 ( // @[NV_NVDLA_CDMA_regfile.scala 133:31:@1591.4]
    .reset(NV_NVDLA_CDMA_dual_reg_1_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_dual_reg_1_io_nvdla_core_clk),
    .io_reg_rd_data(NV_NVDLA_CDMA_dual_reg_1_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CDMA_dual_reg_1_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_en),
    .io_field_data_bank(NV_NVDLA_CDMA_dual_reg_1_io_field_data_bank),
    .io_field_weight_bank(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bank),
    .io_field_batches(NV_NVDLA_CDMA_dual_reg_1_io_field_batches),
    .io_field_batch_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_batch_stride),
    .io_field_conv_x_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_conv_x_stride),
    .io_field_conv_y_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_conv_y_stride),
    .io_field_cvt_en(NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_en),
    .io_field_cvt_truncate(NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_truncate),
    .io_field_cvt_offset(NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_offset),
    .io_field_cvt_scale(NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_scale),
    .io_field_cya(NV_NVDLA_CDMA_dual_reg_1_io_field_cya),
    .io_field_datain_addr_high_0(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_0),
    .io_field_datain_addr_high_1(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_1),
    .io_field_datain_addr_low_0(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_0),
    .io_field_datain_addr_low_1(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_1),
    .io_field_line_packed(NV_NVDLA_CDMA_dual_reg_1_io_field_line_packed),
    .io_field_surf_packed(NV_NVDLA_CDMA_dual_reg_1_io_field_surf_packed),
    .io_field_datain_ram_type(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_ram_type),
    .io_field_datain_format(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_format),
    .io_field_pixel_format(NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_format),
    .io_field_pixel_mapping(NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_mapping),
    .io_field_pixel_sign_override(NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_sign_override),
    .io_field_datain_height(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_height),
    .io_field_datain_width(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_width),
    .io_field_datain_channel(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_channel),
    .io_field_datain_height_ext(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_height_ext),
    .io_field_datain_width_ext(NV_NVDLA_CDMA_dual_reg_1_io_field_datain_width_ext),
    .io_field_entries(NV_NVDLA_CDMA_dual_reg_1_io_field_entries),
    .io_field_grains(NV_NVDLA_CDMA_dual_reg_1_io_field_grains),
    .io_field_line_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_line_stride),
    .io_field_uv_line_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_uv_line_stride),
    .io_field_mean_format(NV_NVDLA_CDMA_dual_reg_1_io_field_mean_format),
    .io_field_mean_gu(NV_NVDLA_CDMA_dual_reg_1_io_field_mean_gu),
    .io_field_mean_ry(NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ry),
    .io_field_mean_ax(NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ax),
    .io_field_mean_bv(NV_NVDLA_CDMA_dual_reg_1_io_field_mean_bv),
    .io_field_conv_mode(NV_NVDLA_CDMA_dual_reg_1_io_field_conv_mode),
    .io_field_data_reuse(NV_NVDLA_CDMA_dual_reg_1_io_field_data_reuse),
    .io_field_in_precision(NV_NVDLA_CDMA_dual_reg_1_io_field_in_precision),
    .io_field_proc_precision(NV_NVDLA_CDMA_dual_reg_1_io_field_proc_precision),
    .io_field_skip_data_rls(NV_NVDLA_CDMA_dual_reg_1_io_field_skip_data_rls),
    .io_field_skip_weight_rls(NV_NVDLA_CDMA_dual_reg_1_io_field_skip_weight_rls),
    .io_field_weight_reuse(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_reuse),
    .io_field_nan_to_zero(NV_NVDLA_CDMA_dual_reg_1_io_field_nan_to_zero),
    .io_field_dma_en(NV_NVDLA_CDMA_dual_reg_1_io_field_dma_en),
    .io_field_pixel_x_offset(NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_x_offset),
    .io_field_pixel_y_offset(NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_y_offset),
    .io_field_rsv_per_line(NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_per_line),
    .io_field_rsv_per_uv_line(NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_per_uv_line),
    .io_field_rsv_height(NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_height),
    .io_field_rsv_y_index(NV_NVDLA_CDMA_dual_reg_1_io_field_rsv_y_index),
    .io_field_surf_stride(NV_NVDLA_CDMA_dual_reg_1_io_field_surf_stride),
    .io_field_weight_addr_high(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_high),
    .io_field_weight_addr_low(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_low),
    .io_field_weight_bytes(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bytes),
    .io_field_weight_format(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_format),
    .io_field_weight_ram_type(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_ram_type),
    .io_field_byte_per_kernel(NV_NVDLA_CDMA_dual_reg_1_io_field_byte_per_kernel),
    .io_field_weight_kernel(NV_NVDLA_CDMA_dual_reg_1_io_field_weight_kernel),
    .io_field_wgs_addr_high(NV_NVDLA_CDMA_dual_reg_1_io_field_wgs_addr_high),
    .io_field_wgs_addr_low(NV_NVDLA_CDMA_dual_reg_1_io_field_wgs_addr_low),
    .io_field_wmb_addr_high(NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_addr_high),
    .io_field_wmb_addr_low(NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_addr_low),
    .io_field_wmb_bytes(NV_NVDLA_CDMA_dual_reg_1_io_field_wmb_bytes),
    .io_field_pad_bottom(NV_NVDLA_CDMA_dual_reg_1_io_field_pad_bottom),
    .io_field_pad_left(NV_NVDLA_CDMA_dual_reg_1_io_field_pad_left),
    .io_field_pad_right(NV_NVDLA_CDMA_dual_reg_1_io_field_pad_right),
    .io_field_pad_top(NV_NVDLA_CDMA_dual_reg_1_io_field_pad_top),
    .io_field_pad_value(NV_NVDLA_CDMA_dual_reg_1_io_field_pad_value),
    .io_op_en_trigger(NV_NVDLA_CDMA_dual_reg_1_io_op_en_trigger),
    .io_inf_data_num(NV_NVDLA_CDMA_dual_reg_1_io_inf_data_num),
    .io_inf_weight_num(NV_NVDLA_CDMA_dual_reg_1_io_inf_weight_num),
    .io_nan_data_num(NV_NVDLA_CDMA_dual_reg_1_io_nan_data_num),
    .io_nan_weight_num(NV_NVDLA_CDMA_dual_reg_1_io_nan_weight_num),
    .io_op_en(NV_NVDLA_CDMA_dual_reg_1_io_op_en),
    .io_dat_rd_latency(NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_latency),
    .io_dat_rd_stall(NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_stall),
    .io_wt_rd_latency(NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_latency),
    .io_wt_rd_stall(NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_stall)
  );
  NV_NVDLA_CSB_LOGIC NV_NVDLA_CSB_LOGIC ( // @[NV_NVDLA_CDMA_regfile.scala 224:27:@1694.4]
    .reset(NV_NVDLA_CSB_LOGIC_reset),
    .io_clk(NV_NVDLA_CSB_LOGIC_io_clk),
    .io_csb2dp_req_valid(NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid),
    .io_csb2dp_req_bits(NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits),
    .io_csb2dp_resp_valid(NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid),
    .io_csb2dp_resp_bits(NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits),
    .io_reg_rd_data(NV_NVDLA_CSB_LOGIC_io_reg_rd_data),
    .io_reg_offset(NV_NVDLA_CSB_LOGIC_io_reg_offset),
    .io_reg_wr_data(NV_NVDLA_CSB_LOGIC_io_reg_wr_data),
    .io_reg_wr_en(NV_NVDLA_CSB_LOGIC_io_reg_wr_en)
  );
  assign _T_275 = ~ _T_203; // @[NV_NVDLA_CDMA_regfile.scala 156:33:@1607.4]
  assign _GEN_0 = io_dp2reg_done ? _T_275 : _T_203; // @[NV_NVDLA_CDMA_regfile.scala 158:25:@1608.4]
  assign _T_277 = _T_221 == 1'h0; // @[NV_NVDLA_CDMA_regfile.scala 169:44:@1612.4]
  assign _T_283 = _T_203 ? 2'h2 : 2'h1; // @[NV_NVDLA_CDMA_regfile.scala 170:27:@1614.4]
  assign _T_284 = _T_277 ? 2'h0 : _T_283; // @[NV_NVDLA_CDMA_regfile.scala 169:27:@1615.4]
  assign _T_286 = _T_250 == 1'h0; // @[NV_NVDLA_CDMA_regfile.scala 173:44:@1617.4]
  assign _T_289 = _T_203 == 1'h0; // @[NV_NVDLA_CDMA_regfile.scala 174:48:@1618.4]
  assign _T_292 = _T_289 ? 2'h2 : 2'h1; // @[NV_NVDLA_CDMA_regfile.scala 174:27:@1619.4]
  assign _T_293 = _T_286 ? 2'h0 : _T_292; // @[NV_NVDLA_CDMA_regfile.scala 173:27:@1620.4]
  assign _T_297 = ~ _T_221; // @[NV_NVDLA_CDMA_regfile.scala 183:33:@1623.4]
  assign _T_298 = _T_297 & NV_NVDLA_CDMA_dual_reg_io_op_en_trigger; // @[NV_NVDLA_CDMA_regfile.scala 183:50:@1624.4]
  assign _T_210 = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 72:27:@1538.4 NV_NVDLA_CDMA_regfile.scala 229:17:@1705.4]
  assign _T_299 = _T_210[0]; // @[NV_NVDLA_CDMA_regfile.scala 183:88:@1625.4]
  assign _T_302 = io_dp2reg_done & _T_289; // @[NV_NVDLA_CDMA_regfile.scala 184:48:@1627.4]
  assign _T_304 = _T_302 ? 1'h0 : _T_221; // @[NV_NVDLA_CDMA_regfile.scala 184:32:@1628.4]
  assign _T_305 = _T_298 ? _T_299 : _T_304; // @[NV_NVDLA_CDMA_regfile.scala 183:32:@1629.4]
  assign _T_306 = ~ _T_250; // @[NV_NVDLA_CDMA_regfile.scala 188:34:@1631.4]
  assign _T_307 = _T_306 & NV_NVDLA_CDMA_dual_reg_1_io_op_en_trigger; // @[NV_NVDLA_CDMA_regfile.scala 188:51:@1632.4]
  assign _T_311 = io_dp2reg_done & _T_203; // @[NV_NVDLA_CDMA_regfile.scala 189:49:@1635.4]
  assign _T_313 = _T_311 ? 1'h0 : _T_250; // @[NV_NVDLA_CDMA_regfile.scala 189:33:@1636.4]
  assign _T_314 = _T_307 ? _T_299 : _T_313; // @[NV_NVDLA_CDMA_regfile.scala 188:33:@1637.4]
  assign _T_315 = _T_203 ? _T_250 : _T_221; // @[NV_NVDLA_CDMA_regfile.scala 193:31:@1639.4]
  assign _T_317 = _T_296[1:0]; // @[NV_NVDLA_CDMA_regfile.scala 194:89:@1640.4]
  assign _T_318 = {_T_317,_T_315}; // @[Cat.scala 30:58:@1641.4]
  assign _T_319 = io_dp2reg_done ? 3'h0 : _T_318; // @[NV_NVDLA_CDMA_regfile.scala 194:33:@1642.4]
  assign _T_208 = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 71:26:@1537.4 NV_NVDLA_CDMA_regfile.scala 227:16:@1703.4]
  assign _GEN_20 = {{20'd0}, _T_208}; // @[NV_NVDLA_CDMA_regfile.scala 207:41:@1663.4]
  assign _T_336 = _GEN_20 < 32'h10; // @[NV_NVDLA_CDMA_regfile.scala 207:41:@1663.4]
  assign _T_342 = _GEN_20 >= 32'h10; // @[NV_NVDLA_CDMA_regfile.scala 208:39:@1666.4]
  assign _T_344 = NV_NVDLA_CDMA_single_reg_io_producer == 1'h0; // @[NV_NVDLA_CDMA_regfile.scala 208:83:@1667.4]
  assign _T_345 = _T_342 & _T_344; // @[NV_NVDLA_CDMA_regfile.scala 208:64:@1668.4]
  assign _T_350 = NV_NVDLA_CDMA_single_reg_io_producer; // @[NV_NVDLA_CDMA_regfile.scala 209:83:@1671.4]
  assign _T_351 = _T_342 & _T_350; // @[NV_NVDLA_CDMA_regfile.scala 209:64:@1672.4]
  assign _T_333 = NV_NVDLA_CSB_LOGIC_io_reg_wr_en; // @[NV_NVDLA_CDMA_regfile.scala 206:25:@1661.4 NV_NVDLA_CDMA_regfile.scala 228:15:@1704.4]
  assign _T_353 = _T_333 & _T_345; // @[NV_NVDLA_CDMA_regfile.scala 212:31:@1675.4]
  assign _T_357 = _T_333 & _T_351; // @[NV_NVDLA_CDMA_regfile.scala 213:31:@1679.4]
  assign _T_364 = _T_336 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@1684.4]
  assign _T_365 = _T_364 & NV_NVDLA_CDMA_single_reg_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 215:43:@1685.4]
  assign _T_369 = _T_345 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@1687.4]
  assign _T_370 = _T_369 & NV_NVDLA_CDMA_dual_reg_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 216:44:@1688.4]
  assign _T_371 = _T_365 | _T_370; // @[NV_NVDLA_CDMA_regfile.scala 215:59:@1689.4]
  assign _T_375 = _T_351 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@1691.4]
  assign _T_376 = _T_375 & NV_NVDLA_CDMA_dual_reg_1_io_reg_rd_data; // @[NV_NVDLA_CDMA_regfile.scala 217:43:@1692.4]
  assign _T_448 = io_dp2reg_wt_flush_done & io_dp2reg_dat_flush_done; // @[NV_NVDLA_CDMA_regfile.scala 251:50:@1777.4]
  assign _T_449 = ~ _T_305; // @[NV_NVDLA_CDMA_regfile.scala 256:43:@1779.4]
  assign _T_450 = _T_221 & _T_449; // @[NV_NVDLA_CDMA_regfile.scala 256:41:@1780.4]
  assign _T_452 = _T_297 & _T_305; // @[NV_NVDLA_CDMA_regfile.scala 257:42:@1782.4]
  assign _T_453 = _T_221 ^ _T_305; // @[NV_NVDLA_CDMA_regfile.scala 258:41:@1783.4]
  assign _T_454 = ~ _T_314; // @[NV_NVDLA_CDMA_regfile.scala 260:43:@1784.4]
  assign _T_455 = _T_250 & _T_454; // @[NV_NVDLA_CDMA_regfile.scala 260:41:@1785.4]
  assign _T_457 = _T_306 & _T_314; // @[NV_NVDLA_CDMA_regfile.scala 261:42:@1787.4]
  assign _T_458 = _T_250 ^ _T_314; // @[NV_NVDLA_CDMA_regfile.scala 262:41:@1788.4]
  assign _T_460 = _T_452 ? 32'h0 : _T_233; // @[NV_NVDLA_CDMA_regfile.scala 269:41:@1789.4]
  assign _T_461 = _T_450 ? 32'h0 : _T_460; // @[NV_NVDLA_CDMA_regfile.scala 268:41:@1790.4]
  assign _T_463 = _T_452 ? 32'h0 : _T_227; // @[NV_NVDLA_CDMA_regfile.scala 272:41:@1791.4]
  assign _T_464 = _T_450 ? 32'h0 : _T_463; // @[NV_NVDLA_CDMA_regfile.scala 271:41:@1792.4]
  assign _T_466 = _T_452 ? 32'h0 : _T_230; // @[NV_NVDLA_CDMA_regfile.scala 275:41:@1793.4]
  assign _T_467 = _T_450 ? 32'h0 : _T_466; // @[NV_NVDLA_CDMA_regfile.scala 274:39:@1794.4]
  assign _T_469 = _T_452 ? 32'h0 : _T_224; // @[NV_NVDLA_CDMA_regfile.scala 278:41:@1795.4]
  assign _T_470 = _T_450 ? 32'h0 : _T_469; // @[NV_NVDLA_CDMA_regfile.scala 277:39:@1796.4]
  assign _GEN_4 = _T_453 ? _T_461 : _T_233; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  assign _GEN_5 = _T_453 ? _T_464 : _T_227; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  assign _GEN_6 = _T_453 ? _T_467 : _T_230; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  assign _GEN_7 = _T_453 ? _T_470 : _T_224; // @[NV_NVDLA_CDMA_regfile.scala 281:24:@1797.4]
  assign _T_472 = _T_457 ? 32'h0 : _T_262; // @[NV_NVDLA_CDMA_regfile.scala 290:41:@1803.4]
  assign _T_473 = _T_455 ? 32'h0 : _T_472; // @[NV_NVDLA_CDMA_regfile.scala 289:41:@1804.4]
  assign _T_475 = _T_457 ? 32'h0 : _T_256; // @[NV_NVDLA_CDMA_regfile.scala 293:41:@1805.4]
  assign _T_476 = _T_455 ? 32'h0 : _T_475; // @[NV_NVDLA_CDMA_regfile.scala 292:41:@1806.4]
  assign _T_478 = _T_457 ? 32'h0 : _T_259; // @[NV_NVDLA_CDMA_regfile.scala 296:41:@1807.4]
  assign _T_479 = _T_455 ? 32'h0 : _T_478; // @[NV_NVDLA_CDMA_regfile.scala 295:39:@1808.4]
  assign _T_481 = _T_457 ? 32'h0 : _T_253; // @[NV_NVDLA_CDMA_regfile.scala 299:41:@1809.4]
  assign _T_482 = _T_455 ? 32'h0 : _T_481; // @[NV_NVDLA_CDMA_regfile.scala 298:39:@1810.4]
  assign _GEN_8 = _T_458 ? _T_473 : _T_262; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  assign _GEN_9 = _T_458 ? _T_476 : _T_256; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  assign _GEN_10 = _T_458 ? _T_479 : _T_259; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  assign _GEN_11 = _T_458 ? _T_482 : _T_253; // @[NV_NVDLA_CDMA_regfile.scala 302:24:@1811.4]
  assign _T_484 = _T_452 ? 32'h0 : _T_245; // @[NV_NVDLA_CDMA_regfile.scala 314:41:@1817.4]
  assign _T_485 = _T_450 ? io_dp2reg_wt_rd_stall : _T_484; // @[NV_NVDLA_CDMA_regfile.scala 313:38:@1818.4]
  assign _T_487 = _T_452 ? 32'h0 : _T_242; // @[NV_NVDLA_CDMA_regfile.scala 317:41:@1819.4]
  assign _T_488 = _T_450 ? 32'h0 : _T_487; // @[NV_NVDLA_CDMA_regfile.scala 316:40:@1820.4]
  assign _T_490 = io_dp2reg_dc_rd_stall | io_dp2reg_img_rd_stall; // @[NV_NVDLA_CDMA_regfile.scala 319:102:@1822.4]
  assign _T_492 = _T_452 ? 32'h0 : _T_239; // @[NV_NVDLA_CDMA_regfile.scala 320:41:@1823.4]
  assign _T_493 = _T_450 ? _T_490 : _T_492; // @[NV_NVDLA_CDMA_regfile.scala 319:39:@1824.4]
  assign _T_495 = io_dp2reg_dc_rd_latency | io_dp2reg_img_rd_latency; // @[NV_NVDLA_CDMA_regfile.scala 322:108:@1826.4]
  assign _T_497 = _T_452 ? 32'h0 : _T_236; // @[NV_NVDLA_CDMA_regfile.scala 323:41:@1827.4]
  assign _T_498 = _T_450 ? _T_495 : _T_497; // @[NV_NVDLA_CDMA_regfile.scala 322:41:@1828.4]
  assign _GEN_12 = _T_453 ? _T_485 : _T_245; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  assign _GEN_13 = _T_453 ? _T_488 : _T_242; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  assign _GEN_14 = _T_453 ? _T_493 : _T_239; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  assign _GEN_15 = _T_453 ? _T_498 : _T_236; // @[NV_NVDLA_CDMA_regfile.scala 326:24:@1829.4]
  assign _T_500 = _T_457 ? 32'h0 : _T_274; // @[NV_NVDLA_CDMA_regfile.scala 334:41:@1835.4]
  assign _T_501 = _T_455 ? io_dp2reg_wt_rd_stall : _T_500; // @[NV_NVDLA_CDMA_regfile.scala 333:38:@1836.4]
  assign _T_503 = _T_457 ? 32'h0 : _T_271; // @[NV_NVDLA_CDMA_regfile.scala 337:41:@1837.4]
  assign _T_504 = _T_455 ? 32'h0 : _T_503; // @[NV_NVDLA_CDMA_regfile.scala 336:40:@1838.4]
  assign _T_508 = _T_457 ? 32'h0 : _T_268; // @[NV_NVDLA_CDMA_regfile.scala 340:41:@1841.4]
  assign _T_509 = _T_455 ? _T_490 : _T_508; // @[NV_NVDLA_CDMA_regfile.scala 339:39:@1842.4]
  assign _T_513 = _T_457 ? 32'h0 : _T_265; // @[NV_NVDLA_CDMA_regfile.scala 343:41:@1845.4]
  assign _T_514 = _T_455 ? _T_495 : _T_513; // @[NV_NVDLA_CDMA_regfile.scala 342:41:@1846.4]
  assign _GEN_16 = _T_458 ? _T_501 : _T_274; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  assign _GEN_17 = _T_458 ? _T_504 : _T_271; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  assign _GEN_18 = _T_458 ? _T_509 : _T_268; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  assign _GEN_19 = _T_458 ? _T_514 : _T_265; // @[NV_NVDLA_CDMA_regfile.scala 346:24:@1847.4]
  assign _T_214 = _T_284[0]; // @[NV_NVDLA_CDMA_regfile.scala 74:31:@1540.4 NV_NVDLA_CDMA_regfile.scala 169:21:@1616.4]
  assign _T_216 = _T_293[0]; // @[NV_NVDLA_CDMA_regfile.scala 75:31:@1541.4 NV_NVDLA_CDMA_regfile.scala 173:21:@1621.4]
  assign io_csb2cdma_resp_valid = NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_valid; // @[NV_NVDLA_CDMA_regfile.scala 226:25:@1699.4]
  assign io_csb2cdma_resp_bits = NV_NVDLA_CSB_LOGIC_io_csb2dp_resp_bits; // @[NV_NVDLA_CDMA_regfile.scala 226:25:@1698.4]
  assign io_dp2reg_consumer = _T_203; // @[NV_NVDLA_CDMA_regfile.scala 162:24:@1611.4]
  assign io_reg2dp_field_data_bank = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_data_bank : NV_NVDLA_CDMA_dual_reg_io_field_data_bank; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1776.4]
  assign io_reg2dp_field_weight_bank = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bank : NV_NVDLA_CDMA_dual_reg_io_field_weight_bank; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1775.4]
  assign io_reg2dp_field_batches = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_batches : NV_NVDLA_CDMA_dual_reg_io_field_batches; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1774.4]
  assign io_reg2dp_field_batch_stride = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_batch_stride : NV_NVDLA_CDMA_dual_reg_io_field_batch_stride; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1773.4]
  assign io_reg2dp_field_cvt_en = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_en : NV_NVDLA_CDMA_dual_reg_io_field_cvt_en; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1770.4]
  assign io_reg2dp_field_cvt_truncate = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_truncate : NV_NVDLA_CDMA_dual_reg_io_field_cvt_truncate; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1769.4]
  assign io_reg2dp_field_cvt_offset = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_offset : NV_NVDLA_CDMA_dual_reg_io_field_cvt_offset; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1768.4]
  assign io_reg2dp_field_cvt_scale = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_cvt_scale : NV_NVDLA_CDMA_dual_reg_io_field_cvt_scale; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1767.4]
  assign io_reg2dp_field_datain_addr_high_0 = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_0 : NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_0; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1765.4]
  assign io_reg2dp_field_datain_addr_high_1 = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_high_1 : NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_high_1; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1764.4]
  assign io_reg2dp_field_datain_addr_low_0 = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_0 : NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_0; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1763.4]
  assign io_reg2dp_field_datain_addr_low_1 = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_addr_low_1 : NV_NVDLA_CDMA_dual_reg_io_field_datain_addr_low_1; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1762.4]
  assign io_reg2dp_field_line_packed = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_line_packed : NV_NVDLA_CDMA_dual_reg_io_field_line_packed; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1761.4]
  assign io_reg2dp_field_surf_packed = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_surf_packed : NV_NVDLA_CDMA_dual_reg_io_field_surf_packed; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1760.4]
  assign io_reg2dp_field_datain_ram_type = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_ram_type : NV_NVDLA_CDMA_dual_reg_io_field_datain_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1759.4]
  assign io_reg2dp_field_datain_format = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_format : NV_NVDLA_CDMA_dual_reg_io_field_datain_format; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1758.4]
  assign io_reg2dp_field_pixel_format = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_format : NV_NVDLA_CDMA_dual_reg_io_field_pixel_format; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1757.4]
  assign io_reg2dp_field_pixel_sign_override = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_sign_override : NV_NVDLA_CDMA_dual_reg_io_field_pixel_sign_override; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1755.4]
  assign io_reg2dp_field_datain_height = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_height : NV_NVDLA_CDMA_dual_reg_io_field_datain_height; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1754.4]
  assign io_reg2dp_field_datain_width = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_width : NV_NVDLA_CDMA_dual_reg_io_field_datain_width; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1753.4]
  assign io_reg2dp_field_datain_channel = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_datain_channel : NV_NVDLA_CDMA_dual_reg_io_field_datain_channel; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1752.4]
  assign io_reg2dp_field_entries = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_entries : NV_NVDLA_CDMA_dual_reg_io_field_entries; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1749.4]
  assign io_reg2dp_field_grains = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_grains : NV_NVDLA_CDMA_dual_reg_io_field_grains; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1748.4]
  assign io_reg2dp_field_line_stride = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_line_stride : NV_NVDLA_CDMA_dual_reg_io_field_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1747.4]
  assign io_reg2dp_field_uv_line_stride = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_uv_line_stride : NV_NVDLA_CDMA_dual_reg_io_field_uv_line_stride; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1746.4]
  assign io_reg2dp_field_mean_format = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_mean_format : NV_NVDLA_CDMA_dual_reg_io_field_mean_format; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1745.4]
  assign io_reg2dp_field_mean_gu = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_mean_gu : NV_NVDLA_CDMA_dual_reg_io_field_mean_gu; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1744.4]
  assign io_reg2dp_field_mean_ry = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ry : NV_NVDLA_CDMA_dual_reg_io_field_mean_ry; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1743.4]
  assign io_reg2dp_field_mean_ax = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_mean_ax : NV_NVDLA_CDMA_dual_reg_io_field_mean_ax; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1742.4]
  assign io_reg2dp_field_mean_bv = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_mean_bv : NV_NVDLA_CDMA_dual_reg_io_field_mean_bv; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1741.4]
  assign io_reg2dp_field_conv_mode = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_conv_mode : NV_NVDLA_CDMA_dual_reg_io_field_conv_mode; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1740.4]
  assign io_reg2dp_field_data_reuse = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_data_reuse : NV_NVDLA_CDMA_dual_reg_io_field_data_reuse; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1739.4]
  assign io_reg2dp_field_proc_precision = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_proc_precision : NV_NVDLA_CDMA_dual_reg_io_field_proc_precision; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1737.4]
  assign io_reg2dp_field_skip_data_rls = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_skip_data_rls : NV_NVDLA_CDMA_dual_reg_io_field_skip_data_rls; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1736.4]
  assign io_reg2dp_field_skip_weight_rls = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_skip_weight_rls : NV_NVDLA_CDMA_dual_reg_io_field_skip_weight_rls; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1735.4]
  assign io_reg2dp_field_weight_reuse = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_reuse : NV_NVDLA_CDMA_dual_reg_io_field_weight_reuse; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1734.4]
  assign io_reg2dp_field_dma_en = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_dma_en : NV_NVDLA_CDMA_dual_reg_io_field_dma_en; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1732.4]
  assign io_reg2dp_field_pixel_x_offset = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pixel_x_offset : NV_NVDLA_CDMA_dual_reg_io_field_pixel_x_offset; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1731.4]
  assign io_reg2dp_field_surf_stride = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_surf_stride : NV_NVDLA_CDMA_dual_reg_io_field_surf_stride; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1725.4]
  assign io_reg2dp_field_weight_addr_high = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_high : NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_high; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1724.4]
  assign io_reg2dp_field_weight_addr_low = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_addr_low : NV_NVDLA_CDMA_dual_reg_io_field_weight_addr_low; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1723.4]
  assign io_reg2dp_field_weight_bytes = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_bytes : NV_NVDLA_CDMA_dual_reg_io_field_weight_bytes; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1722.4]
  assign io_reg2dp_field_weight_ram_type = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_ram_type : NV_NVDLA_CDMA_dual_reg_io_field_weight_ram_type; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1720.4]
  assign io_reg2dp_field_byte_per_kernel = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_byte_per_kernel : NV_NVDLA_CDMA_dual_reg_io_field_byte_per_kernel; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1719.4]
  assign io_reg2dp_field_weight_kernel = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_weight_kernel : NV_NVDLA_CDMA_dual_reg_io_field_weight_kernel; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1718.4]
  assign io_reg2dp_field_pad_left = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pad_left : NV_NVDLA_CDMA_dual_reg_io_field_pad_left; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1711.4]
  assign io_reg2dp_field_pad_right = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pad_right : NV_NVDLA_CDMA_dual_reg_io_field_pad_right; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1710.4]
  assign io_reg2dp_field_pad_value = _T_203 ? NV_NVDLA_CDMA_dual_reg_1_io_field_pad_value : NV_NVDLA_CDMA_dual_reg_io_field_pad_value; // @[NV_NVDLA_CDMA_regfile.scala 237:21:@1708.4]
  assign io_reg2dp_op_en = _T_296[2]; // @[NV_NVDLA_CDMA_regfile.scala 197:21:@1645.4]
  assign NV_NVDLA_CDMA_single_reg_clock = io_nvdla_core_clk; // @[:@1543.4]
  assign NV_NVDLA_CDMA_single_reg_reset = reset; // @[:@1544.4]
  assign NV_NVDLA_CDMA_single_reg_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 80:32:@1546.4]
  assign NV_NVDLA_CDMA_single_reg_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 81:33:@1547.4]
  assign NV_NVDLA_CDMA_single_reg_io_reg_wr_en = _T_333 & _T_336; // @[NV_NVDLA_CDMA_regfile.scala 82:31:@1548.4]
  assign NV_NVDLA_CDMA_single_reg_io_flush_done = _T_206; // @[NV_NVDLA_CDMA_regfile.scala 83:32:@1549.4]
  assign NV_NVDLA_CDMA_single_reg_io_consumer = _T_203; // @[NV_NVDLA_CDMA_regfile.scala 84:30:@1550.4]
  assign NV_NVDLA_CDMA_single_reg_io_status_0 = {{1'd0}, _T_214}; // @[NV_NVDLA_CDMA_regfile.scala 85:30:@1551.4]
  assign NV_NVDLA_CDMA_single_reg_io_status_1 = {{1'd0}, _T_216}; // @[NV_NVDLA_CDMA_regfile.scala 86:30:@1552.4]
  assign NV_NVDLA_CDMA_dual_reg_reset = reset; // @[:@1567.4]
  assign NV_NVDLA_CDMA_dual_reg_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_regfile.scala 105:37:@1568.4]
  assign NV_NVDLA_CDMA_dual_reg_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 106:33:@1569.4]
  assign NV_NVDLA_CDMA_dual_reg_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 107:34:@1570.4]
  assign NV_NVDLA_CDMA_dual_reg_io_reg_wr_en = _T_353 & _T_277; // @[NV_NVDLA_CDMA_regfile.scala 108:32:@1571.4]
  assign NV_NVDLA_CDMA_dual_reg_io_inf_data_num = _T_224; // @[NV_NVDLA_CDMA_regfile.scala 111:35:@1573.4]
  assign NV_NVDLA_CDMA_dual_reg_io_inf_weight_num = _T_227; // @[NV_NVDLA_CDMA_regfile.scala 112:37:@1574.4]
  assign NV_NVDLA_CDMA_dual_reg_io_nan_data_num = _T_230; // @[NV_NVDLA_CDMA_regfile.scala 113:35:@1575.4]
  assign NV_NVDLA_CDMA_dual_reg_io_nan_weight_num = _T_233; // @[NV_NVDLA_CDMA_regfile.scala 114:37:@1576.4]
  assign NV_NVDLA_CDMA_dual_reg_io_op_en = _T_221; // @[NV_NVDLA_CDMA_regfile.scala 110:28:@1572.4]
  assign NV_NVDLA_CDMA_dual_reg_io_dat_rd_latency = _T_236; // @[NV_NVDLA_CDMA_regfile.scala 115:37:@1577.4]
  assign NV_NVDLA_CDMA_dual_reg_io_dat_rd_stall = _T_239; // @[NV_NVDLA_CDMA_regfile.scala 116:35:@1578.4]
  assign NV_NVDLA_CDMA_dual_reg_io_wt_rd_latency = _T_242; // @[NV_NVDLA_CDMA_regfile.scala 117:36:@1579.4]
  assign NV_NVDLA_CDMA_dual_reg_io_wt_rd_stall = _T_245; // @[NV_NVDLA_CDMA_regfile.scala 118:34:@1580.4]
  assign NV_NVDLA_CDMA_dual_reg_1_reset = reset; // @[:@1593.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_regfile.scala 134:37:@1594.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_reg_offset = NV_NVDLA_CSB_LOGIC_io_reg_offset; // @[NV_NVDLA_CDMA_regfile.scala 135:33:@1595.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_data = NV_NVDLA_CSB_LOGIC_io_reg_wr_data; // @[NV_NVDLA_CDMA_regfile.scala 136:34:@1596.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_reg_wr_en = _T_357 & _T_286; // @[NV_NVDLA_CDMA_regfile.scala 137:32:@1597.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_inf_data_num = _T_253; // @[NV_NVDLA_CDMA_regfile.scala 140:35:@1599.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_inf_weight_num = _T_256; // @[NV_NVDLA_CDMA_regfile.scala 141:37:@1600.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_nan_data_num = _T_259; // @[NV_NVDLA_CDMA_regfile.scala 142:35:@1601.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_nan_weight_num = _T_262; // @[NV_NVDLA_CDMA_regfile.scala 143:37:@1602.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_op_en = _T_250; // @[NV_NVDLA_CDMA_regfile.scala 139:28:@1598.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_latency = _T_265; // @[NV_NVDLA_CDMA_regfile.scala 144:37:@1603.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_dat_rd_stall = _T_268; // @[NV_NVDLA_CDMA_regfile.scala 145:35:@1604.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_latency = _T_271; // @[NV_NVDLA_CDMA_regfile.scala 146:36:@1605.4]
  assign NV_NVDLA_CDMA_dual_reg_1_io_wt_rd_stall = _T_274; // @[NV_NVDLA_CDMA_regfile.scala 147:34:@1606.4]
  assign NV_NVDLA_CSB_LOGIC_reset = reset; // @[:@1696.4]
  assign NV_NVDLA_CSB_LOGIC_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_regfile.scala 225:22:@1697.4]
  assign NV_NVDLA_CSB_LOGIC_io_csb2dp_req_valid = io_csb2cdma_req_valid; // @[NV_NVDLA_CDMA_regfile.scala 226:25:@1701.4]
  assign NV_NVDLA_CSB_LOGIC_io_csb2dp_req_bits = io_csb2cdma_req_bits; // @[NV_NVDLA_CDMA_regfile.scala 226:25:@1700.4]
  assign NV_NVDLA_CSB_LOGIC_io_reg_rd_data = _T_371 | _T_376; // @[NV_NVDLA_CDMA_regfile.scala 230:30:@1706.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_203 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_206 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_221 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_224 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_227 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_230 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_233 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_236 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_239 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_242 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_245 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_250 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_253 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_256 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_259 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_262 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_265 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_268 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_271 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_274 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_296 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_203 <= 1'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_203 <= _T_275;
      end
    end
    if (reset) begin
      _T_206 <= 1'h0;
    end else begin
      _T_206 <= _T_448;
    end
    if (reset) begin
      _T_221 <= 1'h0;
    end else begin
      if (_T_298) begin
        _T_221 <= _T_299;
      end else begin
        if (_T_302) begin
          _T_221 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_224 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_224 <= 32'h0;
        end else begin
          if (_T_452) begin
            _T_224 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_227 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_227 <= 32'h0;
        end else begin
          if (_T_452) begin
            _T_227 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_230 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_230 <= 32'h0;
        end else begin
          if (_T_452) begin
            _T_230 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_233 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_233 <= 32'h0;
        end else begin
          if (_T_452) begin
            _T_233 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_236 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_236 <= _T_495;
        end else begin
          if (_T_452) begin
            _T_236 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_239 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_239 <= _T_490;
        end else begin
          if (_T_452) begin
            _T_239 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_242 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_242 <= 32'h0;
        end else begin
          if (_T_452) begin
            _T_242 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_245 <= 32'h0;
    end else begin
      if (_T_453) begin
        if (_T_450) begin
          _T_245 <= io_dp2reg_wt_rd_stall;
        end else begin
          if (_T_452) begin
            _T_245 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_250 <= 1'h0;
    end else begin
      if (_T_307) begin
        _T_250 <= _T_299;
      end else begin
        if (_T_311) begin
          _T_250 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_253 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_253 <= 32'h0;
        end else begin
          if (_T_457) begin
            _T_253 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_256 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_256 <= 32'h0;
        end else begin
          if (_T_457) begin
            _T_256 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_259 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_259 <= 32'h0;
        end else begin
          if (_T_457) begin
            _T_259 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_262 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_262 <= 32'h0;
        end else begin
          if (_T_457) begin
            _T_262 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_265 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_265 <= _T_495;
        end else begin
          if (_T_457) begin
            _T_265 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_268 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_268 <= _T_490;
        end else begin
          if (_T_457) begin
            _T_268 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_271 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_271 <= 32'h0;
        end else begin
          if (_T_457) begin
            _T_271 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_274 <= 32'h0;
    end else begin
      if (_T_458) begin
        if (_T_455) begin
          _T_274 <= io_dp2reg_wt_rd_stall;
        end else begin
          if (_T_457) begin
            _T_274 <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_296 <= 3'h0;
    end else begin
      if (io_dp2reg_done) begin
        _T_296 <= 3'h0;
      end else begin
        _T_296 <= _T_318;
      end
    end
  end
endmodule
module NV_NVDLA_IS_pipe( // @[:@1854.2]
  input         reset, // @[:@1856.4]
  input         io_clk, // @[:@1857.4]
  output [78:0] io_dout, // @[:@1857.4]
  output        io_vo, // @[:@1857.4]
  input         io_ri, // @[:@1857.4]
  input  [78:0] io_di, // @[:@1857.4]
  input         io_vi, // @[:@1857.4]
  output        io_ro // @[:@1857.4]
);
  reg  _T_21; // @[IS_pipe.scala 53:25:@1859.4]
  reg [31:0] _RAND_0;
  reg  _T_24; // @[IS_pipe.scala 54:31:@1860.4]
  reg [31:0] _RAND_1;
  reg  _T_27; // @[IS_pipe.scala 55:31:@1861.4]
  reg [31:0] _RAND_2;
  reg [78:0] _T_29; // @[IS_pipe.scala 56:27:@1862.4]
  reg [95:0] _RAND_3;
  reg  _T_32; // @[IS_pipe.scala 57:31:@1863.4]
  reg [31:0] _RAND_4;
  reg [78:0] _T_34; // @[IS_pipe.scala 58:27:@1864.4]
  reg [95:0] _RAND_5;
  wire  _GEN_0; // @[IS_pipe.scala 70:23:@1873.4]
  wire  _T_48; // @[IS_pipe.scala 75:22:@1878.4]
  wire [78:0] _T_49; // @[IS_pipe.scala 78:19:@1882.4]
  wire  _T_51; // @[IS_pipe.scala 80:32:@1884.4]
  wire  _T_52; // @[IS_pipe.scala 80:29:@1885.4]
  wire  _GEN_2; // @[IS_pipe.scala 82:18:@1887.4]
  wire  _T_53; // @[IS_pipe.scala 86:18:@1890.4]
  assign _GEN_0 = _T_24 ? io_vi : _T_27; // @[IS_pipe.scala 70:23:@1873.4]
  assign _T_48 = _T_24 & io_vi; // @[IS_pipe.scala 75:22:@1878.4]
  assign _T_49 = _T_24 ? io_di : _T_29; // @[IS_pipe.scala 78:19:@1882.4]
  assign _T_51 = _T_32 == 1'h0; // @[IS_pipe.scala 80:32:@1884.4]
  assign _T_52 = io_ri | _T_51; // @[IS_pipe.scala 80:29:@1885.4]
  assign _GEN_2 = _T_52 ? _GEN_0 : _T_32; // @[IS_pipe.scala 82:18:@1887.4]
  assign _T_53 = _T_52 & _GEN_0; // @[IS_pipe.scala 86:18:@1890.4]
  assign io_dout = _T_34; // @[IS_pipe.scala 97:13:@1899.4]
  assign io_vo = _T_32; // @[IS_pipe.scala 96:11:@1898.4]
  assign io_ro = _T_21; // @[IS_pipe.scala 95:11:@1897.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_24 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_27 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  _T_29 = _RAND_3[78:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_32 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  _T_34 = _RAND_5[78:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_21 <= 1'h1;
    end else begin
      _T_21 <= _T_52;
    end
    if (reset) begin
      _T_24 <= 1'h1;
    end else begin
      _T_24 <= _T_52;
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_24) begin
        _T_27 <= io_vi;
      end
    end
    if (_T_48) begin
      _T_29 <= io_di;
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      if (_T_52) begin
        if (_T_24) begin
          _T_32 <= io_vi;
        end else begin
          _T_32 <= _T_27;
        end
      end
    end
    if (_T_53) begin
      if (_T_24) begin
        _T_34 <= io_di;
      end else begin
        _T_34 <= _T_29;
      end
    end
  end
endmodule
module NV_soDLA_DMAIF_rdreq( // @[:@1948.2]
  input         reset, // @[:@1950.4]
  input         io_nvdla_core_clk, // @[:@1951.4]
  output        io_dmaif_rd_req_pd_ready, // @[:@1951.4]
  input         io_dmaif_rd_req_pd_valid, // @[:@1951.4]
  input  [78:0] io_dmaif_rd_req_pd_bits, // @[:@1951.4]
  input         io_mcif_rd_req_pd_ready, // @[:@1951.4]
  output        io_mcif_rd_req_pd_valid, // @[:@1951.4]
  output [78:0] io_mcif_rd_req_pd_bits, // @[:@1951.4]
  input         io_cvif_rd_req_pd_ready, // @[:@1951.4]
  output        io_cvif_rd_req_pd_valid, // @[:@1951.4]
  output [78:0] io_cvif_rd_req_pd_bits, // @[:@1951.4]
  input         io_reg2dp_src_ram_type // @[:@1951.4]
);
  wire  NV_NVDLA_IS_pipe_reset; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_io_clk; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire [78:0] NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_io_vo; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_io_ri; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire [78:0] NV_NVDLA_IS_pipe_io_di; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_io_vi; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_io_ro; // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
  wire  NV_NVDLA_IS_pipe_1_reset; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  NV_NVDLA_IS_pipe_1_io_clk; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire [78:0] NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  NV_NVDLA_IS_pipe_1_io_vo; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  NV_NVDLA_IS_pipe_1_io_ri; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire [78:0] NV_NVDLA_IS_pipe_1_io_di; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  NV_NVDLA_IS_pipe_1_io_vi; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  NV_NVDLA_IS_pipe_1_io_ro; // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
  wire  _T_38; // @[NV_NVDLA_DMAIF_rdreq.scala 54:44:@1965.4]
  wire  _T_40; // @[NV_NVDLA_DMAIF_rdreq.scala 61:78:@1970.4]
  wire  _T_44; // @[NV_NVDLA_DMAIF_rdreq.scala 68:48:@1978.4]
  NV_NVDLA_IS_pipe NV_NVDLA_IS_pipe ( // @[NV_NVDLA_DMAIF_rdreq.scala 45:26:@1953.4]
    .reset(NV_NVDLA_IS_pipe_reset),
    .io_clk(NV_NVDLA_IS_pipe_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_io_ri),
    .io_di(NV_NVDLA_IS_pipe_io_di),
    .io_vi(NV_NVDLA_IS_pipe_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_io_ro)
  );
  NV_NVDLA_IS_pipe NV_NVDLA_IS_pipe_1 ( // @[NV_NVDLA_DMAIF_rdreq.scala 59:30:@1966.4]
    .reset(NV_NVDLA_IS_pipe_1_reset),
    .io_clk(NV_NVDLA_IS_pipe_1_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_1_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_1_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_1_io_ri),
    .io_di(NV_NVDLA_IS_pipe_1_io_di),
    .io_vi(NV_NVDLA_IS_pipe_1_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_1_io_ro)
  );
  assign _T_38 = NV_NVDLA_IS_pipe_io_ro & io_reg2dp_src_ram_type; // @[NV_NVDLA_DMAIF_rdreq.scala 54:44:@1965.4]
  assign _T_40 = io_reg2dp_src_ram_type == 1'h0; // @[NV_NVDLA_DMAIF_rdreq.scala 61:78:@1970.4]
  assign _T_44 = NV_NVDLA_IS_pipe_1_io_ro & _T_40; // @[NV_NVDLA_DMAIF_rdreq.scala 68:48:@1978.4]
  assign io_dmaif_rd_req_pd_ready = _T_38 | _T_44; // @[NV_NVDLA_DMAIF_rdreq.scala 69:34:@1980.4]
  assign io_mcif_rd_req_pd_valid = NV_NVDLA_IS_pipe_io_vo; // @[NV_NVDLA_DMAIF_rdreq.scala 50:29:@1961.4]
  assign io_mcif_rd_req_pd_bits = NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_DMAIF_rdreq.scala 52:28:@1963.4]
  assign io_cvif_rd_req_pd_valid = NV_NVDLA_IS_pipe_1_io_vo; // @[NV_NVDLA_DMAIF_rdreq.scala 64:37:@1974.4]
  assign io_cvif_rd_req_pd_bits = NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_DMAIF_rdreq.scala 66:36:@1976.4]
  assign NV_NVDLA_IS_pipe_reset = reset; // @[:@1955.4]
  assign NV_NVDLA_IS_pipe_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_DMAIF_rdreq.scala 46:21:@1956.4]
  assign NV_NVDLA_IS_pipe_io_ri = io_mcif_rd_req_pd_ready; // @[NV_NVDLA_DMAIF_rdreq.scala 51:20:@1962.4]
  assign NV_NVDLA_IS_pipe_io_di = io_dmaif_rd_req_pd_bits; // @[NV_NVDLA_DMAIF_rdreq.scala 49:20:@1960.4]
  assign NV_NVDLA_IS_pipe_io_vi = io_dmaif_rd_req_pd_valid & io_reg2dp_src_ram_type; // @[NV_NVDLA_DMAIF_rdreq.scala 47:20:@1959.4]
  assign NV_NVDLA_IS_pipe_1_reset = reset; // @[:@1968.4]
  assign NV_NVDLA_IS_pipe_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_DMAIF_rdreq.scala 60:25:@1969.4]
  assign NV_NVDLA_IS_pipe_1_io_ri = io_cvif_rd_req_pd_ready; // @[NV_NVDLA_DMAIF_rdreq.scala 65:24:@1975.4]
  assign NV_NVDLA_IS_pipe_1_io_di = io_dmaif_rd_req_pd_bits; // @[NV_NVDLA_DMAIF_rdreq.scala 63:24:@1973.4]
  assign NV_NVDLA_IS_pipe_1_io_vi = io_dmaif_rd_req_pd_valid & _T_40; // @[NV_NVDLA_DMAIF_rdreq.scala 61:24:@1972.4]
endmodule
module NV_NVDLA_IS_pipe_2( // @[:@1982.2]
  input          reset, // @[:@1984.4]
  input          io_clk, // @[:@1985.4]
  output [256:0] io_dout, // @[:@1985.4]
  output         io_vo, // @[:@1985.4]
  input          io_ri, // @[:@1985.4]
  input  [256:0] io_di, // @[:@1985.4]
  input          io_vi, // @[:@1985.4]
  output         io_ro // @[:@1985.4]
);
  reg  _T_21; // @[IS_pipe.scala 53:25:@1987.4]
  reg [31:0] _RAND_0;
  reg  _T_24; // @[IS_pipe.scala 54:31:@1988.4]
  reg [31:0] _RAND_1;
  reg  _T_27; // @[IS_pipe.scala 55:31:@1989.4]
  reg [31:0] _RAND_2;
  reg [256:0] _T_29; // @[IS_pipe.scala 56:27:@1990.4]
  reg [287:0] _RAND_3;
  reg  _T_32; // @[IS_pipe.scala 57:31:@1991.4]
  reg [31:0] _RAND_4;
  reg [256:0] _T_34; // @[IS_pipe.scala 58:27:@1992.4]
  reg [287:0] _RAND_5;
  wire  _GEN_0; // @[IS_pipe.scala 70:23:@2001.4]
  wire  _T_48; // @[IS_pipe.scala 75:22:@2006.4]
  wire [256:0] _T_49; // @[IS_pipe.scala 78:19:@2010.4]
  wire  _T_51; // @[IS_pipe.scala 80:32:@2012.4]
  wire  _T_52; // @[IS_pipe.scala 80:29:@2013.4]
  wire  _GEN_2; // @[IS_pipe.scala 82:18:@2015.4]
  wire  _T_53; // @[IS_pipe.scala 86:18:@2018.4]
  assign _GEN_0 = _T_24 ? io_vi : _T_27; // @[IS_pipe.scala 70:23:@2001.4]
  assign _T_48 = _T_24 & io_vi; // @[IS_pipe.scala 75:22:@2006.4]
  assign _T_49 = _T_24 ? io_di : _T_29; // @[IS_pipe.scala 78:19:@2010.4]
  assign _T_51 = _T_32 == 1'h0; // @[IS_pipe.scala 80:32:@2012.4]
  assign _T_52 = io_ri | _T_51; // @[IS_pipe.scala 80:29:@2013.4]
  assign _GEN_2 = _T_52 ? _GEN_0 : _T_32; // @[IS_pipe.scala 82:18:@2015.4]
  assign _T_53 = _T_52 & _GEN_0; // @[IS_pipe.scala 86:18:@2018.4]
  assign io_dout = _T_34; // @[IS_pipe.scala 97:13:@2027.4]
  assign io_vo = _T_32; // @[IS_pipe.scala 96:11:@2026.4]
  assign io_ro = _T_21; // @[IS_pipe.scala 95:11:@2025.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_24 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_27 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {9{`RANDOM}};
  _T_29 = _RAND_3[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_32 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {9{`RANDOM}};
  _T_34 = _RAND_5[256:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_21 <= 1'h1;
    end else begin
      _T_21 <= _T_52;
    end
    if (reset) begin
      _T_24 <= 1'h1;
    end else begin
      _T_24 <= _T_52;
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_24) begin
        _T_27 <= io_vi;
      end
    end
    if (_T_48) begin
      _T_29 <= io_di;
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      if (_T_52) begin
        if (_T_24) begin
          _T_32 <= io_vi;
        end else begin
          _T_32 <= _T_27;
        end
      end
    end
    if (_T_53) begin
      if (_T_24) begin
        _T_34 <= io_di;
      end else begin
        _T_34 <= _T_29;
      end
    end
  end
endmodule
module NV_soDLA_DMAIF_rdrsp( // @[:@2123.2]
  input          reset, // @[:@2125.4]
  input          io_nvdla_core_clk, // @[:@2126.4]
  output         io_mcif_rd_rsp_pd_ready, // @[:@2126.4]
  input          io_mcif_rd_rsp_pd_valid, // @[:@2126.4]
  input  [256:0] io_mcif_rd_rsp_pd_bits, // @[:@2126.4]
  output         io_cvif_rd_rsp_pd_ready, // @[:@2126.4]
  input          io_cvif_rd_rsp_pd_valid, // @[:@2126.4]
  input  [256:0] io_cvif_rd_rsp_pd_bits, // @[:@2126.4]
  input          io_dmaif_rd_rsp_pd_ready, // @[:@2126.4]
  output         io_dmaif_rd_rsp_pd_valid, // @[:@2126.4]
  output [256:0] io_dmaif_rd_rsp_pd_bits // @[:@2126.4]
);
  wire  NV_NVDLA_IS_pipe_reset; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_io_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire [256:0] NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_io_vo; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_io_ri; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire [256:0] NV_NVDLA_IS_pipe_io_di; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_io_vi; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
  wire  NV_NVDLA_IS_pipe_1_reset; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_1_io_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire [256:0] NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_1_io_vo; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_1_io_ri; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire [256:0] NV_NVDLA_IS_pipe_1_io_di; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_1_io_vi; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_1_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
  wire  NV_NVDLA_IS_pipe_2_reset; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  NV_NVDLA_IS_pipe_2_io_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire [256:0] NV_NVDLA_IS_pipe_2_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  NV_NVDLA_IS_pipe_2_io_vo; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  NV_NVDLA_IS_pipe_2_io_ri; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire [256:0] NV_NVDLA_IS_pipe_2_io_di; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  NV_NVDLA_IS_pipe_2_io_vi; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  NV_NVDLA_IS_pipe_2_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
  wire  _T_44; // @[Bitwise.scala 72:15:@2149.4]
  wire [256:0] _T_47; // @[Bitwise.scala 72:12:@2150.4]
  wire [256:0] _T_48; // @[NV_NVDLA_DMAIF_rdrsp.scala 71:61:@2151.4]
  wire  _T_49; // @[Bitwise.scala 72:15:@2152.4]
  wire [256:0] _T_52; // @[Bitwise.scala 72:12:@2153.4]
  wire [256:0] _T_53; // @[NV_NVDLA_DMAIF_rdrsp.scala 72:61:@2154.4]
  NV_NVDLA_IS_pipe_2 NV_NVDLA_IS_pipe ( // @[NV_NVDLA_DMAIF_rdrsp.scala 49:26:@2131.4]
    .reset(NV_NVDLA_IS_pipe_reset),
    .io_clk(NV_NVDLA_IS_pipe_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_io_ri),
    .io_di(NV_NVDLA_IS_pipe_io_di),
    .io_vi(NV_NVDLA_IS_pipe_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_io_ro)
  );
  NV_NVDLA_IS_pipe_2 NV_NVDLA_IS_pipe_1 ( // @[NV_NVDLA_DMAIF_rdrsp.scala 59:30:@2139.4]
    .reset(NV_NVDLA_IS_pipe_1_reset),
    .io_clk(NV_NVDLA_IS_pipe_1_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_1_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_1_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_1_io_ri),
    .io_di(NV_NVDLA_IS_pipe_1_io_di),
    .io_vi(NV_NVDLA_IS_pipe_1_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_1_io_ro)
  );
  NV_NVDLA_IS_pipe_2 NV_NVDLA_IS_pipe_2 ( // @[NV_NVDLA_DMAIF_rdrsp.scala 85:26:@2157.4]
    .reset(NV_NVDLA_IS_pipe_2_reset),
    .io_clk(NV_NVDLA_IS_pipe_2_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_2_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_2_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_2_io_ri),
    .io_di(NV_NVDLA_IS_pipe_2_io_di),
    .io_vi(NV_NVDLA_IS_pipe_2_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_2_io_ro)
  );
  assign _T_44 = NV_NVDLA_IS_pipe_io_vo; // @[Bitwise.scala 72:15:@2149.4]
  assign _T_47 = _T_44 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@2150.4]
  assign _T_48 = _T_47 & NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 71:61:@2151.4]
  assign _T_49 = NV_NVDLA_IS_pipe_1_io_vo; // @[Bitwise.scala 72:15:@2152.4]
  assign _T_52 = _T_49 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@2153.4]
  assign _T_53 = _T_52 & NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 72:61:@2154.4]
  assign io_mcif_rd_rsp_pd_ready = NV_NVDLA_IS_pipe_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 52:29:@2136.4]
  assign io_cvif_rd_rsp_pd_ready = NV_NVDLA_IS_pipe_1_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 62:37:@2144.4]
  assign io_dmaif_rd_rsp_pd_valid = NV_NVDLA_IS_pipe_2_io_vo; // @[NV_NVDLA_DMAIF_rdrsp.scala 90:30:@2164.4]
  assign io_dmaif_rd_rsp_pd_bits = NV_NVDLA_IS_pipe_2_io_dout; // @[NV_NVDLA_DMAIF_rdrsp.scala 92:28:@2166.4]
  assign NV_NVDLA_IS_pipe_reset = reset; // @[:@2133.4]
  assign NV_NVDLA_IS_pipe_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 50:21:@2134.4]
  assign NV_NVDLA_IS_pipe_io_ri = NV_NVDLA_IS_pipe_2_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 55:20:@2138.4]
  assign NV_NVDLA_IS_pipe_io_di = io_mcif_rd_rsp_pd_bits; // @[NV_NVDLA_DMAIF_rdrsp.scala 53:20:@2137.4]
  assign NV_NVDLA_IS_pipe_io_vi = io_mcif_rd_rsp_pd_valid; // @[NV_NVDLA_DMAIF_rdrsp.scala 51:20:@2135.4]
  assign NV_NVDLA_IS_pipe_1_reset = reset; // @[:@2141.4]
  assign NV_NVDLA_IS_pipe_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 60:25:@2142.4]
  assign NV_NVDLA_IS_pipe_1_io_ri = NV_NVDLA_IS_pipe_2_io_ro; // @[NV_NVDLA_DMAIF_rdrsp.scala 65:24:@2146.4]
  assign NV_NVDLA_IS_pipe_1_io_di = io_cvif_rd_rsp_pd_bits; // @[NV_NVDLA_DMAIF_rdrsp.scala 63:24:@2145.4]
  assign NV_NVDLA_IS_pipe_1_io_vi = io_cvif_rd_rsp_pd_valid; // @[NV_NVDLA_DMAIF_rdrsp.scala 61:24:@2143.4]
  assign NV_NVDLA_IS_pipe_2_reset = reset; // @[:@2159.4]
  assign NV_NVDLA_IS_pipe_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_DMAIF_rdrsp.scala 86:21:@2160.4]
  assign NV_NVDLA_IS_pipe_2_io_ri = io_dmaif_rd_rsp_pd_ready; // @[NV_NVDLA_DMAIF_rdrsp.scala 91:20:@2165.4]
  assign NV_NVDLA_IS_pipe_2_io_di = _T_48 | _T_53; // @[NV_NVDLA_DMAIF_rdrsp.scala 89:20:@2163.4]
  assign NV_NVDLA_IS_pipe_2_io_vi = NV_NVDLA_IS_pipe_io_vo | NV_NVDLA_IS_pipe_1_io_vo; // @[NV_NVDLA_DMAIF_rdrsp.scala 87:20:@2161.4]
endmodule
module nv_ram_rwsp( // @[:@2199.2]
  input          io_clk, // @[:@2202.4]
  input          io_re, // @[:@2202.4]
  input          io_we, // @[:@2202.4]
  input          io_ore, // @[:@2202.4]
  input  [2:0]   io_ra, // @[:@2202.4]
  input  [2:0]   io_wa, // @[:@2202.4]
  input  [256:0] io_di, // @[:@2202.4]
  output [256:0] io_dout // @[:@2202.4]
);
  reg [256:0] _T_26_0; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_0;
  reg [256:0] _T_26_1; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_1;
  reg [256:0] _T_26_2; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_2;
  reg [256:0] _T_26_3; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_3;
  reg [256:0] _T_26_4; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_4;
  reg [256:0] _T_26_5; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_5;
  reg [256:0] _T_26_6; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_6;
  reg [256:0] _T_26_7; // @[nv_ram_rwsp.scala 31:18:@2204.4]
  reg [287:0] _RAND_7;
  reg [2:0] _T_38; // @[nv_ram_rwsp.scala 32:19:@2205.4]
  reg [31:0] _RAND_8;
  reg [256:0] _T_40; // @[nv_ram_rwsp.scala 33:21:@2206.4]
  reg [287:0] _RAND_9;
  wire [256:0] _GEN_0; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_1; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_2; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_3; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_4; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_5; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_6; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_7; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  wire [256:0] _GEN_18; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_19; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_20; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_21; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_22; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_23; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  wire [256:0] _GEN_24; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_0 = 3'h0 == io_wa ? io_di : _T_26_0; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_1 = 3'h1 == io_wa ? io_di : _T_26_1; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_2 = 3'h2 == io_wa ? io_di : _T_26_2; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_3 = 3'h3 == io_wa ? io_di : _T_26_3; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_4 = 3'h4 == io_wa ? io_di : _T_26_4; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_5 = 3'h5 == io_wa ? io_di : _T_26_5; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_6 = 3'h6 == io_wa ? io_di : _T_26_6; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_7 = 3'h7 == io_wa ? io_di : _T_26_7; // @[nv_ram_rwsp.scala 36:20:@2208.6]
  assign _GEN_18 = 3'h1 == _T_38 ? _T_26_1 : _T_26_0; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_19 = 3'h2 == _T_38 ? _T_26_2 : _GEN_18; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_20 = 3'h3 == _T_38 ? _T_26_3 : _GEN_19; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_21 = 3'h4 == _T_38 ? _T_26_4 : _GEN_20; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_22 = 3'h5 == _T_38 ? _T_26_5 : _GEN_21; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_23 = 3'h6 == _T_38 ? _T_26_6 : _GEN_22; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign _GEN_24 = 3'h7 == _T_38 ? _T_26_7 : _GEN_23; // @[nv_ram_rwsp.scala 43:16:@2214.6]
  assign io_dout = _T_40; // @[nv_ram_rwsp.scala 45:13:@2216.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {9{`RANDOM}};
  _T_26_0 = _RAND_0[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {9{`RANDOM}};
  _T_26_1 = _RAND_1[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {9{`RANDOM}};
  _T_26_2 = _RAND_2[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {9{`RANDOM}};
  _T_26_3 = _RAND_3[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {9{`RANDOM}};
  _T_26_4 = _RAND_4[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {9{`RANDOM}};
  _T_26_5 = _RAND_5[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {9{`RANDOM}};
  _T_26_6 = _RAND_6[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {9{`RANDOM}};
  _T_26_7 = _RAND_7[256:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_38 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {9{`RANDOM}};
  _T_40 = _RAND_9[256:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (3'h0 == io_wa) begin
        _T_26_0 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h1 == io_wa) begin
        _T_26_1 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h2 == io_wa) begin
        _T_26_2 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h3 == io_wa) begin
        _T_26_3 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h4 == io_wa) begin
        _T_26_4 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h5 == io_wa) begin
        _T_26_5 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h6 == io_wa) begin
        _T_26_6 <= io_di;
      end
    end
    if (io_we) begin
      if (3'h7 == io_wa) begin
        _T_26_7 <= io_di;
      end
    end
    if (io_re) begin
      _T_38 <= io_ra;
    end
    if (io_ore) begin
      if (3'h7 == _T_38) begin
        _T_40 <= _T_26_7;
      end else begin
        if (3'h6 == _T_38) begin
          _T_40 <= _T_26_6;
        end else begin
          if (3'h5 == _T_38) begin
            _T_40 <= _T_26_5;
          end else begin
            if (3'h4 == _T_38) begin
              _T_40 <= _T_26_4;
            end else begin
              if (3'h3 == _T_38) begin
                _T_40 <= _T_26_3;
              end else begin
                if (3'h2 == _T_38) begin
                  _T_40 <= _T_26_2;
                end else begin
                  if (3'h1 == _T_38) begin
                    _T_40 <= _T_26_1;
                  end else begin
                    _T_40 <= _T_26_0;
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_fifo( // @[:@2218.2]
  input          clock, // @[:@2219.4]
  input          reset, // @[:@2220.4]
  input          io_clk, // @[:@2221.4]
  input          io_wr_pvld, // @[:@2221.4]
  output         io_wr_prdy, // @[:@2221.4]
  input  [256:0] io_wr_pd, // @[:@2221.4]
  output         io_rd_pvld, // @[:@2221.4]
  input          io_rd_prdy, // @[:@2221.4]
  output [256:0] io_rd_pd // @[:@2221.4]
);
  wire  nv_ram_rwsp_io_clk; // @[FIFO.scala 270:29:@2275.4]
  wire  nv_ram_rwsp_io_re; // @[FIFO.scala 270:29:@2275.4]
  wire  nv_ram_rwsp_io_we; // @[FIFO.scala 270:29:@2275.4]
  wire  nv_ram_rwsp_io_ore; // @[FIFO.scala 270:29:@2275.4]
  wire [2:0] nv_ram_rwsp_io_ra; // @[FIFO.scala 270:29:@2275.4]
  wire [2:0] nv_ram_rwsp_io_wa; // @[FIFO.scala 270:29:@2275.4]
  wire [256:0] nv_ram_rwsp_io_di; // @[FIFO.scala 270:29:@2275.4]
  wire [256:0] nv_ram_rwsp_io_dout; // @[FIFO.scala 270:29:@2275.4]
  reg  _T_26; // @[FIFO.scala 156:56:@2230.4]
  reg [31:0] _RAND_0;
  wire  _T_30; // @[FIFO.scala 182:23:@2232.4]
  wire  _T_33; // @[FIFO.scala 183:36:@2235.4]
  reg [3:0] _T_38; // @[FIFO.scala 186:53:@2238.4]
  reg [31:0] _RAND_1;
  wire [4:0] _T_40; // @[FIFO.scala 190:76:@2239.4]
  wire [4:0] _T_41; // @[FIFO.scala 190:76:@2240.4]
  wire [3:0] _T_42; // @[FIFO.scala 190:76:@2241.4]
  wire [3:0] _T_43; // @[FIFO.scala 190:43:@2242.4]
  wire [4:0] _T_45; // @[FIFO.scala 191:69:@2243.4]
  wire [3:0] _T_46; // @[FIFO.scala 191:69:@2244.4]
  wire [3:0] _T_47; // @[FIFO.scala 191:46:@2245.4]
  wire  _T_103; // @[FIFO.scala 331:38:@2306.4]
  wire [3:0] _T_48; // @[FIFO.scala 192:32:@2246.4]
  wire  _T_50; // @[FIFO.scala 194:80:@2247.4]
  wire  _T_52; // @[FIFO.scala 195:40:@2248.4]
  wire  _T_60; // @[FIFO.scala 202:27:@2256.4]
  wire [3:0] _GEN_0; // @[FIFO.scala 202:40:@2257.4]
  reg [2:0] _T_63; // @[FIFO.scala 215:68:@2260.4]
  reg [31:0] _RAND_2;
  wire [3:0] _T_65; // @[FIFO.scala 217:42:@2261.4]
  wire [2:0] _T_66; // @[FIFO.scala 217:42:@2262.4]
  wire [2:0] _GEN_1; // @[FIFO.scala 218:29:@2263.4]
  reg [2:0] _T_71; // @[FIFO.scala 224:63:@2267.4]
  reg [31:0] _RAND_3;
  wire [3:0] _T_73; // @[FIFO.scala 225:42:@2268.4]
  wire [2:0] _T_74; // @[FIFO.scala 225:42:@2269.4]
  wire [2:0] _GEN_2; // @[FIFO.scala 227:29:@2270.4]
  reg  _T_82; // @[FIFO.scala 289:73:@2289.4]
  reg [31:0] _RAND_4;
  reg  _T_85; // @[FIFO.scala 295:72:@2291.4]
  reg [31:0] _RAND_5;
  reg  _T_88; // @[FIFO.scala 297:97:@2292.4]
  reg [31:0] _RAND_6;
  reg [3:0] _T_91; // @[FIFO.scala 299:53:@2293.4]
  reg [31:0] _RAND_7;
  wire [4:0] _T_93; // @[FIFO.scala 300:74:@2294.4]
  wire [4:0] _T_94; // @[FIFO.scala 300:74:@2295.4]
  wire [3:0] _T_95; // @[FIFO.scala 300:74:@2296.4]
  wire [3:0] _T_96; // @[FIFO.scala 300:43:@2297.4]
  wire [4:0] _T_98; // @[FIFO.scala 301:68:@2298.4]
  wire [3:0] _T_99; // @[FIFO.scala 301:68:@2299.4]
  wire [3:0] _T_100; // @[FIFO.scala 301:46:@2300.4]
  wire [3:0] _T_101; // @[FIFO.scala 302:32:@2301.4]
  wire  _T_102; // @[FIFO.scala 303:25:@2302.4]
  wire [3:0] _GEN_3; // @[FIFO.scala 303:39:@2303.4]
  wire  _T_105; // @[FIFO.scala 333:77:@2308.4]
  wire  _T_107; // @[FIFO.scala 334:83:@2309.4]
  wire  _T_108; // @[FIFO.scala 335:44:@2310.4]
  wire  _T_109; // @[FIFO.scala 336:60:@2311.4]
  wire  _T_111; // @[FIFO.scala 336:81:@2313.4]
  wire  _GEN_4; // @[FIFO.scala 338:43:@2317.4]
  wire  _T_115; // @[FIFO.scala 341:66:@2320.4]
  wire  _T_116; // @[FIFO.scala 341:63:@2321.4]
  wire  _T_117; // @[FIFO.scala 341:43:@2322.4]
  nv_ram_rwsp nv_ram_rwsp ( // @[FIFO.scala 270:29:@2275.4]
    .io_clk(nv_ram_rwsp_io_clk),
    .io_re(nv_ram_rwsp_io_re),
    .io_we(nv_ram_rwsp_io_we),
    .io_ore(nv_ram_rwsp_io_ore),
    .io_ra(nv_ram_rwsp_io_ra),
    .io_wa(nv_ram_rwsp_io_wa),
    .io_di(nv_ram_rwsp_io_di),
    .io_dout(nv_ram_rwsp_io_dout)
  );
  assign _T_30 = _T_26 == 1'h0; // @[FIFO.scala 182:23:@2232.4]
  assign _T_33 = io_wr_pvld & _T_30; // @[FIFO.scala 183:36:@2235.4]
  assign _T_40 = _T_38 - 4'h1; // @[FIFO.scala 190:76:@2239.4]
  assign _T_41 = $unsigned(_T_40); // @[FIFO.scala 190:76:@2240.4]
  assign _T_42 = _T_41[3:0]; // @[FIFO.scala 190:76:@2241.4]
  assign _T_43 = _T_33 ? _T_38 : _T_42; // @[FIFO.scala 190:43:@2242.4]
  assign _T_45 = _T_38 + 4'h1; // @[FIFO.scala 191:69:@2243.4]
  assign _T_46 = _T_38 + 4'h1; // @[FIFO.scala 191:69:@2244.4]
  assign _T_47 = _T_33 ? _T_46 : _T_38; // @[FIFO.scala 191:46:@2245.4]
  assign _T_103 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 331:38:@2306.4]
  assign _T_48 = _T_103 ? _T_43 : _T_47; // @[FIFO.scala 192:32:@2246.4]
  assign _T_50 = _T_47 == 4'h8; // @[FIFO.scala 194:80:@2247.4]
  assign _T_52 = _T_103 ? 1'h0 : _T_50; // @[FIFO.scala 195:40:@2248.4]
  assign _T_60 = _T_33 ^ _T_103; // @[FIFO.scala 202:27:@2256.4]
  assign _GEN_0 = _T_60 ? _T_48 : _T_38; // @[FIFO.scala 202:40:@2257.4]
  assign _T_65 = _T_63 + 3'h1; // @[FIFO.scala 217:42:@2261.4]
  assign _T_66 = _T_63 + 3'h1; // @[FIFO.scala 217:42:@2262.4]
  assign _GEN_1 = _T_33 ? _T_66 : _T_63; // @[FIFO.scala 218:29:@2263.4]
  assign _T_73 = _T_71 + 3'h1; // @[FIFO.scala 225:42:@2268.4]
  assign _T_74 = _T_71 + 3'h1; // @[FIFO.scala 225:42:@2269.4]
  assign _GEN_2 = _T_103 ? _T_74 : _T_71; // @[FIFO.scala 227:29:@2270.4]
  assign _T_93 = _T_91 - 4'h1; // @[FIFO.scala 300:74:@2294.4]
  assign _T_94 = $unsigned(_T_93); // @[FIFO.scala 300:74:@2295.4]
  assign _T_95 = _T_94[3:0]; // @[FIFO.scala 300:74:@2296.4]
  assign _T_96 = _T_82 ? _T_91 : _T_95; // @[FIFO.scala 300:43:@2297.4]
  assign _T_98 = _T_91 + 4'h1; // @[FIFO.scala 301:68:@2298.4]
  assign _T_99 = _T_91 + 4'h1; // @[FIFO.scala 301:68:@2299.4]
  assign _T_100 = _T_82 ? _T_99 : _T_91; // @[FIFO.scala 301:46:@2300.4]
  assign _T_101 = _T_103 ? _T_96 : _T_100; // @[FIFO.scala 302:32:@2301.4]
  assign _T_102 = _T_82 | _T_103; // @[FIFO.scala 303:25:@2302.4]
  assign _GEN_3 = _T_102 ? _T_101 : _T_91; // @[FIFO.scala 303:39:@2303.4]
  assign _T_105 = _T_96 != 4'h0; // @[FIFO.scala 333:77:@2308.4]
  assign _T_107 = _T_100 != 4'h0; // @[FIFO.scala 334:83:@2309.4]
  assign _T_108 = _T_103 ? _T_105 : _T_107; // @[FIFO.scala 335:44:@2310.4]
  assign _T_109 = ~ _T_85; // @[FIFO.scala 336:60:@2311.4]
  assign _T_111 = _T_109 | _T_103; // @[FIFO.scala 336:81:@2313.4]
  assign _GEN_4 = _T_102 ? _T_108 : _T_85; // @[FIFO.scala 338:43:@2317.4]
  assign _T_115 = io_rd_prdy == 1'h0; // @[FIFO.scala 341:66:@2320.4]
  assign _T_116 = _T_88 & _T_115; // @[FIFO.scala 341:63:@2321.4]
  assign _T_117 = _T_85 | _T_116; // @[FIFO.scala 341:43:@2322.4]
  assign io_wr_prdy = _T_26 == 1'h0; // @[FIFO.scala 182:20:@2233.4]
  assign io_rd_pvld = _T_88; // @[FIFO.scala 344:24:@2324.4]
  assign io_rd_pd = nv_ram_rwsp_io_dout; // @[FIFO.scala 345:22:@2325.4]
  assign nv_ram_rwsp_io_clk = io_clk; // @[FIFO.scala 271:24:@2278.4]
  assign nv_ram_rwsp_io_re = _T_108 & _T_111; // @[FIFO.scala 279:23:@2285.4]
  assign nv_ram_rwsp_io_we = io_wr_pvld & _T_30; // @[FIFO.scala 276:23:@2281.4]
  assign nv_ram_rwsp_io_ore = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 280:24:@2286.4]
  assign nv_ram_rwsp_io_ra = _T_103 ? _T_74 : _T_71; // @[FIFO.scala 278:23:@2284.4]
  assign nv_ram_rwsp_io_wa = _T_63; // @[FIFO.scala 274:27:@2280.4]
  assign nv_ram_rwsp_io_di = io_wr_pd; // @[FIFO.scala 277:23:@2282.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_38 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_63 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_71 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_82 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_85 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_88 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_91 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_103) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_50;
      end
    end
    if (reset) begin
      _T_38 <= 4'h0;
    end else begin
      if (_T_60) begin
        if (_T_103) begin
          if (!(_T_33)) begin
            _T_38 <= _T_42;
          end
        end else begin
          if (_T_33) begin
            _T_38 <= _T_46;
          end
        end
      end
    end
    if (reset) begin
      _T_63 <= 3'h0;
    end else begin
      if (_T_33) begin
        _T_63 <= _T_66;
      end
    end
    if (reset) begin
      _T_71 <= 3'h0;
    end else begin
      if (_T_103) begin
        _T_71 <= _T_74;
      end
    end
    if (reset) begin
      _T_82 <= 1'h0;
    end else begin
      _T_82 <= _T_33;
    end
    if (reset) begin
      _T_85 <= 1'h0;
    end else begin
      if (_T_102) begin
        if (_T_103) begin
          _T_85 <= _T_105;
        end else begin
          _T_85 <= _T_107;
        end
      end
    end
    if (reset) begin
      _T_88 <= 1'h0;
    end else begin
      _T_88 <= _T_117;
    end
    if (reset) begin
      _T_91 <= 4'h0;
    end else begin
      if (_T_102) begin
        if (_T_103) begin
          if (!(_T_82)) begin
            _T_91 <= _T_95;
          end
        end else begin
          if (_T_82) begin
            _T_91 <= _T_99;
          end
        end
      end
    end
  end
endmodule
module nv_ram_rwsp_1( // @[:@2372.2]
  input        io_clk, // @[:@2375.4]
  input        io_re, // @[:@2375.4]
  input        io_we, // @[:@2375.4]
  input        io_ore, // @[:@2375.4]
  input  [6:0] io_ra, // @[:@2375.4]
  input  [6:0] io_wa, // @[:@2375.4]
  input  [5:0] io_di, // @[:@2375.4]
  output [5:0] io_dout // @[:@2375.4]
);
  reg [5:0] _T_26_0; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_26_1; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_1;
  reg [5:0] _T_26_2; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_2;
  reg [5:0] _T_26_3; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_3;
  reg [5:0] _T_26_4; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_4;
  reg [5:0] _T_26_5; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_5;
  reg [5:0] _T_26_6; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_6;
  reg [5:0] _T_26_7; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_7;
  reg [5:0] _T_26_8; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_8;
  reg [5:0] _T_26_9; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_9;
  reg [5:0] _T_26_10; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_10;
  reg [5:0] _T_26_11; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_26_12; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_12;
  reg [5:0] _T_26_13; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_13;
  reg [5:0] _T_26_14; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_14;
  reg [5:0] _T_26_15; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_15;
  reg [5:0] _T_26_16; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_16;
  reg [5:0] _T_26_17; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_17;
  reg [5:0] _T_26_18; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_18;
  reg [5:0] _T_26_19; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_19;
  reg [5:0] _T_26_20; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_20;
  reg [5:0] _T_26_21; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_21;
  reg [5:0] _T_26_22; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_22;
  reg [5:0] _T_26_23; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_23;
  reg [5:0] _T_26_24; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_24;
  reg [5:0] _T_26_25; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_25;
  reg [5:0] _T_26_26; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_26;
  reg [5:0] _T_26_27; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_27;
  reg [5:0] _T_26_28; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_28;
  reg [5:0] _T_26_29; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_29;
  reg [5:0] _T_26_30; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_30;
  reg [5:0] _T_26_31; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_31;
  reg [5:0] _T_26_32; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_32;
  reg [5:0] _T_26_33; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_33;
  reg [5:0] _T_26_34; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_34;
  reg [5:0] _T_26_35; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_26_36; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_26_37; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_37;
  reg [5:0] _T_26_38; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_38;
  reg [5:0] _T_26_39; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_39;
  reg [5:0] _T_26_40; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_40;
  reg [5:0] _T_26_41; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_41;
  reg [5:0] _T_26_42; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_42;
  reg [5:0] _T_26_43; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_43;
  reg [5:0] _T_26_44; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_44;
  reg [5:0] _T_26_45; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_45;
  reg [5:0] _T_26_46; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_46;
  reg [5:0] _T_26_47; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_47;
  reg [5:0] _T_26_48; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_48;
  reg [5:0] _T_26_49; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_49;
  reg [5:0] _T_26_50; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_50;
  reg [5:0] _T_26_51; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_51;
  reg [5:0] _T_26_52; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_52;
  reg [5:0] _T_26_53; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_53;
  reg [5:0] _T_26_54; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_54;
  reg [5:0] _T_26_55; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_55;
  reg [5:0] _T_26_56; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_56;
  reg [5:0] _T_26_57; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_57;
  reg [5:0] _T_26_58; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_58;
  reg [5:0] _T_26_59; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_59;
  reg [5:0] _T_26_60; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_60;
  reg [5:0] _T_26_61; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_61;
  reg [5:0] _T_26_62; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_62;
  reg [5:0] _T_26_63; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_63;
  reg [5:0] _T_26_64; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_64;
  reg [5:0] _T_26_65; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_65;
  reg [5:0] _T_26_66; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_66;
  reg [5:0] _T_26_67; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_67;
  reg [5:0] _T_26_68; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_68;
  reg [5:0] _T_26_69; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_69;
  reg [5:0] _T_26_70; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_70;
  reg [5:0] _T_26_71; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_71;
  reg [5:0] _T_26_72; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_72;
  reg [5:0] _T_26_73; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_73;
  reg [5:0] _T_26_74; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_74;
  reg [5:0] _T_26_75; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_75;
  reg [5:0] _T_26_76; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_76;
  reg [5:0] _T_26_77; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_77;
  reg [5:0] _T_26_78; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_78;
  reg [5:0] _T_26_79; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_79;
  reg [5:0] _T_26_80; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_80;
  reg [5:0] _T_26_81; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_81;
  reg [5:0] _T_26_82; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_82;
  reg [5:0] _T_26_83; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_83;
  reg [5:0] _T_26_84; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_84;
  reg [5:0] _T_26_85; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_85;
  reg [5:0] _T_26_86; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_86;
  reg [5:0] _T_26_87; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_87;
  reg [5:0] _T_26_88; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_88;
  reg [5:0] _T_26_89; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_89;
  reg [5:0] _T_26_90; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_90;
  reg [5:0] _T_26_91; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_91;
  reg [5:0] _T_26_92; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_92;
  reg [5:0] _T_26_93; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_93;
  reg [5:0] _T_26_94; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_94;
  reg [5:0] _T_26_95; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_95;
  reg [5:0] _T_26_96; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_96;
  reg [5:0] _T_26_97; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_97;
  reg [5:0] _T_26_98; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_98;
  reg [5:0] _T_26_99; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_99;
  reg [5:0] _T_26_100; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_100;
  reg [5:0] _T_26_101; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_101;
  reg [5:0] _T_26_102; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_102;
  reg [5:0] _T_26_103; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_103;
  reg [5:0] _T_26_104; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_104;
  reg [5:0] _T_26_105; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_105;
  reg [5:0] _T_26_106; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_106;
  reg [5:0] _T_26_107; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_107;
  reg [5:0] _T_26_108; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_108;
  reg [5:0] _T_26_109; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_109;
  reg [5:0] _T_26_110; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_110;
  reg [5:0] _T_26_111; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_111;
  reg [5:0] _T_26_112; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_112;
  reg [5:0] _T_26_113; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_113;
  reg [5:0] _T_26_114; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_114;
  reg [5:0] _T_26_115; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_115;
  reg [5:0] _T_26_116; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_116;
  reg [5:0] _T_26_117; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_117;
  reg [5:0] _T_26_118; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_118;
  reg [5:0] _T_26_119; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_119;
  reg [5:0] _T_26_120; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_120;
  reg [5:0] _T_26_121; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_121;
  reg [5:0] _T_26_122; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_122;
  reg [5:0] _T_26_123; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_123;
  reg [5:0] _T_26_124; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_124;
  reg [5:0] _T_26_125; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_125;
  reg [5:0] _T_26_126; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_126;
  reg [5:0] _T_26_127; // @[nv_ram_rwsp.scala 31:18:@2377.4]
  reg [31:0] _RAND_127;
  reg [6:0] _T_158; // @[nv_ram_rwsp.scala 32:19:@2378.4]
  reg [31:0] _RAND_128;
  reg [5:0] _T_160; // @[nv_ram_rwsp.scala 33:21:@2379.4]
  reg [31:0] _RAND_129;
  wire [5:0] _GEN_0; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_1; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_2; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_3; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_4; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_5; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_6; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_7; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_8; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_9; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_10; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_11; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_12; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_13; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_14; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_15; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_16; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_17; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_18; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_19; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_20; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_21; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_22; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_23; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_24; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_25; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_26; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_27; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_28; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_29; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_30; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_31; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_32; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_33; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_34; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_35; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_36; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_37; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_38; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_39; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_40; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_41; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_42; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_43; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_44; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_45; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_46; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_47; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_48; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_49; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_50; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_51; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_52; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_53; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_54; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_55; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_56; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_57; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_58; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_59; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_60; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_61; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_62; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_63; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_64; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_65; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_66; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_67; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_68; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_69; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_70; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_71; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_72; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_73; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_74; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_75; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_76; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_77; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_78; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_79; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_80; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_81; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_82; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_83; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_84; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_85; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_86; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_87; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_88; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_89; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_90; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_91; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_92; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_93; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_94; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_95; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_96; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_97; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_98; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_99; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_100; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_101; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_102; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_103; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_104; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_105; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_106; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_107; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_108; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_109; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_110; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_111; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_112; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_113; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_114; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_115; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_116; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_117; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_118; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_119; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_120; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_121; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_122; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_123; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_124; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_125; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_126; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_127; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  wire [5:0] _GEN_258; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_259; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_260; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_261; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_262; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_263; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_264; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_265; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_266; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_267; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_268; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_269; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_270; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_271; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_272; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_273; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_274; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_275; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_276; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_277; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_278; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_279; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_280; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_281; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_282; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_283; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_284; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_285; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_286; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_287; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_288; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_289; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_290; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_291; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_292; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_293; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_294; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_295; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_296; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_297; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_298; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_299; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_300; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_301; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_302; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_303; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_304; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_305; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_306; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_307; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_308; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_309; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_310; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_311; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_312; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_313; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_314; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_315; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_316; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_317; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_318; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_319; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_320; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_321; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_322; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_323; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_324; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_325; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_326; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_327; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_328; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_329; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_330; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_331; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_332; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_333; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_334; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_335; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_336; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_337; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_338; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_339; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_340; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_341; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_342; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_343; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_344; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_345; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_346; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_347; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_348; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_349; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_350; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_351; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_352; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_353; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_354; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_355; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_356; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_357; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_358; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_359; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_360; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_361; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_362; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_363; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_364; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_365; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_366; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_367; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_368; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_369; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_370; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_371; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_372; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_373; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_374; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_375; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_376; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_377; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_378; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_379; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_380; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_381; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_382; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_383; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  wire [5:0] _GEN_384; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_0 = 7'h0 == io_wa ? io_di : _T_26_0; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_1 = 7'h1 == io_wa ? io_di : _T_26_1; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_2 = 7'h2 == io_wa ? io_di : _T_26_2; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_3 = 7'h3 == io_wa ? io_di : _T_26_3; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_4 = 7'h4 == io_wa ? io_di : _T_26_4; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_5 = 7'h5 == io_wa ? io_di : _T_26_5; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_6 = 7'h6 == io_wa ? io_di : _T_26_6; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_7 = 7'h7 == io_wa ? io_di : _T_26_7; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_8 = 7'h8 == io_wa ? io_di : _T_26_8; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_9 = 7'h9 == io_wa ? io_di : _T_26_9; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_10 = 7'ha == io_wa ? io_di : _T_26_10; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_11 = 7'hb == io_wa ? io_di : _T_26_11; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_12 = 7'hc == io_wa ? io_di : _T_26_12; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_13 = 7'hd == io_wa ? io_di : _T_26_13; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_14 = 7'he == io_wa ? io_di : _T_26_14; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_15 = 7'hf == io_wa ? io_di : _T_26_15; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_16 = 7'h10 == io_wa ? io_di : _T_26_16; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_17 = 7'h11 == io_wa ? io_di : _T_26_17; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_18 = 7'h12 == io_wa ? io_di : _T_26_18; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_19 = 7'h13 == io_wa ? io_di : _T_26_19; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_20 = 7'h14 == io_wa ? io_di : _T_26_20; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_21 = 7'h15 == io_wa ? io_di : _T_26_21; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_22 = 7'h16 == io_wa ? io_di : _T_26_22; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_23 = 7'h17 == io_wa ? io_di : _T_26_23; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_24 = 7'h18 == io_wa ? io_di : _T_26_24; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_25 = 7'h19 == io_wa ? io_di : _T_26_25; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_26 = 7'h1a == io_wa ? io_di : _T_26_26; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_27 = 7'h1b == io_wa ? io_di : _T_26_27; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_28 = 7'h1c == io_wa ? io_di : _T_26_28; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_29 = 7'h1d == io_wa ? io_di : _T_26_29; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_30 = 7'h1e == io_wa ? io_di : _T_26_30; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_31 = 7'h1f == io_wa ? io_di : _T_26_31; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_32 = 7'h20 == io_wa ? io_di : _T_26_32; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_33 = 7'h21 == io_wa ? io_di : _T_26_33; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_34 = 7'h22 == io_wa ? io_di : _T_26_34; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_35 = 7'h23 == io_wa ? io_di : _T_26_35; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_36 = 7'h24 == io_wa ? io_di : _T_26_36; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_37 = 7'h25 == io_wa ? io_di : _T_26_37; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_38 = 7'h26 == io_wa ? io_di : _T_26_38; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_39 = 7'h27 == io_wa ? io_di : _T_26_39; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_40 = 7'h28 == io_wa ? io_di : _T_26_40; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_41 = 7'h29 == io_wa ? io_di : _T_26_41; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_42 = 7'h2a == io_wa ? io_di : _T_26_42; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_43 = 7'h2b == io_wa ? io_di : _T_26_43; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_44 = 7'h2c == io_wa ? io_di : _T_26_44; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_45 = 7'h2d == io_wa ? io_di : _T_26_45; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_46 = 7'h2e == io_wa ? io_di : _T_26_46; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_47 = 7'h2f == io_wa ? io_di : _T_26_47; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_48 = 7'h30 == io_wa ? io_di : _T_26_48; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_49 = 7'h31 == io_wa ? io_di : _T_26_49; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_50 = 7'h32 == io_wa ? io_di : _T_26_50; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_51 = 7'h33 == io_wa ? io_di : _T_26_51; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_52 = 7'h34 == io_wa ? io_di : _T_26_52; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_53 = 7'h35 == io_wa ? io_di : _T_26_53; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_54 = 7'h36 == io_wa ? io_di : _T_26_54; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_55 = 7'h37 == io_wa ? io_di : _T_26_55; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_56 = 7'h38 == io_wa ? io_di : _T_26_56; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_57 = 7'h39 == io_wa ? io_di : _T_26_57; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_58 = 7'h3a == io_wa ? io_di : _T_26_58; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_59 = 7'h3b == io_wa ? io_di : _T_26_59; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_60 = 7'h3c == io_wa ? io_di : _T_26_60; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_61 = 7'h3d == io_wa ? io_di : _T_26_61; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_62 = 7'h3e == io_wa ? io_di : _T_26_62; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_63 = 7'h3f == io_wa ? io_di : _T_26_63; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_64 = 7'h40 == io_wa ? io_di : _T_26_64; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_65 = 7'h41 == io_wa ? io_di : _T_26_65; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_66 = 7'h42 == io_wa ? io_di : _T_26_66; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_67 = 7'h43 == io_wa ? io_di : _T_26_67; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_68 = 7'h44 == io_wa ? io_di : _T_26_68; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_69 = 7'h45 == io_wa ? io_di : _T_26_69; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_70 = 7'h46 == io_wa ? io_di : _T_26_70; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_71 = 7'h47 == io_wa ? io_di : _T_26_71; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_72 = 7'h48 == io_wa ? io_di : _T_26_72; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_73 = 7'h49 == io_wa ? io_di : _T_26_73; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_74 = 7'h4a == io_wa ? io_di : _T_26_74; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_75 = 7'h4b == io_wa ? io_di : _T_26_75; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_76 = 7'h4c == io_wa ? io_di : _T_26_76; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_77 = 7'h4d == io_wa ? io_di : _T_26_77; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_78 = 7'h4e == io_wa ? io_di : _T_26_78; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_79 = 7'h4f == io_wa ? io_di : _T_26_79; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_80 = 7'h50 == io_wa ? io_di : _T_26_80; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_81 = 7'h51 == io_wa ? io_di : _T_26_81; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_82 = 7'h52 == io_wa ? io_di : _T_26_82; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_83 = 7'h53 == io_wa ? io_di : _T_26_83; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_84 = 7'h54 == io_wa ? io_di : _T_26_84; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_85 = 7'h55 == io_wa ? io_di : _T_26_85; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_86 = 7'h56 == io_wa ? io_di : _T_26_86; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_87 = 7'h57 == io_wa ? io_di : _T_26_87; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_88 = 7'h58 == io_wa ? io_di : _T_26_88; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_89 = 7'h59 == io_wa ? io_di : _T_26_89; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_90 = 7'h5a == io_wa ? io_di : _T_26_90; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_91 = 7'h5b == io_wa ? io_di : _T_26_91; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_92 = 7'h5c == io_wa ? io_di : _T_26_92; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_93 = 7'h5d == io_wa ? io_di : _T_26_93; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_94 = 7'h5e == io_wa ? io_di : _T_26_94; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_95 = 7'h5f == io_wa ? io_di : _T_26_95; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_96 = 7'h60 == io_wa ? io_di : _T_26_96; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_97 = 7'h61 == io_wa ? io_di : _T_26_97; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_98 = 7'h62 == io_wa ? io_di : _T_26_98; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_99 = 7'h63 == io_wa ? io_di : _T_26_99; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_100 = 7'h64 == io_wa ? io_di : _T_26_100; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_101 = 7'h65 == io_wa ? io_di : _T_26_101; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_102 = 7'h66 == io_wa ? io_di : _T_26_102; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_103 = 7'h67 == io_wa ? io_di : _T_26_103; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_104 = 7'h68 == io_wa ? io_di : _T_26_104; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_105 = 7'h69 == io_wa ? io_di : _T_26_105; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_106 = 7'h6a == io_wa ? io_di : _T_26_106; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_107 = 7'h6b == io_wa ? io_di : _T_26_107; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_108 = 7'h6c == io_wa ? io_di : _T_26_108; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_109 = 7'h6d == io_wa ? io_di : _T_26_109; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_110 = 7'h6e == io_wa ? io_di : _T_26_110; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_111 = 7'h6f == io_wa ? io_di : _T_26_111; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_112 = 7'h70 == io_wa ? io_di : _T_26_112; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_113 = 7'h71 == io_wa ? io_di : _T_26_113; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_114 = 7'h72 == io_wa ? io_di : _T_26_114; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_115 = 7'h73 == io_wa ? io_di : _T_26_115; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_116 = 7'h74 == io_wa ? io_di : _T_26_116; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_117 = 7'h75 == io_wa ? io_di : _T_26_117; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_118 = 7'h76 == io_wa ? io_di : _T_26_118; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_119 = 7'h77 == io_wa ? io_di : _T_26_119; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_120 = 7'h78 == io_wa ? io_di : _T_26_120; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_121 = 7'h79 == io_wa ? io_di : _T_26_121; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_122 = 7'h7a == io_wa ? io_di : _T_26_122; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_123 = 7'h7b == io_wa ? io_di : _T_26_123; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_124 = 7'h7c == io_wa ? io_di : _T_26_124; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_125 = 7'h7d == io_wa ? io_di : _T_26_125; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_126 = 7'h7e == io_wa ? io_di : _T_26_126; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_127 = 7'h7f == io_wa ? io_di : _T_26_127; // @[nv_ram_rwsp.scala 36:20:@2381.6]
  assign _GEN_258 = 7'h1 == _T_158 ? _T_26_1 : _T_26_0; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_259 = 7'h2 == _T_158 ? _T_26_2 : _GEN_258; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_260 = 7'h3 == _T_158 ? _T_26_3 : _GEN_259; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_261 = 7'h4 == _T_158 ? _T_26_4 : _GEN_260; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_262 = 7'h5 == _T_158 ? _T_26_5 : _GEN_261; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_263 = 7'h6 == _T_158 ? _T_26_6 : _GEN_262; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_264 = 7'h7 == _T_158 ? _T_26_7 : _GEN_263; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_265 = 7'h8 == _T_158 ? _T_26_8 : _GEN_264; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_266 = 7'h9 == _T_158 ? _T_26_9 : _GEN_265; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_267 = 7'ha == _T_158 ? _T_26_10 : _GEN_266; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_268 = 7'hb == _T_158 ? _T_26_11 : _GEN_267; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_269 = 7'hc == _T_158 ? _T_26_12 : _GEN_268; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_270 = 7'hd == _T_158 ? _T_26_13 : _GEN_269; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_271 = 7'he == _T_158 ? _T_26_14 : _GEN_270; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_272 = 7'hf == _T_158 ? _T_26_15 : _GEN_271; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_273 = 7'h10 == _T_158 ? _T_26_16 : _GEN_272; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_274 = 7'h11 == _T_158 ? _T_26_17 : _GEN_273; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_275 = 7'h12 == _T_158 ? _T_26_18 : _GEN_274; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_276 = 7'h13 == _T_158 ? _T_26_19 : _GEN_275; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_277 = 7'h14 == _T_158 ? _T_26_20 : _GEN_276; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_278 = 7'h15 == _T_158 ? _T_26_21 : _GEN_277; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_279 = 7'h16 == _T_158 ? _T_26_22 : _GEN_278; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_280 = 7'h17 == _T_158 ? _T_26_23 : _GEN_279; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_281 = 7'h18 == _T_158 ? _T_26_24 : _GEN_280; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_282 = 7'h19 == _T_158 ? _T_26_25 : _GEN_281; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_283 = 7'h1a == _T_158 ? _T_26_26 : _GEN_282; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_284 = 7'h1b == _T_158 ? _T_26_27 : _GEN_283; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_285 = 7'h1c == _T_158 ? _T_26_28 : _GEN_284; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_286 = 7'h1d == _T_158 ? _T_26_29 : _GEN_285; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_287 = 7'h1e == _T_158 ? _T_26_30 : _GEN_286; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_288 = 7'h1f == _T_158 ? _T_26_31 : _GEN_287; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_289 = 7'h20 == _T_158 ? _T_26_32 : _GEN_288; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_290 = 7'h21 == _T_158 ? _T_26_33 : _GEN_289; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_291 = 7'h22 == _T_158 ? _T_26_34 : _GEN_290; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_292 = 7'h23 == _T_158 ? _T_26_35 : _GEN_291; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_293 = 7'h24 == _T_158 ? _T_26_36 : _GEN_292; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_294 = 7'h25 == _T_158 ? _T_26_37 : _GEN_293; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_295 = 7'h26 == _T_158 ? _T_26_38 : _GEN_294; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_296 = 7'h27 == _T_158 ? _T_26_39 : _GEN_295; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_297 = 7'h28 == _T_158 ? _T_26_40 : _GEN_296; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_298 = 7'h29 == _T_158 ? _T_26_41 : _GEN_297; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_299 = 7'h2a == _T_158 ? _T_26_42 : _GEN_298; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_300 = 7'h2b == _T_158 ? _T_26_43 : _GEN_299; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_301 = 7'h2c == _T_158 ? _T_26_44 : _GEN_300; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_302 = 7'h2d == _T_158 ? _T_26_45 : _GEN_301; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_303 = 7'h2e == _T_158 ? _T_26_46 : _GEN_302; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_304 = 7'h2f == _T_158 ? _T_26_47 : _GEN_303; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_305 = 7'h30 == _T_158 ? _T_26_48 : _GEN_304; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_306 = 7'h31 == _T_158 ? _T_26_49 : _GEN_305; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_307 = 7'h32 == _T_158 ? _T_26_50 : _GEN_306; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_308 = 7'h33 == _T_158 ? _T_26_51 : _GEN_307; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_309 = 7'h34 == _T_158 ? _T_26_52 : _GEN_308; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_310 = 7'h35 == _T_158 ? _T_26_53 : _GEN_309; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_311 = 7'h36 == _T_158 ? _T_26_54 : _GEN_310; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_312 = 7'h37 == _T_158 ? _T_26_55 : _GEN_311; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_313 = 7'h38 == _T_158 ? _T_26_56 : _GEN_312; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_314 = 7'h39 == _T_158 ? _T_26_57 : _GEN_313; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_315 = 7'h3a == _T_158 ? _T_26_58 : _GEN_314; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_316 = 7'h3b == _T_158 ? _T_26_59 : _GEN_315; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_317 = 7'h3c == _T_158 ? _T_26_60 : _GEN_316; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_318 = 7'h3d == _T_158 ? _T_26_61 : _GEN_317; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_319 = 7'h3e == _T_158 ? _T_26_62 : _GEN_318; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_320 = 7'h3f == _T_158 ? _T_26_63 : _GEN_319; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_321 = 7'h40 == _T_158 ? _T_26_64 : _GEN_320; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_322 = 7'h41 == _T_158 ? _T_26_65 : _GEN_321; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_323 = 7'h42 == _T_158 ? _T_26_66 : _GEN_322; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_324 = 7'h43 == _T_158 ? _T_26_67 : _GEN_323; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_325 = 7'h44 == _T_158 ? _T_26_68 : _GEN_324; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_326 = 7'h45 == _T_158 ? _T_26_69 : _GEN_325; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_327 = 7'h46 == _T_158 ? _T_26_70 : _GEN_326; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_328 = 7'h47 == _T_158 ? _T_26_71 : _GEN_327; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_329 = 7'h48 == _T_158 ? _T_26_72 : _GEN_328; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_330 = 7'h49 == _T_158 ? _T_26_73 : _GEN_329; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_331 = 7'h4a == _T_158 ? _T_26_74 : _GEN_330; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_332 = 7'h4b == _T_158 ? _T_26_75 : _GEN_331; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_333 = 7'h4c == _T_158 ? _T_26_76 : _GEN_332; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_334 = 7'h4d == _T_158 ? _T_26_77 : _GEN_333; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_335 = 7'h4e == _T_158 ? _T_26_78 : _GEN_334; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_336 = 7'h4f == _T_158 ? _T_26_79 : _GEN_335; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_337 = 7'h50 == _T_158 ? _T_26_80 : _GEN_336; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_338 = 7'h51 == _T_158 ? _T_26_81 : _GEN_337; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_339 = 7'h52 == _T_158 ? _T_26_82 : _GEN_338; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_340 = 7'h53 == _T_158 ? _T_26_83 : _GEN_339; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_341 = 7'h54 == _T_158 ? _T_26_84 : _GEN_340; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_342 = 7'h55 == _T_158 ? _T_26_85 : _GEN_341; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_343 = 7'h56 == _T_158 ? _T_26_86 : _GEN_342; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_344 = 7'h57 == _T_158 ? _T_26_87 : _GEN_343; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_345 = 7'h58 == _T_158 ? _T_26_88 : _GEN_344; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_346 = 7'h59 == _T_158 ? _T_26_89 : _GEN_345; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_347 = 7'h5a == _T_158 ? _T_26_90 : _GEN_346; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_348 = 7'h5b == _T_158 ? _T_26_91 : _GEN_347; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_349 = 7'h5c == _T_158 ? _T_26_92 : _GEN_348; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_350 = 7'h5d == _T_158 ? _T_26_93 : _GEN_349; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_351 = 7'h5e == _T_158 ? _T_26_94 : _GEN_350; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_352 = 7'h5f == _T_158 ? _T_26_95 : _GEN_351; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_353 = 7'h60 == _T_158 ? _T_26_96 : _GEN_352; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_354 = 7'h61 == _T_158 ? _T_26_97 : _GEN_353; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_355 = 7'h62 == _T_158 ? _T_26_98 : _GEN_354; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_356 = 7'h63 == _T_158 ? _T_26_99 : _GEN_355; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_357 = 7'h64 == _T_158 ? _T_26_100 : _GEN_356; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_358 = 7'h65 == _T_158 ? _T_26_101 : _GEN_357; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_359 = 7'h66 == _T_158 ? _T_26_102 : _GEN_358; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_360 = 7'h67 == _T_158 ? _T_26_103 : _GEN_359; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_361 = 7'h68 == _T_158 ? _T_26_104 : _GEN_360; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_362 = 7'h69 == _T_158 ? _T_26_105 : _GEN_361; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_363 = 7'h6a == _T_158 ? _T_26_106 : _GEN_362; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_364 = 7'h6b == _T_158 ? _T_26_107 : _GEN_363; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_365 = 7'h6c == _T_158 ? _T_26_108 : _GEN_364; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_366 = 7'h6d == _T_158 ? _T_26_109 : _GEN_365; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_367 = 7'h6e == _T_158 ? _T_26_110 : _GEN_366; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_368 = 7'h6f == _T_158 ? _T_26_111 : _GEN_367; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_369 = 7'h70 == _T_158 ? _T_26_112 : _GEN_368; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_370 = 7'h71 == _T_158 ? _T_26_113 : _GEN_369; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_371 = 7'h72 == _T_158 ? _T_26_114 : _GEN_370; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_372 = 7'h73 == _T_158 ? _T_26_115 : _GEN_371; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_373 = 7'h74 == _T_158 ? _T_26_116 : _GEN_372; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_374 = 7'h75 == _T_158 ? _T_26_117 : _GEN_373; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_375 = 7'h76 == _T_158 ? _T_26_118 : _GEN_374; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_376 = 7'h77 == _T_158 ? _T_26_119 : _GEN_375; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_377 = 7'h78 == _T_158 ? _T_26_120 : _GEN_376; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_378 = 7'h79 == _T_158 ? _T_26_121 : _GEN_377; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_379 = 7'h7a == _T_158 ? _T_26_122 : _GEN_378; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_380 = 7'h7b == _T_158 ? _T_26_123 : _GEN_379; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_381 = 7'h7c == _T_158 ? _T_26_124 : _GEN_380; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_382 = 7'h7d == _T_158 ? _T_26_125 : _GEN_381; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_383 = 7'h7e == _T_158 ? _T_26_126 : _GEN_382; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign _GEN_384 = 7'h7f == _T_158 ? _T_26_127 : _GEN_383; // @[nv_ram_rwsp.scala 43:16:@2387.6]
  assign io_dout = _T_160; // @[nv_ram_rwsp.scala 45:13:@2389.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26_0 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26_1 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_26_2 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26_3 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_26_4 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_26_5 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_26_6 = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_26_7 = _RAND_7[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_26_8 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_26_9 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_26_10 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_26_11 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_26_12 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_26_13 = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_26_14 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_26_15 = _RAND_15[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_26_16 = _RAND_16[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_26_17 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_26_18 = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_26_19 = _RAND_19[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_26_20 = _RAND_20[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_26_21 = _RAND_21[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_26_22 = _RAND_22[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_26_23 = _RAND_23[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_26_24 = _RAND_24[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_26_25 = _RAND_25[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26_26 = _RAND_26[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_26_27 = _RAND_27[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_26_28 = _RAND_28[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_26_29 = _RAND_29[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_26_30 = _RAND_30[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_26_31 = _RAND_31[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_26_32 = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_26_33 = _RAND_33[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_26_34 = _RAND_34[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_26_35 = _RAND_35[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_26_36 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_26_37 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_26_38 = _RAND_38[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_26_39 = _RAND_39[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_26_40 = _RAND_40[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_26_41 = _RAND_41[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_26_42 = _RAND_42[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_26_43 = _RAND_43[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_26_44 = _RAND_44[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_26_45 = _RAND_45[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_26_46 = _RAND_46[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_26_47 = _RAND_47[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_26_48 = _RAND_48[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_26_49 = _RAND_49[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_26_50 = _RAND_50[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_26_51 = _RAND_51[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_26_52 = _RAND_52[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_26_53 = _RAND_53[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_26_54 = _RAND_54[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_26_55 = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_26_56 = _RAND_56[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_26_57 = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_26_58 = _RAND_58[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_26_59 = _RAND_59[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_26_60 = _RAND_60[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_26_61 = _RAND_61[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_26_62 = _RAND_62[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_26_63 = _RAND_63[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_26_64 = _RAND_64[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_26_65 = _RAND_65[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_26_66 = _RAND_66[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_26_67 = _RAND_67[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_26_68 = _RAND_68[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_26_69 = _RAND_69[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_26_70 = _RAND_70[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_26_71 = _RAND_71[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_26_72 = _RAND_72[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_26_73 = _RAND_73[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_26_74 = _RAND_74[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_26_75 = _RAND_75[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_26_76 = _RAND_76[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_26_77 = _RAND_77[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_26_78 = _RAND_78[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_26_79 = _RAND_79[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_26_80 = _RAND_80[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_26_81 = _RAND_81[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_26_82 = _RAND_82[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_26_83 = _RAND_83[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_26_84 = _RAND_84[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_26_85 = _RAND_85[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_26_86 = _RAND_86[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_26_87 = _RAND_87[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_26_88 = _RAND_88[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_26_89 = _RAND_89[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_26_90 = _RAND_90[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_26_91 = _RAND_91[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_26_92 = _RAND_92[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_26_93 = _RAND_93[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_26_94 = _RAND_94[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_26_95 = _RAND_95[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_26_96 = _RAND_96[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_26_97 = _RAND_97[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_26_98 = _RAND_98[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_26_99 = _RAND_99[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_26_100 = _RAND_100[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_26_101 = _RAND_101[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_26_102 = _RAND_102[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_26_103 = _RAND_103[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_26_104 = _RAND_104[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_26_105 = _RAND_105[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_26_106 = _RAND_106[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_26_107 = _RAND_107[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_26_108 = _RAND_108[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_26_109 = _RAND_109[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_26_110 = _RAND_110[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_26_111 = _RAND_111[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_26_112 = _RAND_112[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_26_113 = _RAND_113[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_26_114 = _RAND_114[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_26_115 = _RAND_115[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_26_116 = _RAND_116[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_26_117 = _RAND_117[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_26_118 = _RAND_118[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_26_119 = _RAND_119[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_26_120 = _RAND_120[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_26_121 = _RAND_121[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_26_122 = _RAND_122[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_26_123 = _RAND_123[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_26_124 = _RAND_124[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_26_125 = _RAND_125[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_26_126 = _RAND_126[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_26_127 = _RAND_127[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_158 = _RAND_128[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_160 = _RAND_129[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (7'h0 == io_wa) begin
        _T_26_0 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1 == io_wa) begin
        _T_26_1 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2 == io_wa) begin
        _T_26_2 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3 == io_wa) begin
        _T_26_3 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4 == io_wa) begin
        _T_26_4 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5 == io_wa) begin
        _T_26_5 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6 == io_wa) begin
        _T_26_6 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7 == io_wa) begin
        _T_26_7 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h8 == io_wa) begin
        _T_26_8 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h9 == io_wa) begin
        _T_26_9 <= io_di;
      end
    end
    if (io_we) begin
      if (7'ha == io_wa) begin
        _T_26_10 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hb == io_wa) begin
        _T_26_11 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hc == io_wa) begin
        _T_26_12 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hd == io_wa) begin
        _T_26_13 <= io_di;
      end
    end
    if (io_we) begin
      if (7'he == io_wa) begin
        _T_26_14 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hf == io_wa) begin
        _T_26_15 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h10 == io_wa) begin
        _T_26_16 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h11 == io_wa) begin
        _T_26_17 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h12 == io_wa) begin
        _T_26_18 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h13 == io_wa) begin
        _T_26_19 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h14 == io_wa) begin
        _T_26_20 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h15 == io_wa) begin
        _T_26_21 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h16 == io_wa) begin
        _T_26_22 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h17 == io_wa) begin
        _T_26_23 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h18 == io_wa) begin
        _T_26_24 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h19 == io_wa) begin
        _T_26_25 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1a == io_wa) begin
        _T_26_26 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1b == io_wa) begin
        _T_26_27 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1c == io_wa) begin
        _T_26_28 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1d == io_wa) begin
        _T_26_29 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1e == io_wa) begin
        _T_26_30 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1f == io_wa) begin
        _T_26_31 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h20 == io_wa) begin
        _T_26_32 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h21 == io_wa) begin
        _T_26_33 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h22 == io_wa) begin
        _T_26_34 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h23 == io_wa) begin
        _T_26_35 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h24 == io_wa) begin
        _T_26_36 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h25 == io_wa) begin
        _T_26_37 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h26 == io_wa) begin
        _T_26_38 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h27 == io_wa) begin
        _T_26_39 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h28 == io_wa) begin
        _T_26_40 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h29 == io_wa) begin
        _T_26_41 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2a == io_wa) begin
        _T_26_42 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2b == io_wa) begin
        _T_26_43 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2c == io_wa) begin
        _T_26_44 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2d == io_wa) begin
        _T_26_45 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2e == io_wa) begin
        _T_26_46 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2f == io_wa) begin
        _T_26_47 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h30 == io_wa) begin
        _T_26_48 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h31 == io_wa) begin
        _T_26_49 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h32 == io_wa) begin
        _T_26_50 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h33 == io_wa) begin
        _T_26_51 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h34 == io_wa) begin
        _T_26_52 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h35 == io_wa) begin
        _T_26_53 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h36 == io_wa) begin
        _T_26_54 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h37 == io_wa) begin
        _T_26_55 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h38 == io_wa) begin
        _T_26_56 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h39 == io_wa) begin
        _T_26_57 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3a == io_wa) begin
        _T_26_58 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3b == io_wa) begin
        _T_26_59 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3c == io_wa) begin
        _T_26_60 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3d == io_wa) begin
        _T_26_61 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3e == io_wa) begin
        _T_26_62 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3f == io_wa) begin
        _T_26_63 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h40 == io_wa) begin
        _T_26_64 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h41 == io_wa) begin
        _T_26_65 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h42 == io_wa) begin
        _T_26_66 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h43 == io_wa) begin
        _T_26_67 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h44 == io_wa) begin
        _T_26_68 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h45 == io_wa) begin
        _T_26_69 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h46 == io_wa) begin
        _T_26_70 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h47 == io_wa) begin
        _T_26_71 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h48 == io_wa) begin
        _T_26_72 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h49 == io_wa) begin
        _T_26_73 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4a == io_wa) begin
        _T_26_74 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4b == io_wa) begin
        _T_26_75 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4c == io_wa) begin
        _T_26_76 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4d == io_wa) begin
        _T_26_77 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4e == io_wa) begin
        _T_26_78 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4f == io_wa) begin
        _T_26_79 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h50 == io_wa) begin
        _T_26_80 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h51 == io_wa) begin
        _T_26_81 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h52 == io_wa) begin
        _T_26_82 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h53 == io_wa) begin
        _T_26_83 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h54 == io_wa) begin
        _T_26_84 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h55 == io_wa) begin
        _T_26_85 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h56 == io_wa) begin
        _T_26_86 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h57 == io_wa) begin
        _T_26_87 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h58 == io_wa) begin
        _T_26_88 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h59 == io_wa) begin
        _T_26_89 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5a == io_wa) begin
        _T_26_90 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5b == io_wa) begin
        _T_26_91 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5c == io_wa) begin
        _T_26_92 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5d == io_wa) begin
        _T_26_93 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5e == io_wa) begin
        _T_26_94 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5f == io_wa) begin
        _T_26_95 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h60 == io_wa) begin
        _T_26_96 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h61 == io_wa) begin
        _T_26_97 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h62 == io_wa) begin
        _T_26_98 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h63 == io_wa) begin
        _T_26_99 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h64 == io_wa) begin
        _T_26_100 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h65 == io_wa) begin
        _T_26_101 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h66 == io_wa) begin
        _T_26_102 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h67 == io_wa) begin
        _T_26_103 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h68 == io_wa) begin
        _T_26_104 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h69 == io_wa) begin
        _T_26_105 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6a == io_wa) begin
        _T_26_106 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6b == io_wa) begin
        _T_26_107 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6c == io_wa) begin
        _T_26_108 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6d == io_wa) begin
        _T_26_109 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6e == io_wa) begin
        _T_26_110 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6f == io_wa) begin
        _T_26_111 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h70 == io_wa) begin
        _T_26_112 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h71 == io_wa) begin
        _T_26_113 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h72 == io_wa) begin
        _T_26_114 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h73 == io_wa) begin
        _T_26_115 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h74 == io_wa) begin
        _T_26_116 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h75 == io_wa) begin
        _T_26_117 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h76 == io_wa) begin
        _T_26_118 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h77 == io_wa) begin
        _T_26_119 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h78 == io_wa) begin
        _T_26_120 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h79 == io_wa) begin
        _T_26_121 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7a == io_wa) begin
        _T_26_122 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7b == io_wa) begin
        _T_26_123 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7c == io_wa) begin
        _T_26_124 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7d == io_wa) begin
        _T_26_125 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7e == io_wa) begin
        _T_26_126 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7f == io_wa) begin
        _T_26_127 <= io_di;
      end
    end
    if (io_re) begin
      _T_158 <= io_ra;
    end
    if (io_ore) begin
      if (7'h7f == _T_158) begin
        _T_160 <= _T_26_127;
      end else begin
        if (7'h7e == _T_158) begin
          _T_160 <= _T_26_126;
        end else begin
          if (7'h7d == _T_158) begin
            _T_160 <= _T_26_125;
          end else begin
            if (7'h7c == _T_158) begin
              _T_160 <= _T_26_124;
            end else begin
              if (7'h7b == _T_158) begin
                _T_160 <= _T_26_123;
              end else begin
                if (7'h7a == _T_158) begin
                  _T_160 <= _T_26_122;
                end else begin
                  if (7'h79 == _T_158) begin
                    _T_160 <= _T_26_121;
                  end else begin
                    if (7'h78 == _T_158) begin
                      _T_160 <= _T_26_120;
                    end else begin
                      if (7'h77 == _T_158) begin
                        _T_160 <= _T_26_119;
                      end else begin
                        if (7'h76 == _T_158) begin
                          _T_160 <= _T_26_118;
                        end else begin
                          if (7'h75 == _T_158) begin
                            _T_160 <= _T_26_117;
                          end else begin
                            if (7'h74 == _T_158) begin
                              _T_160 <= _T_26_116;
                            end else begin
                              if (7'h73 == _T_158) begin
                                _T_160 <= _T_26_115;
                              end else begin
                                if (7'h72 == _T_158) begin
                                  _T_160 <= _T_26_114;
                                end else begin
                                  if (7'h71 == _T_158) begin
                                    _T_160 <= _T_26_113;
                                  end else begin
                                    if (7'h70 == _T_158) begin
                                      _T_160 <= _T_26_112;
                                    end else begin
                                      if (7'h6f == _T_158) begin
                                        _T_160 <= _T_26_111;
                                      end else begin
                                        if (7'h6e == _T_158) begin
                                          _T_160 <= _T_26_110;
                                        end else begin
                                          if (7'h6d == _T_158) begin
                                            _T_160 <= _T_26_109;
                                          end else begin
                                            if (7'h6c == _T_158) begin
                                              _T_160 <= _T_26_108;
                                            end else begin
                                              if (7'h6b == _T_158) begin
                                                _T_160 <= _T_26_107;
                                              end else begin
                                                if (7'h6a == _T_158) begin
                                                  _T_160 <= _T_26_106;
                                                end else begin
                                                  if (7'h69 == _T_158) begin
                                                    _T_160 <= _T_26_105;
                                                  end else begin
                                                    if (7'h68 == _T_158) begin
                                                      _T_160 <= _T_26_104;
                                                    end else begin
                                                      if (7'h67 == _T_158) begin
                                                        _T_160 <= _T_26_103;
                                                      end else begin
                                                        if (7'h66 == _T_158) begin
                                                          _T_160 <= _T_26_102;
                                                        end else begin
                                                          if (7'h65 == _T_158) begin
                                                            _T_160 <= _T_26_101;
                                                          end else begin
                                                            if (7'h64 == _T_158) begin
                                                              _T_160 <= _T_26_100;
                                                            end else begin
                                                              if (7'h63 == _T_158) begin
                                                                _T_160 <= _T_26_99;
                                                              end else begin
                                                                if (7'h62 == _T_158) begin
                                                                  _T_160 <= _T_26_98;
                                                                end else begin
                                                                  if (7'h61 == _T_158) begin
                                                                    _T_160 <= _T_26_97;
                                                                  end else begin
                                                                    if (7'h60 == _T_158) begin
                                                                      _T_160 <= _T_26_96;
                                                                    end else begin
                                                                      if (7'h5f == _T_158) begin
                                                                        _T_160 <= _T_26_95;
                                                                      end else begin
                                                                        if (7'h5e == _T_158) begin
                                                                          _T_160 <= _T_26_94;
                                                                        end else begin
                                                                          if (7'h5d == _T_158) begin
                                                                            _T_160 <= _T_26_93;
                                                                          end else begin
                                                                            if (7'h5c == _T_158) begin
                                                                              _T_160 <= _T_26_92;
                                                                            end else begin
                                                                              if (7'h5b == _T_158) begin
                                                                                _T_160 <= _T_26_91;
                                                                              end else begin
                                                                                if (7'h5a == _T_158) begin
                                                                                  _T_160 <= _T_26_90;
                                                                                end else begin
                                                                                  if (7'h59 == _T_158) begin
                                                                                    _T_160 <= _T_26_89;
                                                                                  end else begin
                                                                                    if (7'h58 == _T_158) begin
                                                                                      _T_160 <= _T_26_88;
                                                                                    end else begin
                                                                                      if (7'h57 == _T_158) begin
                                                                                        _T_160 <= _T_26_87;
                                                                                      end else begin
                                                                                        if (7'h56 == _T_158) begin
                                                                                          _T_160 <= _T_26_86;
                                                                                        end else begin
                                                                                          if (7'h55 == _T_158) begin
                                                                                            _T_160 <= _T_26_85;
                                                                                          end else begin
                                                                                            if (7'h54 == _T_158) begin
                                                                                              _T_160 <= _T_26_84;
                                                                                            end else begin
                                                                                              if (7'h53 == _T_158) begin
                                                                                                _T_160 <= _T_26_83;
                                                                                              end else begin
                                                                                                if (7'h52 == _T_158) begin
                                                                                                  _T_160 <= _T_26_82;
                                                                                                end else begin
                                                                                                  if (7'h51 == _T_158) begin
                                                                                                    _T_160 <= _T_26_81;
                                                                                                  end else begin
                                                                                                    if (7'h50 == _T_158) begin
                                                                                                      _T_160 <= _T_26_80;
                                                                                                    end else begin
                                                                                                      if (7'h4f == _T_158) begin
                                                                                                        _T_160 <= _T_26_79;
                                                                                                      end else begin
                                                                                                        if (7'h4e == _T_158) begin
                                                                                                          _T_160 <= _T_26_78;
                                                                                                        end else begin
                                                                                                          if (7'h4d == _T_158) begin
                                                                                                            _T_160 <= _T_26_77;
                                                                                                          end else begin
                                                                                                            if (7'h4c == _T_158) begin
                                                                                                              _T_160 <= _T_26_76;
                                                                                                            end else begin
                                                                                                              if (7'h4b == _T_158) begin
                                                                                                                _T_160 <= _T_26_75;
                                                                                                              end else begin
                                                                                                                if (7'h4a == _T_158) begin
                                                                                                                  _T_160 <= _T_26_74;
                                                                                                                end else begin
                                                                                                                  if (7'h49 == _T_158) begin
                                                                                                                    _T_160 <= _T_26_73;
                                                                                                                  end else begin
                                                                                                                    if (7'h48 == _T_158) begin
                                                                                                                      _T_160 <= _T_26_72;
                                                                                                                    end else begin
                                                                                                                      if (7'h47 == _T_158) begin
                                                                                                                        _T_160 <= _T_26_71;
                                                                                                                      end else begin
                                                                                                                        if (7'h46 == _T_158) begin
                                                                                                                          _T_160 <= _T_26_70;
                                                                                                                        end else begin
                                                                                                                          if (7'h45 == _T_158) begin
                                                                                                                            _T_160 <= _T_26_69;
                                                                                                                          end else begin
                                                                                                                            if (7'h44 == _T_158) begin
                                                                                                                              _T_160 <= _T_26_68;
                                                                                                                            end else begin
                                                                                                                              if (7'h43 == _T_158) begin
                                                                                                                                _T_160 <= _T_26_67;
                                                                                                                              end else begin
                                                                                                                                if (7'h42 == _T_158) begin
                                                                                                                                  _T_160 <= _T_26_66;
                                                                                                                                end else begin
                                                                                                                                  if (7'h41 == _T_158) begin
                                                                                                                                    _T_160 <= _T_26_65;
                                                                                                                                  end else begin
                                                                                                                                    if (7'h40 == _T_158) begin
                                                                                                                                      _T_160 <= _T_26_64;
                                                                                                                                    end else begin
                                                                                                                                      if (7'h3f == _T_158) begin
                                                                                                                                        _T_160 <= _T_26_63;
                                                                                                                                      end else begin
                                                                                                                                        if (7'h3e == _T_158) begin
                                                                                                                                          _T_160 <= _T_26_62;
                                                                                                                                        end else begin
                                                                                                                                          if (7'h3d == _T_158) begin
                                                                                                                                            _T_160 <= _T_26_61;
                                                                                                                                          end else begin
                                                                                                                                            if (7'h3c == _T_158) begin
                                                                                                                                              _T_160 <= _T_26_60;
                                                                                                                                            end else begin
                                                                                                                                              if (7'h3b == _T_158) begin
                                                                                                                                                _T_160 <= _T_26_59;
                                                                                                                                              end else begin
                                                                                                                                                if (7'h3a == _T_158) begin
                                                                                                                                                  _T_160 <= _T_26_58;
                                                                                                                                                end else begin
                                                                                                                                                  if (7'h39 == _T_158) begin
                                                                                                                                                    _T_160 <= _T_26_57;
                                                                                                                                                  end else begin
                                                                                                                                                    if (7'h38 == _T_158) begin
                                                                                                                                                      _T_160 <= _T_26_56;
                                                                                                                                                    end else begin
                                                                                                                                                      if (7'h37 == _T_158) begin
                                                                                                                                                        _T_160 <= _T_26_55;
                                                                                                                                                      end else begin
                                                                                                                                                        if (7'h36 == _T_158) begin
                                                                                                                                                          _T_160 <= _T_26_54;
                                                                                                                                                        end else begin
                                                                                                                                                          if (7'h35 == _T_158) begin
                                                                                                                                                            _T_160 <= _T_26_53;
                                                                                                                                                          end else begin
                                                                                                                                                            if (7'h34 == _T_158) begin
                                                                                                                                                              _T_160 <= _T_26_52;
                                                                                                                                                            end else begin
                                                                                                                                                              if (7'h33 == _T_158) begin
                                                                                                                                                                _T_160 <= _T_26_51;
                                                                                                                                                              end else begin
                                                                                                                                                                if (7'h32 == _T_158) begin
                                                                                                                                                                  _T_160 <= _T_26_50;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (7'h31 == _T_158) begin
                                                                                                                                                                    _T_160 <= _T_26_49;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (7'h30 == _T_158) begin
                                                                                                                                                                      _T_160 <= _T_26_48;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (7'h2f == _T_158) begin
                                                                                                                                                                        _T_160 <= _T_26_47;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (7'h2e == _T_158) begin
                                                                                                                                                                          _T_160 <= _T_26_46;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (7'h2d == _T_158) begin
                                                                                                                                                                            _T_160 <= _T_26_45;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (7'h2c == _T_158) begin
                                                                                                                                                                              _T_160 <= _T_26_44;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (7'h2b == _T_158) begin
                                                                                                                                                                                _T_160 <= _T_26_43;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (7'h2a == _T_158) begin
                                                                                                                                                                                  _T_160 <= _T_26_42;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (7'h29 == _T_158) begin
                                                                                                                                                                                    _T_160 <= _T_26_41;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (7'h28 == _T_158) begin
                                                                                                                                                                                      _T_160 <= _T_26_40;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (7'h27 == _T_158) begin
                                                                                                                                                                                        _T_160 <= _T_26_39;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (7'h26 == _T_158) begin
                                                                                                                                                                                          _T_160 <= _T_26_38;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (7'h25 == _T_158) begin
                                                                                                                                                                                            _T_160 <= _T_26_37;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (7'h24 == _T_158) begin
                                                                                                                                                                                              _T_160 <= _T_26_36;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (7'h23 == _T_158) begin
                                                                                                                                                                                                _T_160 <= _T_26_35;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (7'h22 == _T_158) begin
                                                                                                                                                                                                  _T_160 <= _T_26_34;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (7'h21 == _T_158) begin
                                                                                                                                                                                                    _T_160 <= _T_26_33;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (7'h20 == _T_158) begin
                                                                                                                                                                                                      _T_160 <= _T_26_32;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (7'h1f == _T_158) begin
                                                                                                                                                                                                        _T_160 <= _T_26_31;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (7'h1e == _T_158) begin
                                                                                                                                                                                                          _T_160 <= _T_26_30;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (7'h1d == _T_158) begin
                                                                                                                                                                                                            _T_160 <= _T_26_29;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (7'h1c == _T_158) begin
                                                                                                                                                                                                              _T_160 <= _T_26_28;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (7'h1b == _T_158) begin
                                                                                                                                                                                                                _T_160 <= _T_26_27;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (7'h1a == _T_158) begin
                                                                                                                                                                                                                  _T_160 <= _T_26_26;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (7'h19 == _T_158) begin
                                                                                                                                                                                                                    _T_160 <= _T_26_25;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (7'h18 == _T_158) begin
                                                                                                                                                                                                                      _T_160 <= _T_26_24;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (7'h17 == _T_158) begin
                                                                                                                                                                                                                        _T_160 <= _T_26_23;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (7'h16 == _T_158) begin
                                                                                                                                                                                                                          _T_160 <= _T_26_22;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (7'h15 == _T_158) begin
                                                                                                                                                                                                                            _T_160 <= _T_26_21;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (7'h14 == _T_158) begin
                                                                                                                                                                                                                              _T_160 <= _T_26_20;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (7'h13 == _T_158) begin
                                                                                                                                                                                                                                _T_160 <= _T_26_19;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (7'h12 == _T_158) begin
                                                                                                                                                                                                                                  _T_160 <= _T_26_18;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (7'h11 == _T_158) begin
                                                                                                                                                                                                                                    _T_160 <= _T_26_17;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (7'h10 == _T_158) begin
                                                                                                                                                                                                                                      _T_160 <= _T_26_16;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (7'hf == _T_158) begin
                                                                                                                                                                                                                                        _T_160 <= _T_26_15;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (7'he == _T_158) begin
                                                                                                                                                                                                                                          _T_160 <= _T_26_14;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (7'hd == _T_158) begin
                                                                                                                                                                                                                                            _T_160 <= _T_26_13;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (7'hc == _T_158) begin
                                                                                                                                                                                                                                              _T_160 <= _T_26_12;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (7'hb == _T_158) begin
                                                                                                                                                                                                                                                _T_160 <= _T_26_11;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (7'ha == _T_158) begin
                                                                                                                                                                                                                                                  _T_160 <= _T_26_10;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (7'h9 == _T_158) begin
                                                                                                                                                                                                                                                    _T_160 <= _T_26_9;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (7'h8 == _T_158) begin
                                                                                                                                                                                                                                                      _T_160 <= _T_26_8;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (7'h7 == _T_158) begin
                                                                                                                                                                                                                                                        _T_160 <= _T_26_7;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (7'h6 == _T_158) begin
                                                                                                                                                                                                                                                          _T_160 <= _T_26_6;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (7'h5 == _T_158) begin
                                                                                                                                                                                                                                                            _T_160 <= _T_26_5;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (7'h4 == _T_158) begin
                                                                                                                                                                                                                                                              _T_160 <= _T_26_4;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (7'h3 == _T_158) begin
                                                                                                                                                                                                                                                                _T_160 <= _T_26_3;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (7'h2 == _T_158) begin
                                                                                                                                                                                                                                                                  _T_160 <= _T_26_2;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  if (7'h1 == _T_158) begin
                                                                                                                                                                                                                                                                    _T_160 <= _T_26_1;
                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                    _T_160 <= _T_26_0;
                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_fifo_1( // @[:@2391.2]
  input        clock, // @[:@2392.4]
  input        reset, // @[:@2393.4]
  input        io_clk, // @[:@2394.4]
  input        io_wr_pvld, // @[:@2394.4]
  output       io_wr_prdy, // @[:@2394.4]
  input  [5:0] io_wr_pd, // @[:@2394.4]
  output       io_rd_pvld, // @[:@2394.4]
  input        io_rd_prdy, // @[:@2394.4]
  output [5:0] io_rd_pd // @[:@2394.4]
);
  wire  nv_ram_rwsp_io_clk; // @[FIFO.scala 270:29:@2468.4]
  wire  nv_ram_rwsp_io_re; // @[FIFO.scala 270:29:@2468.4]
  wire  nv_ram_rwsp_io_we; // @[FIFO.scala 270:29:@2468.4]
  wire  nv_ram_rwsp_io_ore; // @[FIFO.scala 270:29:@2468.4]
  wire [6:0] nv_ram_rwsp_io_ra; // @[FIFO.scala 270:29:@2468.4]
  wire [6:0] nv_ram_rwsp_io_wa; // @[FIFO.scala 270:29:@2468.4]
  wire [5:0] nv_ram_rwsp_io_di; // @[FIFO.scala 270:29:@2468.4]
  wire [5:0] nv_ram_rwsp_io_dout; // @[FIFO.scala 270:29:@2468.4]
  reg  _T_26; // @[FIFO.scala 156:56:@2403.4]
  reg [31:0] _RAND_0;
  reg  _T_29; // @[FIFO.scala 158:52:@2404.4]
  reg [31:0] _RAND_1;
  reg [5:0] _T_31; // @[FIFO.scala 159:64:@2405.4]
  reg [31:0] _RAND_2;
  reg  _T_34; // @[FIFO.scala 160:52:@2406.4]
  reg [31:0] _RAND_3;
  wire  _T_125; // @[FIFO.scala 331:38:@2499.4]
  wire  _T_54; // @[FIFO.scala 183:39:@2427.4]
  wire  _T_55; // @[FIFO.scala 183:36:@2428.4]
  reg [7:0] _T_60; // @[FIFO.scala 186:53:@2431.4]
  reg [31:0] _RAND_4;
  wire [8:0] _T_67; // @[FIFO.scala 191:69:@2436.4]
  wire [7:0] _T_68; // @[FIFO.scala 191:69:@2437.4]
  wire [7:0] _T_69; // @[FIFO.scala 191:46:@2438.4]
  wire  _T_72; // @[FIFO.scala 194:80:@2440.4]
  wire  _T_74; // @[FIFO.scala 195:40:@2441.4]
  wire [8:0] _T_62; // @[FIFO.scala 190:76:@2432.4]
  wire [8:0] _T_63; // @[FIFO.scala 190:76:@2433.4]
  wire [7:0] _T_64; // @[FIFO.scala 190:76:@2434.4]
  wire [7:0] _T_65; // @[FIFO.scala 190:43:@2435.4]
  wire [7:0] _T_70; // @[FIFO.scala 192:32:@2439.4]
  wire  _T_37; // @[FIFO.scala 166:60:@2408.4]
  wire  _T_39; // @[FIFO.scala 166:80:@2409.4]
  wire  _T_40; // @[FIFO.scala 166:77:@2410.4]
  wire  _T_41; // @[FIFO.scala 167:38:@2411.4]
  wire  _T_42; // @[FIFO.scala 168:45:@2412.4]
  wire  _T_44; // @[FIFO.scala 171:18:@2414.4]
  wire  _T_46; // @[FIFO.scala 172:45:@2416.6]
  wire  _T_47; // @[FIFO.scala 172:42:@2417.6]
  wire  _GEN_0; // @[FIFO.scala 171:34:@2415.4]
  wire  _T_50; // @[FIFO.scala 176:34:@2421.4]
  wire  _T_82; // @[FIFO.scala 202:27:@2449.4]
  wire [7:0] _GEN_2; // @[FIFO.scala 202:40:@2450.4]
  reg [6:0] _T_85; // @[FIFO.scala 215:68:@2453.4]
  reg [31:0] _RAND_5;
  wire [7:0] _T_87; // @[FIFO.scala 217:42:@2454.4]
  wire [6:0] _T_88; // @[FIFO.scala 217:42:@2455.4]
  wire [6:0] _GEN_3; // @[FIFO.scala 218:29:@2456.4]
  reg [6:0] _T_93; // @[FIFO.scala 224:63:@2460.4]
  reg [31:0] _RAND_6;
  wire [7:0] _T_95; // @[FIFO.scala 225:42:@2461.4]
  wire [6:0] _T_96; // @[FIFO.scala 225:42:@2462.4]
  wire [6:0] _GEN_4; // @[FIFO.scala 227:29:@2463.4]
  reg  _T_104; // @[FIFO.scala 289:73:@2482.4]
  reg [31:0] _RAND_7;
  reg  _T_107; // @[FIFO.scala 295:72:@2484.4]
  reg [31:0] _RAND_8;
  reg  _T_110; // @[FIFO.scala 297:97:@2485.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_113; // @[FIFO.scala 299:53:@2486.4]
  reg [31:0] _RAND_10;
  wire [8:0] _T_115; // @[FIFO.scala 300:74:@2487.4]
  wire [8:0] _T_116; // @[FIFO.scala 300:74:@2488.4]
  wire [7:0] _T_117; // @[FIFO.scala 300:74:@2489.4]
  wire [7:0] _T_118; // @[FIFO.scala 300:43:@2490.4]
  wire [8:0] _T_120; // @[FIFO.scala 301:68:@2491.4]
  wire [7:0] _T_121; // @[FIFO.scala 301:68:@2492.4]
  wire [7:0] _T_122; // @[FIFO.scala 301:46:@2493.4]
  wire [7:0] _T_123; // @[FIFO.scala 302:32:@2494.4]
  wire  _T_124; // @[FIFO.scala 303:25:@2495.4]
  wire [7:0] _GEN_5; // @[FIFO.scala 303:39:@2496.4]
  wire  _T_127; // @[FIFO.scala 333:77:@2501.4]
  wire  _T_129; // @[FIFO.scala 334:83:@2502.4]
  wire  _T_130; // @[FIFO.scala 335:44:@2503.4]
  wire  _T_131; // @[FIFO.scala 336:60:@2504.4]
  wire  _T_133; // @[FIFO.scala 336:81:@2506.4]
  wire  _GEN_6; // @[FIFO.scala 338:43:@2510.4]
  wire  _T_137; // @[FIFO.scala 341:66:@2513.4]
  wire  _T_138; // @[FIFO.scala 341:63:@2514.4]
  wire  _T_139; // @[FIFO.scala 341:43:@2515.4]
  nv_ram_rwsp_1 nv_ram_rwsp ( // @[FIFO.scala 270:29:@2468.4]
    .io_clk(nv_ram_rwsp_io_clk),
    .io_re(nv_ram_rwsp_io_re),
    .io_we(nv_ram_rwsp_io_we),
    .io_ore(nv_ram_rwsp_io_ore),
    .io_ra(nv_ram_rwsp_io_ra),
    .io_wa(nv_ram_rwsp_io_wa),
    .io_di(nv_ram_rwsp_io_di),
    .io_dout(nv_ram_rwsp_io_dout)
  );
  assign _T_125 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 331:38:@2499.4]
  assign _T_54 = _T_26 == 1'h0; // @[FIFO.scala 183:39:@2427.4]
  assign _T_55 = _T_29 & _T_54; // @[FIFO.scala 183:36:@2428.4]
  assign _T_67 = _T_60 + 8'h1; // @[FIFO.scala 191:69:@2436.4]
  assign _T_68 = _T_60 + 8'h1; // @[FIFO.scala 191:69:@2437.4]
  assign _T_69 = _T_55 ? _T_68 : _T_60; // @[FIFO.scala 191:46:@2438.4]
  assign _T_72 = _T_69 == 8'h80; // @[FIFO.scala 194:80:@2440.4]
  assign _T_74 = _T_125 ? 1'h0 : _T_72; // @[FIFO.scala 195:40:@2441.4]
  assign _T_62 = _T_60 - 8'h1; // @[FIFO.scala 190:76:@2432.4]
  assign _T_63 = $unsigned(_T_62); // @[FIFO.scala 190:76:@2433.4]
  assign _T_64 = _T_63[7:0]; // @[FIFO.scala 190:76:@2434.4]
  assign _T_65 = _T_55 ? _T_60 : _T_64; // @[FIFO.scala 190:43:@2435.4]
  assign _T_70 = _T_125 ? _T_65 : _T_69; // @[FIFO.scala 192:32:@2439.4]
  assign _T_37 = _T_29 & _T_74; // @[FIFO.scala 166:60:@2408.4]
  assign _T_39 = _T_55 == 1'h0; // @[FIFO.scala 166:80:@2409.4]
  assign _T_40 = _T_37 & _T_39; // @[FIFO.scala 166:77:@2410.4]
  assign _T_41 = io_wr_pvld ? _T_74 : _T_40; // @[FIFO.scala 167:38:@2411.4]
  assign _T_42 = _T_29 & _T_26; // @[FIFO.scala 168:45:@2412.4]
  assign _T_44 = _T_42 == 1'h0; // @[FIFO.scala 171:18:@2414.4]
  assign _T_46 = _T_34 == 1'h0; // @[FIFO.scala 172:45:@2416.6]
  assign _T_47 = io_wr_pvld & _T_46; // @[FIFO.scala 172:42:@2417.6]
  assign _GEN_0 = _T_44 ? _T_47 : _T_29; // @[FIFO.scala 171:34:@2415.4]
  assign _T_50 = _T_46 & io_wr_pvld; // @[FIFO.scala 176:34:@2421.4]
  assign _T_82 = _T_55 ^ _T_125; // @[FIFO.scala 202:27:@2449.4]
  assign _GEN_2 = _T_82 ? _T_70 : _T_60; // @[FIFO.scala 202:40:@2450.4]
  assign _T_87 = _T_85 + 7'h1; // @[FIFO.scala 217:42:@2454.4]
  assign _T_88 = _T_85 + 7'h1; // @[FIFO.scala 217:42:@2455.4]
  assign _GEN_3 = _T_55 ? _T_88 : _T_85; // @[FIFO.scala 218:29:@2456.4]
  assign _T_95 = _T_93 + 7'h1; // @[FIFO.scala 225:42:@2461.4]
  assign _T_96 = _T_93 + 7'h1; // @[FIFO.scala 225:42:@2462.4]
  assign _GEN_4 = _T_125 ? _T_96 : _T_93; // @[FIFO.scala 227:29:@2463.4]
  assign _T_115 = _T_113 - 8'h1; // @[FIFO.scala 300:74:@2487.4]
  assign _T_116 = $unsigned(_T_115); // @[FIFO.scala 300:74:@2488.4]
  assign _T_117 = _T_116[7:0]; // @[FIFO.scala 300:74:@2489.4]
  assign _T_118 = _T_104 ? _T_113 : _T_117; // @[FIFO.scala 300:43:@2490.4]
  assign _T_120 = _T_113 + 8'h1; // @[FIFO.scala 301:68:@2491.4]
  assign _T_121 = _T_113 + 8'h1; // @[FIFO.scala 301:68:@2492.4]
  assign _T_122 = _T_104 ? _T_121 : _T_113; // @[FIFO.scala 301:46:@2493.4]
  assign _T_123 = _T_125 ? _T_118 : _T_122; // @[FIFO.scala 302:32:@2494.4]
  assign _T_124 = _T_104 | _T_125; // @[FIFO.scala 303:25:@2495.4]
  assign _GEN_5 = _T_124 ? _T_123 : _T_113; // @[FIFO.scala 303:39:@2496.4]
  assign _T_127 = _T_118 != 8'h0; // @[FIFO.scala 333:77:@2501.4]
  assign _T_129 = _T_122 != 8'h0; // @[FIFO.scala 334:83:@2502.4]
  assign _T_130 = _T_125 ? _T_127 : _T_129; // @[FIFO.scala 335:44:@2503.4]
  assign _T_131 = ~ _T_107; // @[FIFO.scala 336:60:@2504.4]
  assign _T_133 = _T_131 | _T_125; // @[FIFO.scala 336:81:@2506.4]
  assign _GEN_6 = _T_124 ? _T_130 : _T_107; // @[FIFO.scala 338:43:@2510.4]
  assign _T_137 = io_rd_prdy == 1'h0; // @[FIFO.scala 341:66:@2513.4]
  assign _T_138 = _T_110 & _T_137; // @[FIFO.scala 341:63:@2514.4]
  assign _T_139 = _T_107 | _T_138; // @[FIFO.scala 341:43:@2515.4]
  assign io_wr_prdy = _T_34 == 1'h0; // @[FIFO.scala 182:20:@2426.4]
  assign io_rd_pvld = _T_110; // @[FIFO.scala 344:24:@2517.4]
  assign io_rd_pd = nv_ram_rwsp_io_dout; // @[FIFO.scala 345:22:@2518.4]
  assign nv_ram_rwsp_io_clk = io_clk; // @[FIFO.scala 271:24:@2471.4]
  assign nv_ram_rwsp_io_re = _T_130 & _T_133; // @[FIFO.scala 279:23:@2478.4]
  assign nv_ram_rwsp_io_we = _T_29 & _T_54; // @[FIFO.scala 276:23:@2474.4]
  assign nv_ram_rwsp_io_ore = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 280:24:@2479.4]
  assign nv_ram_rwsp_io_ra = _T_125 ? _T_96 : _T_93; // @[FIFO.scala 278:23:@2477.4]
  assign nv_ram_rwsp_io_wa = _T_85; // @[FIFO.scala 274:27:@2473.4]
  assign nv_ram_rwsp_io_di = _T_31; // @[FIFO.scala 277:23:@2475.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_31 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_34 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_60 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_85 = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_93 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_104 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_107 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_110 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_113 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_125) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_72;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_29 <= _T_47;
      end
    end
    if (_T_50) begin
      _T_31 <= io_wr_pd;
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (io_wr_pvld) begin
        if (_T_125) begin
          _T_34 <= 1'h0;
        end else begin
          _T_34 <= _T_72;
        end
      end else begin
        _T_34 <= _T_40;
      end
    end
    if (reset) begin
      _T_60 <= 8'h0;
    end else begin
      if (_T_82) begin
        if (_T_125) begin
          if (!(_T_55)) begin
            _T_60 <= _T_64;
          end
        end else begin
          if (_T_55) begin
            _T_60 <= _T_68;
          end
        end
      end
    end
    if (reset) begin
      _T_85 <= 7'h0;
    end else begin
      if (_T_55) begin
        _T_85 <= _T_88;
      end
    end
    if (reset) begin
      _T_93 <= 7'h0;
    end else begin
      if (_T_125) begin
        _T_93 <= _T_96;
      end
    end
    if (reset) begin
      _T_104 <= 1'h0;
    end else begin
      _T_104 <= _T_55;
    end
    if (reset) begin
      _T_107 <= 1'h0;
    end else begin
      if (_T_124) begin
        if (_T_125) begin
          _T_107 <= _T_127;
        end else begin
          _T_107 <= _T_129;
        end
      end
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      _T_110 <= _T_139;
    end
    if (reset) begin
      _T_113 <= 8'h0;
    end else begin
      if (_T_124) begin
        if (_T_125) begin
          if (!(_T_104)) begin
            _T_113 <= _T_117;
          end
        end else begin
          if (_T_104) begin
            _T_113 <= _T_121;
          end
        end
      end
    end
  end
endmodule
module NV_COUNTER_STAGE_histogram( // @[:@2534.2]
  input         reset, // @[:@2536.4]
  input         io_clk, // @[:@2537.4]
  input         io_rd_stall_inc, // @[:@2537.4]
  input         io_rd_stall_clr, // @[:@2537.4]
  input         io_rd_stall_cen, // @[:@2537.4]
  output [31:0] io_cnt_cur // @[:@2537.4]
);
  reg [31:0] _T_20; // @[Perf_Counter.scala 47:30:@2540.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_34; // @[Perf_Counter.scala 56:28:@2548.4]
  wire [33:0] _T_22; // @[Perf_Counter.scala 48:23:@2541.4 Perf_Counter.scala 55:13:@2547.4]
  wire [33:0] _T_24; // @[Perf_Counter.scala 49:23:@2542.4 Perf_Counter.scala 56:13:@2549.4]
  wire [33:0] _T_45; // @[Perf_Counter.scala 58:19:@2558.4]
  wire [33:0] _T_46; // @[Perf_Counter.scala 61:19:@2560.4]
  wire [33:0] _T_48; // @[Perf_Counter.scala 62:19:@2562.4]
  wire [33:0] _GEN_0; // @[Perf_Counter.scala 65:26:@2564.4]
  assign _T_34 = _T_20 + 32'h1; // @[Perf_Counter.scala 56:28:@2548.4]
  assign _T_22 = {{2'd0}, _T_20}; // @[Perf_Counter.scala 48:23:@2541.4 Perf_Counter.scala 55:13:@2547.4]
  assign _T_24 = {{1'd0}, _T_34}; // @[Perf_Counter.scala 49:23:@2542.4 Perf_Counter.scala 56:13:@2549.4]
  assign _T_45 = io_rd_stall_inc ? _T_24 : _T_22; // @[Perf_Counter.scala 58:19:@2558.4]
  assign _T_46 = io_rd_stall_inc ? _T_45 : _T_22; // @[Perf_Counter.scala 61:19:@2560.4]
  assign _T_48 = io_rd_stall_clr ? 34'h0 : _T_46; // @[Perf_Counter.scala 62:19:@2562.4]
  assign _GEN_0 = io_rd_stall_cen ? _T_48 : {{2'd0}, _T_20}; // @[Perf_Counter.scala 65:26:@2564.4]
  assign io_cnt_cur = _T_20; // @[Perf_Counter.scala 69:16:@2567.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_20 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_20 <= 32'h0;
    end else begin
      _T_20 <= _GEN_0[31:0];
    end
  end
endmodule
module NV_COUNTER_STAGE_histogram_1( // @[:@2569.2]
  input        reset, // @[:@2571.4]
  input        io_clk, // @[:@2572.4]
  input        io_rd_stall_inc, // @[:@2572.4]
  input        io_rd_stall_dec, // @[:@2572.4]
  input        io_rd_stall_clr, // @[:@2572.4]
  input        io_rd_stall_cen, // @[:@2572.4]
  output [8:0] io_cnt_cur // @[:@2572.4]
);
  wire  _T_17; // @[Perf_Counter.scala 44:31:@2574.4]
  reg [8:0] _T_20; // @[Perf_Counter.scala 47:30:@2575.4]
  reg [31:0] _RAND_0;
  wire [9:0] _T_34; // @[Perf_Counter.scala 56:28:@2583.4]
  wire [9:0] _T_36; // @[Perf_Counter.scala 57:28:@2585.4]
  wire [9:0] _T_37; // @[Perf_Counter.scala 57:28:@2586.4]
  wire  _T_39; // @[Perf_Counter.scala 58:39:@2588.4]
  wire  _T_40; // @[Perf_Counter.scala 58:36:@2589.4]
  wire  _T_42; // @[Perf_Counter.scala 59:23:@2590.4]
  wire  _T_43; // @[Perf_Counter.scala 59:40:@2591.4]
  wire [10:0] _T_26; // @[Perf_Counter.scala 50:23:@2578.4 Perf_Counter.scala 57:13:@2587.4]
  wire [10:0] _T_22; // @[Perf_Counter.scala 48:23:@2576.4 Perf_Counter.scala 55:13:@2582.4]
  wire [10:0] _T_44; // @[Perf_Counter.scala 59:22:@2592.4]
  wire [10:0] _T_24; // @[Perf_Counter.scala 49:23:@2577.4 Perf_Counter.scala 56:13:@2584.4]
  wire [10:0] _T_45; // @[Perf_Counter.scala 58:19:@2593.4]
  wire [10:0] _T_46; // @[Perf_Counter.scala 61:19:@2595.4]
  wire [10:0] _T_48; // @[Perf_Counter.scala 62:19:@2597.4]
  wire [10:0] _GEN_0; // @[Perf_Counter.scala 65:26:@2599.4]
  assign _T_17 = io_rd_stall_inc ^ io_rd_stall_dec; // @[Perf_Counter.scala 44:31:@2574.4]
  assign _T_34 = _T_20 + 9'h1; // @[Perf_Counter.scala 56:28:@2583.4]
  assign _T_36 = _T_20 - 9'h1; // @[Perf_Counter.scala 57:28:@2585.4]
  assign _T_37 = $unsigned(_T_36); // @[Perf_Counter.scala 57:28:@2586.4]
  assign _T_39 = io_rd_stall_dec == 1'h0; // @[Perf_Counter.scala 58:39:@2588.4]
  assign _T_40 = io_rd_stall_inc & _T_39; // @[Perf_Counter.scala 58:36:@2589.4]
  assign _T_42 = io_rd_stall_inc == 1'h0; // @[Perf_Counter.scala 59:23:@2590.4]
  assign _T_43 = _T_42 & io_rd_stall_dec; // @[Perf_Counter.scala 59:40:@2591.4]
  assign _T_26 = {{1'd0}, _T_37}; // @[Perf_Counter.scala 50:23:@2578.4 Perf_Counter.scala 57:13:@2587.4]
  assign _T_22 = {{2'd0}, _T_20}; // @[Perf_Counter.scala 48:23:@2576.4 Perf_Counter.scala 55:13:@2582.4]
  assign _T_44 = _T_43 ? _T_26 : _T_22; // @[Perf_Counter.scala 59:22:@2592.4]
  assign _T_24 = {{1'd0}, _T_34}; // @[Perf_Counter.scala 49:23:@2577.4 Perf_Counter.scala 56:13:@2584.4]
  assign _T_45 = _T_40 ? _T_24 : _T_44; // @[Perf_Counter.scala 58:19:@2593.4]
  assign _T_46 = _T_17 ? _T_45 : _T_22; // @[Perf_Counter.scala 61:19:@2595.4]
  assign _T_48 = io_rd_stall_clr ? 11'h0 : _T_46; // @[Perf_Counter.scala 62:19:@2597.4]
  assign _GEN_0 = io_rd_stall_cen ? _T_48 : {{2'd0}, _T_20}; // @[Perf_Counter.scala 65:26:@2599.4]
  assign io_cnt_cur = _T_20; // @[Perf_Counter.scala 69:16:@2602.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_20 = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_20 <= 9'h0;
    end else begin
      _T_20 <= _GEN_0[8:0];
    end
  end
endmodule
module NV_NVDLA_CDMA_wt( // @[:@2604.2]
  input          reset, // @[:@2606.4]
  input          io_nvdla_core_clk, // @[:@2607.4]
  input          io_nvdla_core_ng_clk, // @[:@2607.4]
  input          io_cdma_wt2mcif_rd_req_pd_ready, // @[:@2607.4]
  output         io_cdma_wt2mcif_rd_req_pd_valid, // @[:@2607.4]
  output [78:0]  io_cdma_wt2mcif_rd_req_pd_bits, // @[:@2607.4]
  output         io_mcif2cdma_wt_rd_rsp_pd_ready, // @[:@2607.4]
  input          io_mcif2cdma_wt_rd_rsp_pd_valid, // @[:@2607.4]
  input  [256:0] io_mcif2cdma_wt_rd_rsp_pd_bits, // @[:@2607.4]
  input          io_cdma_wt2cvif_rd_req_pd_ready, // @[:@2607.4]
  output         io_cdma_wt2cvif_rd_req_pd_valid, // @[:@2607.4]
  output [78:0]  io_cdma_wt2cvif_rd_req_pd_bits, // @[:@2607.4]
  output         io_cvif2cdma_wt_rd_rsp_pd_ready, // @[:@2607.4]
  input          io_cvif2cdma_wt_rd_rsp_pd_valid, // @[:@2607.4]
  input  [256:0] io_cvif2cdma_wt_rd_rsp_pd_bits, // @[:@2607.4]
  output [1:0]   io_cdma2buf_wt_wr_sel, // @[:@2607.4]
  output         io_cdma2buf_wt_wr_addr_valid, // @[:@2607.4]
  output [16:0]  io_cdma2buf_wt_wr_addr_bits, // @[:@2607.4]
  output [255:0] io_cdma2buf_wt_wr_data, // @[:@2607.4]
  input          io_status2dma_fsm_switch, // @[:@2607.4]
  output [1:0]   io_wt2status_state, // @[:@2607.4]
  output         io_cdma2sc_wt_updt_valid, // @[:@2607.4]
  output [14:0]  io_cdma2sc_wt_updt_bits_entries, // @[:@2607.4]
  output [13:0]  io_cdma2sc_wt_updt_bits_kernels, // @[:@2607.4]
  output         io_cdma2sc_wt_pending_ack, // @[:@2607.4]
  input          io_sc2cdma_wt_updt_valid, // @[:@2607.4]
  input  [14:0]  io_sc2cdma_wt_updt_bits_entries, // @[:@2607.4]
  input          io_sc2cdma_wt_pending_req, // @[:@2607.4]
  input          io_reg2dp_op_en, // @[:@2607.4]
  input          io_reg2dp_weight_reuse, // @[:@2607.4]
  input          io_reg2dp_skip_weight_rls, // @[:@2607.4]
  input  [17:0]  io_reg2dp_byte_per_kernel, // @[:@2607.4]
  input  [12:0]  io_reg2dp_weight_kernel, // @[:@2607.4]
  input          io_reg2dp_weight_ram_type, // @[:@2607.4]
  input  [26:0]  io_reg2dp_weight_addr_low, // @[:@2607.4]
  input  [31:0]  io_reg2dp_weight_addr_high, // @[:@2607.4]
  input  [31:0]  io_reg2dp_weight_bytes, // @[:@2607.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@2607.4]
  input  [4:0]   io_reg2dp_weight_bank, // @[:@2607.4]
  input          io_reg2dp_dma_en, // @[:@2607.4]
  output         io_dp2reg_wt_flush_done, // @[:@2607.4]
  output [31:0]  io_dp2reg_wt_rd_stall // @[:@2607.4]
);
  wire  NV_NVDLA_DMAIF_rdreq_reset; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type; // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
  wire  NV_NVDLA_DMAIF_rdrsp_reset; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
  wire  NV_NVDLA_fifo_clock; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_reset; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_io_clk; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_io_wr_pvld; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire [256:0] NV_NVDLA_fifo_io_wr_pd; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_io_rd_prdy; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire [256:0] NV_NVDLA_fifo_io_rd_pd; // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
  wire  NV_NVDLA_fifo_1_clock; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_reset; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_io_clk; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_io_wr_pvld; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_io_wr_prdy; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire [5:0] NV_NVDLA_fifo_1_io_wr_pd; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_io_rd_pvld; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_NVDLA_fifo_1_io_rd_prdy; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire [5:0] NV_NVDLA_fifo_1_io_rd_pd; // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
  wire  NV_COUNTER_STAGE_histogram_reset; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire  NV_COUNTER_STAGE_histogram_io_clk; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_inc; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_clr; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_cen; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire [31:0] NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
  wire  NV_COUNTER_STAGE_histogram_1_reset; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_clk; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  wire [8:0] NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
  reg  _T_83; // @[NV_NVDLA_CDMA_wt.scala 97:39:@2612.4]
  reg [31:0] _RAND_0;
  reg [1:0] _T_89; // @[NV_NVDLA_CDMA_wt.scala 99:28:@2613.4]
  reg [31:0] _RAND_1;
  wire  _T_92; // @[Conditional.scala 37:30:@2616.4]
  reg [4:0] _T_105; // @[NV_NVDLA_CDMA_wt.scala 122:33:@2656.4]
  reg [31:0] _RAND_2;
  wire  _T_135; // @[NV_NVDLA_CDMA_wt.scala 133:38:@2672.4]
  reg [4:0] _T_112; // @[NV_NVDLA_CDMA_wt.scala 123:35:@2658.4]
  reg [31:0] _RAND_3;
  wire  _T_136; // @[NV_NVDLA_CDMA_wt.scala 133:83:@2673.4]
  wire  _T_137; // @[NV_NVDLA_CDMA_wt.scala 133:63:@2674.4]
  wire  _T_93; // @[NV_NVDLA_CDMA_wt.scala 104:31:@2618.6]
  wire  _T_94; // @[NV_NVDLA_CDMA_wt.scala 105:36:@2623.8]
  wire  _T_95; // @[NV_NVDLA_CDMA_wt.scala 105:61:@2624.8]
  wire [1:0] _GEN_0; // @[NV_NVDLA_CDMA_wt.scala 106:37:@2629.10]
  wire [1:0] _GEN_1; // @[NV_NVDLA_CDMA_wt.scala 105:85:@2625.8]
  wire [1:0] _GEN_2; // @[NV_NVDLA_CDMA_wt.scala 104:47:@2619.6]
  wire  _T_96; // @[Conditional.scala 37:30:@2634.6]
  reg  _T_147; // @[NV_NVDLA_CDMA_wt.scala 143:33:@2682.4]
  reg [31:0] _RAND_4;
  reg  _T_144; // @[NV_NVDLA_CDMA_wt.scala 142:30:@2681.4]
  reg [31:0] _RAND_5;
  wire  _T_157; // @[NV_NVDLA_CDMA_wt.scala 153:41:@2692.4]
  wire  _T_158; // @[NV_NVDLA_CDMA_wt.scala 153:39:@2693.4]
  wire [1:0] _GEN_3; // @[NV_NVDLA_CDMA_wt.scala 109:32:@2636.8]
  wire  _T_97; // @[Conditional.scala 37:30:@2641.8]
  reg  _T_119; // @[NV_NVDLA_CDMA_wt.scala 126:30:@2661.4]
  reg [31:0] _RAND_6;
  reg [3:0] _T_122; // @[NV_NVDLA_CDMA_wt.scala 127:34:@2662.4]
  reg [31:0] _RAND_7;
  wire  _T_133; // @[NV_NVDLA_CDMA_wt.scala 132:50:@2669.4]
  wire  _T_134; // @[NV_NVDLA_CDMA_wt.scala 132:31:@2670.4]
  wire [1:0] _GEN_4; // @[NV_NVDLA_CDMA_wt.scala 112:27:@2643.10]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@2642.8]
  wire [1:0] _GEN_8; // @[Conditional.scala 39:67:@2635.6]
  wire [1:0] _GEN_9; // @[Conditional.scala 40:58:@2617.4]
  wire  _T_125; // @[NV_NVDLA_CDMA_wt.scala 130:64:@2663.4]
  wire  _T_126; // @[NV_NVDLA_CDMA_wt.scala 130:45:@2664.4]
  wire [4:0] _T_128; // @[NV_NVDLA_CDMA_wt.scala 130:103:@2665.4]
  wire [3:0] _T_129; // @[NV_NVDLA_CDMA_wt.scala 130:103:@2666.4]
  wire [3:0] _T_130; // @[NV_NVDLA_CDMA_wt.scala 130:32:@2667.4]
  wire  _T_151; // @[NV_NVDLA_CDMA_wt.scala 146:47:@2684.4]
  wire  _T_152; // @[NV_NVDLA_CDMA_wt.scala 146:33:@2685.4]
  wire [3:0] _T_131; // @[NV_NVDLA_CDMA_wt.scala 129:32:@2668.4]
  wire  _T_153; // @[NV_NVDLA_CDMA_wt.scala 148:30:@2687.4]
  wire  _T_138; // @[NV_NVDLA_CDMA_wt.scala 135:19:@2676.4]
  wire [3:0] _GEN_10; // @[NV_NVDLA_CDMA_wt.scala 135:32:@2677.4]
  reg [1:0] _T_141; // @[NV_NVDLA_CDMA_wt.scala 141:38:@2680.4]
  reg [31:0] _RAND_8;
  reg  _T_150; // @[NV_NVDLA_CDMA_wt.scala 144:30:@2683.4]
  reg [31:0] _RAND_9;
  wire  _T_154; // @[NV_NVDLA_CDMA_wt.scala 149:33:@2689.4]
  wire  _T_155; // @[NV_NVDLA_CDMA_wt.scala 150:33:@2690.4]
  wire  _T_156; // @[NV_NVDLA_CDMA_wt.scala 151:37:@2691.4]
  wire [4:0] _GEN_11; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  wire [4:0] _GEN_12; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  wire  _GEN_13; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  reg [11:0] _T_168; // @[NV_NVDLA_CDMA_wt.scala 176:24:@2709.4]
  reg [31:0] _RAND_10;
  reg [5:0] _T_175; // @[NV_NVDLA_CDMA_wt.scala 177:30:@2711.4]
  reg [31:0] _RAND_11;
  reg [6:0] _T_182; // @[NV_NVDLA_CDMA_wt.scala 178:34:@2713.4]
  reg [31:0] _RAND_12;
  wire [18:0] _T_187; // @[NV_NVDLA_CDMA_wt.scala 181:63:@2715.4]
  reg [18:0] _T_189; // @[Reg.scala 11:16:@2716.4]
  reg [31:0] _RAND_13;
  wire [6:0] _T_192; // @[NV_NVDLA_CDMA_wt.scala 184:43:@2720.4]
  wire [7:0] _T_194; // @[NV_NVDLA_CDMA_wt.scala 185:28:@2721.4]
  wire [5:0] _T_196; // @[NV_NVDLA_CDMA_wt.scala 186:43:@2722.4]
  wire [5:0] _T_198; // @[NV_NVDLA_CDMA_wt.scala 187:47:@2723.4]
  wire [6:0] _T_199; // @[NV_NVDLA_CDMA_wt.scala 188:43:@2724.4]
  wire [11:0] _GEN_15; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  wire [5:0] _GEN_16; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  wire [6:0] _GEN_17; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  reg [3:0] _T_209; // @[NV_NVDLA_CDMA_wt.scala 205:33:@2734.4]
  reg [31:0] _RAND_14;
  reg [28:0] _T_212; // @[NV_NVDLA_CDMA_wt.scala 206:38:@2735.4]
  reg [31:0] _RAND_15;
  reg  _T_215; // @[NV_NVDLA_CDMA_wt.scala 207:38:@2736.4]
  reg [31:0] _RAND_16;
  wire [28:0] _GEN_63; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2738.4]
  wire [29:0] _T_218; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2738.4]
  wire [29:0] _T_219; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2739.4]
  wire [28:0] _T_220; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2740.4]
  wire [26:0] _T_221; // @[NV_NVDLA_CDMA_wt.scala 212:66:@2741.4]
  wire [28:0] _T_222; // @[NV_NVDLA_CDMA_wt.scala 212:33:@2742.4]
  wire [2:0] _T_224; // @[NV_NVDLA_CDMA_wt.scala 213:92:@2743.4]
  wire [3:0] _GEN_64; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2744.4]
  wire [4:0] _T_225; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2744.4]
  wire [4:0] _T_226; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2745.4]
  wire [3:0] _T_227; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2746.4]
  wire [3:0] _T_229; // @[NV_NVDLA_CDMA_wt.scala 213:37:@2747.4]
  wire [28:0] _GEN_65; // @[NV_NVDLA_CDMA_wt.scala 214:52:@2748.4]
  wire  _T_230; // @[NV_NVDLA_CDMA_wt.scala 214:52:@2748.4]
  wire [3:0] _T_231; // @[NV_NVDLA_CDMA_wt.scala 214:92:@2749.4]
  wire [3:0] _T_232; // @[NV_NVDLA_CDMA_wt.scala 214:28:@2750.4]
  reg  _T_272; // @[NV_NVDLA_CDMA_wt.scala 246:32:@2784.4]
  reg [31:0] _RAND_17;
  wire  _T_308; // @[NV_NVDLA_CDMA_wt.scala 275:48:@2810.4]
  wire  _T_313; // @[NV_NVDLA_CDMA_wt.scala 277:30:@2815.4 NV_NVDLA_CDMA_wt.scala 309:20:@2841.4]
  wire  _T_315; // @[NV_NVDLA_CDMA_wt.scala 278:34:@2816.4 NV_NVDLA_CDMA_wt.scala 399:24:@2936.4]
  wire  _T_316; // @[NV_NVDLA_CDMA_wt.scala 279:41:@2817.4]
  reg [13:0] _T_289; // @[NV_NVDLA_CDMA_wt.scala 266:64:@2798.4]
  reg [31:0] _RAND_18;
  reg [16:0] _T_292; // @[NV_NVDLA_CDMA_wt.scala 267:65:@2799.4]
  reg [31:0] _RAND_19;
  wire [16:0] _GEN_66; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2801.4]
  wire [17:0] _T_296; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2801.4]
  wire [16:0] _T_297; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2802.4]
  reg [16:0] _T_295; // @[NV_NVDLA_CDMA_wt.scala 268:62:@2800.4]
  reg [31:0] _RAND_20;
  wire [17:0] _T_298; // @[NV_NVDLA_CDMA_wt.scala 269:53:@2803.4]
  wire [16:0] _T_299; // @[NV_NVDLA_CDMA_wt.scala 269:53:@2804.4]
  wire [15:0] _T_301; // @[Cat.scala 30:58:@2805.4]
  wire [16:0] _T_303; // @[NV_NVDLA_CDMA_wt.scala 270:115:@2806.4]
  wire  _T_304; // @[NV_NVDLA_CDMA_wt.scala 270:53:@2807.4]
  wire  _T_305; // @[NV_NVDLA_CDMA_wt.scala 270:38:@2808.4]
  wire  _T_317; // @[NV_NVDLA_CDMA_wt.scala 280:42:@2818.4]
  wire  _T_318; // @[NV_NVDLA_CDMA_wt.scala 280:40:@2819.4]
  reg  _T_284; // @[NV_NVDLA_CDMA_wt.scala 250:33:@2788.4]
  reg [31:0] _RAND_21;
  wire  _T_319; // @[NV_NVDLA_CDMA_wt.scala 280:64:@2820.4]
  wire  _T_320; // @[NV_NVDLA_CDMA_wt.scala 280:62:@2821.4]
  wire  _T_321; // @[NV_NVDLA_CDMA_wt.scala 281:34:@2822.4]
  wire  _T_309; // @[NV_NVDLA_CDMA_wt.scala 275:63:@2811.4]
  wire  _T_310; // @[NV_NVDLA_CDMA_wt.scala 275:45:@2812.4]
  wire  _T_311; // @[NV_NVDLA_CDMA_wt.scala 275:31:@2813.4]
  wire [3:0] _GEN_19; // @[NV_NVDLA_CDMA_wt.scala 216:27:@2751.4]
  wire [28:0] _GEN_20; // @[NV_NVDLA_CDMA_wt.scala 216:27:@2751.4]
  reg [58:0] _T_235; // @[NV_NVDLA_CDMA_wt.scala 223:33:@2756.4]
  reg [63:0] _RAND_22;
  reg [3:0] _T_238; // @[NV_NVDLA_CDMA_wt.scala 224:33:@2757.4]
  reg [31:0] _RAND_23;
  reg [2:0] _T_241; // @[NV_NVDLA_CDMA_wt.scala 225:37:@2758.4]
  reg [31:0] _RAND_24;
  reg  _T_244; // @[NV_NVDLA_CDMA_wt.scala 226:33:@2759.4]
  reg [31:0] _RAND_25;
  reg  _T_247; // @[NV_NVDLA_CDMA_wt.scala 227:33:@2760.4]
  reg [31:0] _RAND_26;
  reg  _T_250; // @[NV_NVDLA_CDMA_wt.scala 228:38:@2761.4]
  reg [31:0] _RAND_27;
  wire  _T_251; // @[NV_NVDLA_CDMA_wt.scala 231:69:@2762.4]
  wire  _T_252; // @[NV_NVDLA_CDMA_wt.scala 231:45:@2763.4]
  wire [55:0] _T_253; // @[NV_NVDLA_CDMA_wt.scala 232:41:@2764.4]
  wire [56:0] _T_255; // @[NV_NVDLA_CDMA_wt.scala 232:61:@2765.4]
  wire  _T_256; // @[NV_NVDLA_CDMA_wt.scala 233:29:@2766.4]
  wire [58:0] _T_257; // @[Cat.scala 30:58:@2767.4]
  wire [59:0] _T_259; // @[Cat.scala 30:58:@2768.4]
  wire [59:0] _T_260; // @[NV_NVDLA_CDMA_wt.scala 233:28:@2769.4]
  wire [2:0] _T_261; // @[NV_NVDLA_CDMA_wt.scala 234:43:@2770.4]
  wire [3:0] _T_263; // @[NV_NVDLA_CDMA_wt.scala 234:50:@2771.4]
  wire [3:0] _T_264; // @[NV_NVDLA_CDMA_wt.scala 234:50:@2772.4]
  wire  _T_267; // @[NV_NVDLA_CDMA_wt.scala 235:51:@2773.4]
  wire  _T_268; // @[NV_NVDLA_CDMA_wt.scala 235:28:@2774.4]
  wire [59:0] _GEN_21; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  wire [3:0] _GEN_23; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  wire  _GEN_24; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  wire  _GEN_25; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  wire  _T_269; // @[NV_NVDLA_CDMA_wt.scala 244:48:@2782.4]
  reg [58:0] _T_275; // @[NV_NVDLA_CDMA_wt.scala 247:33:@2785.4]
  reg [63:0] _RAND_28;
  reg [3:0] _T_278; // @[NV_NVDLA_CDMA_wt.scala 248:33:@2786.4]
  reg [31:0] _RAND_29;
  reg [2:0] _T_281; // @[NV_NVDLA_CDMA_wt.scala 249:37:@2787.4]
  reg [31:0] _RAND_30;
  wire  _T_285; // @[NV_NVDLA_CDMA_wt.scala 253:39:@2789.4]
  wire  _T_286; // @[NV_NVDLA_CDMA_wt.scala 260:39:@2795.6]
  wire [58:0] _GEN_26; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  wire [3:0] _GEN_27; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  wire [2:0] _GEN_28; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  wire  _GEN_29; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  wire [14:0] _T_337; // @[Cat.scala 30:58:@2868.4]
  wire [63:0] _T_335; // @[Cat.scala 30:58:@2866.4]
  wire  _T_333; // @[NV_NVDLA_CDMA_wt.scala 337:38:@2864.4]
  reg [3:0] _T_342; // @[NV_NVDLA_CDMA_wt.scala 345:72:@2871.4]
  reg [31:0] _RAND_31;
  wire  _T_344; // @[NV_NVDLA_CDMA_wt.scala 348:44:@2873.6]
  wire [4:0] _T_347; // @[NV_NVDLA_CDMA_wt.scala 352:72:@2878.8]
  wire [3:0] _T_348; // @[NV_NVDLA_CDMA_wt.scala 352:72:@2879.8]
  wire [3:0] _GEN_30; // @[NV_NVDLA_CDMA_wt.scala 348:76:@2874.6]
  reg [16:0] _T_357; // @[NV_NVDLA_CDMA_wt.scala 359:34:@2885.4]
  reg [31:0] _RAND_32;
  wire [14:0] _T_385; // @[Cat.scala 30:58:@2924.4]
  wire [16:0] _GEN_68; // @[NV_NVDLA_CDMA_wt.scala 387:40:@2925.4]
  wire  _T_386; // @[NV_NVDLA_CDMA_wt.scala 387:40:@2925.4]
  wire  _T_411; // @[NV_NVDLA_CDMA_wt.scala 421:40:@2957.4]
  wire [1:0] _T_401; // @[NV_NVDLA_CDMA_wt.scala 416:40:@2947.4]
  wire  _T_412; // @[NV_NVDLA_CDMA_wt.scala 421:72:@2958.4]
  wire  _T_413; // @[NV_NVDLA_CDMA_wt.scala 421:57:@2959.4]
  wire [3:0] _GEN_31; // @[NV_NVDLA_CDMA_wt.scala 347:31:@2872.4]
  reg  _T_351; // @[NV_NVDLA_CDMA_wt.scala 357:61:@2883.4]
  reg [31:0] _RAND_33;
  reg [14:0] _T_354; // @[NV_NVDLA_CDMA_wt.scala 358:64:@2884.4]
  reg [31:0] _RAND_34;
  wire  _T_359; // @[NV_NVDLA_CDMA_wt.scala 360:30:@2886.4]
  wire  _T_360; // @[NV_NVDLA_CDMA_wt.scala 360:27:@2887.4]
  wire [17:0] _T_364; // @[NV_NVDLA_CDMA_wt.scala 366:52:@2891.8]
  wire [16:0] _T_365; // @[NV_NVDLA_CDMA_wt.scala 366:52:@2892.8]
  wire [16:0] _GEN_32; // @[NV_NVDLA_CDMA_wt.scala 365:76:@2890.6]
  wire  _T_366; // @[NV_NVDLA_CDMA_wt.scala 370:32:@2897.6]
  wire [16:0] _GEN_69; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2903.10]
  wire [17:0] _T_372; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2903.10]
  wire [17:0] _T_373; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2904.10]
  wire [16:0] _T_374; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2905.10]
  wire [17:0] _T_375; // @[NV_NVDLA_CDMA_wt.scala 379:52:@2909.10]
  wire [17:0] _T_376; // @[NV_NVDLA_CDMA_wt.scala 379:52:@2910.10]
  wire [16:0] _T_377; // @[NV_NVDLA_CDMA_wt.scala 379:52:@2911.10]
  wire [16:0] _GEN_33; // @[NV_NVDLA_CDMA_wt.scala 375:76:@2900.8]
  wire  _T_379; // @[NV_NVDLA_CDMA_wt.scala 383:15:@2916.8]
  wire  _T_380; // @[NV_NVDLA_CDMA_wt.scala 383:33:@2917.8]
  wire [16:0] _GEN_34; // @[NV_NVDLA_CDMA_wt.scala 383:46:@2918.8]
  wire [16:0] _GEN_35; // @[NV_NVDLA_CDMA_wt.scala 370:45:@2898.6]
  wire [16:0] _GEN_36; // @[NV_NVDLA_CDMA_wt.scala 360:43:@2888.4]
  reg [3:0] _T_397; // @[NV_NVDLA_CDMA_wt.scala 411:35:@2943.4]
  reg [31:0] _RAND_35;
  wire [255:0] _T_398; // @[NV_NVDLA_CDMA_wt.scala 413:40:@2944.4]
  wire  _T_399; // @[NV_NVDLA_CDMA_wt.scala 414:40:@2945.4]
  wire [3:0] _T_400; // @[NV_NVDLA_CDMA_wt.scala 415:41:@2946.4]
  wire [3:0] _GEN_72; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2949.4]
  wire [4:0] _T_403; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2949.4]
  wire [3:0] _T_404; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2950.4]
  wire  _T_405; // @[NV_NVDLA_CDMA_wt.scala 419:55:@2951.4]
  wire [3:0] _T_407; // @[NV_NVDLA_CDMA_wt.scala 419:33:@2952.4]
  wire  _T_410; // @[NV_NVDLA_CDMA_wt.scala 420:60:@2955.4]
  wire [3:0] _GEN_37; // @[NV_NVDLA_CDMA_wt.scala 425:42:@2961.4]
  reg [16:0] _T_422; // @[NV_NVDLA_CDMA_wt.scala 434:33:@2966.4]
  reg [31:0] _RAND_36;
  wire [17:0] _T_437; // @[NV_NVDLA_CDMA_wt.scala 477:45:@2978.4]
  wire [16:0] _T_438; // @[NV_NVDLA_CDMA_wt.scala 477:45:@2979.4]
  wire  _T_440; // @[NV_NVDLA_CDMA_wt.scala 478:59:@2980.4]
  wire  _T_441; // @[NV_NVDLA_CDMA_wt.scala 478:42:@2981.4]
  wire  _T_442; // @[NV_NVDLA_CDMA_wt.scala 478:40:@2982.4]
  wire [16:0] _T_444; // @[Cat.scala 30:58:@2983.4]
  wire  _T_445; // @[NV_NVDLA_CDMA_wt.scala 480:51:@2984.4]
  wire  _T_446; // @[NV_NVDLA_CDMA_wt.scala 481:42:@2985.4]
  wire  _T_447; // @[NV_NVDLA_CDMA_wt.scala 481:63:@2986.4]
  wire [15:0] _T_449; // @[Cat.scala 30:58:@2987.4]
  wire [16:0] _T_451; // @[NV_NVDLA_CDMA_wt.scala 481:31:@2989.4]
  wire  _T_452; // @[NV_NVDLA_CDMA_wt.scala 490:29:@2996.4]
  wire  _T_453; // @[NV_NVDLA_CDMA_wt.scala 490:41:@2997.4]
  wire [16:0] _GEN_40; // @[NV_NVDLA_CDMA_wt.scala 490:60:@2998.4]
  reg [17:0] _T_456; // @[NV_NVDLA_CDMA_wt.scala 500:68:@3001.4]
  reg [31:0] _RAND_37;
  wire [18:0] _T_458; // @[NV_NVDLA_CDMA_wt.scala 501:49:@3002.4]
  wire [17:0] _T_459; // @[NV_NVDLA_CDMA_wt.scala 501:49:@3003.4]
  wire  _T_460; // @[NV_NVDLA_CDMA_wt.scala 502:49:@3004.4]
  wire  _T_461; // @[NV_NVDLA_CDMA_wt.scala 502:31:@3005.4]
  wire [17:0] _GEN_41; // @[NV_NVDLA_CDMA_wt.scala 506:30:@3008.4]
  wire  _T_463; // @[NV_NVDLA_CDMA_wt.scala 510:48:@3011.4]
  reg [1:0] _T_468; // @[NV_NVDLA_CDMA_wt.scala 513:77:@3013.4]
  reg [31:0] _RAND_38;
  wire [15:0] _T_471; // @[NV_NVDLA_CDMA_wt.scala 518:70:@3015.4]
  wire [15:0] _T_473; // @[NV_NVDLA_CDMA_wt.scala 519:118:@3016.4]
  wire [16:0] _T_474; // @[NV_NVDLA_CDMA_wt.scala 519:99:@3017.4]
  wire [15:0] _T_475; // @[NV_NVDLA_CDMA_wt.scala 519:99:@3018.4]
  wire [15:0] _T_476; // @[NV_NVDLA_CDMA_wt.scala 518:37:@3019.4]
  wire  _T_477; // @[NV_NVDLA_CDMA_wt.scala 520:73:@3021.4]
  wire  _T_478; // @[NV_NVDLA_CDMA_wt.scala 520:129:@3022.4]
  wire  _T_479; // @[NV_NVDLA_CDMA_wt.scala 520:40:@3023.4]
  wire [1:0] _GEN_73; // @[NV_NVDLA_CDMA_wt.scala 522:118:@3026.6]
  wire  _T_481; // @[NV_NVDLA_CDMA_wt.scala 522:118:@3026.6]
  wire [1:0] _T_492; // @[NV_NVDLA_CDMA_wt.scala 522:150:@3031.6]
  wire [1:0] _GEN_42; // @[NV_NVDLA_CDMA_wt.scala 521:34:@3025.4]
  wire [255:0] _T_494; // @[NV_NVDLA_CDMA_wt.scala 531:36:@3035.4]
  reg  _T_497; // @[NV_NVDLA_CDMA_wt.scala 532:76:@3036.4]
  reg [31:0] _RAND_39;
  reg [16:0] _T_500; // @[Reg.scala 19:20:@3039.4]
  reg [31:0] _RAND_40;
  wire [16:0] _T_465; // @[NV_NVDLA_CDMA_wt.scala 511:37:@3012.4 NV_NVDLA_CDMA_wt.scala 518:31:@3020.4]
  wire [16:0] _GEN_43; // @[Reg.scala 20:19:@3040.4]
  reg [255:0] _T_503; // @[Reg.scala 19:20:@3044.4]
  reg [255:0] _RAND_41;
  wire [255:0] _GEN_44; // @[Reg.scala 20:19:@3045.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CDMA_wt.scala 548:35:@3052.4]
  wire  _T_514; // @[NV_NVDLA_CDMA_wt.scala 556:50:@3059.4]
  wire  _T_515; // @[NV_NVDLA_CDMA_wt.scala 556:74:@3060.4]
  wire  _T_516; // @[NV_NVDLA_CDMA_wt.scala 556:72:@3061.4]
  wire [3:0] _T_518; // @[NV_NVDLA_CDMA_wt.scala 556:32:@3062.4]
  wire [2:0] _T_521; // @[NV_NVDLA_CDMA_wt.scala 557:32:@3063.4]
  reg [25:0] _T_560; // @[NV_NVDLA_CDMA_wt.scala 591:33:@3102.4]
  reg [31:0] _RAND_42;
  reg [25:0] _T_615; // @[NV_NVDLA_CDMA_wt.scala 642:37:@3150.4]
  reg [31:0] _RAND_43;
  wire [26:0] _T_624; // @[NV_NVDLA_CDMA_wt.scala 647:39:@3154.4]
  wire [26:0] _T_625; // @[NV_NVDLA_CDMA_wt.scala 647:39:@3155.4]
  wire [25:0] _T_626; // @[NV_NVDLA_CDMA_wt.scala 647:39:@3156.4]
  wire [14:0] _T_627; // @[NV_NVDLA_CDMA_wt.scala 652:41:@3157.4]
  wire [15:0] _T_523; // @[Cat.scala 30:58:@3064.4]
  reg  _T_563; // @[NV_NVDLA_CDMA_wt.scala 592:33:@3103.4]
  reg [31:0] _RAND_44;
  wire  _T_605; // @[NV_NVDLA_CDMA_wt.scala 622:26:@3136.4]
  wire [33:0] _T_597; // @[Cat.scala 30:58:@3129.4]
  reg [31:0] _T_566; // @[NV_NVDLA_CDMA_wt.scala 593:36:@3104.4]
  reg [31:0] _RAND_45;
  wire [33:0] _GEN_75; // @[NV_NVDLA_CDMA_wt.scala 618:95:@3130.4]
  wire  _T_598; // @[NV_NVDLA_CDMA_wt.scala 618:95:@3130.4]
  wire  _T_599; // @[NV_NVDLA_CDMA_wt.scala 618:35:@3131.4]
  wire [1:0] _T_600; // @[NV_NVDLA_CDMA_wt.scala 619:40:@3132.4]
  wire  _T_602; // @[NV_NVDLA_CDMA_wt.scala 619:70:@3133.4]
  wire  _T_603; // @[NV_NVDLA_CDMA_wt.scala 619:24:@3134.4]
  wire  _T_604; // @[NV_NVDLA_CDMA_wt.scala 618:117:@3135.4]
  wire  _T_607; // @[NV_NVDLA_CDMA_wt.scala 622:25:@3137.4]
  wire [16:0] _T_525; // @[NV_NVDLA_CDMA_wt.scala 563:34:@3065.4]
  wire [15:0] _T_527; // @[Cat.scala 30:58:@3067.4]
  wire [16:0] _T_529; // @[NV_NVDLA_CDMA_wt.scala 564:31:@3068.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3070.4]
  wire [14:0] _T_530; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3070.4]
  wire [13:0] _T_531; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3071.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3072.4]
  wire [14:0] _T_532; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3072.4]
  wire [14:0] _T_533; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3073.4]
  wire [13:0] _T_534; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3074.4]
  wire [16:0] _GEN_78; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3075.4]
  wire [17:0] _T_535; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3075.4]
  wire [16:0] _T_536; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3076.4]
  wire [17:0] _T_537; // @[NV_NVDLA_CDMA_wt.scala 572:63:@3077.4]
  wire [17:0] _T_538; // @[NV_NVDLA_CDMA_wt.scala 572:63:@3078.4]
  wire [16:0] _T_539; // @[NV_NVDLA_CDMA_wt.scala 572:63:@3079.4]
  wire [17:0] _T_541; // @[NV_NVDLA_CDMA_wt.scala 573:57:@3080.4]
  wire [16:0] _T_542; // @[NV_NVDLA_CDMA_wt.scala 573:57:@3081.4]
  wire [17:0] _T_543; // @[NV_NVDLA_CDMA_wt.scala 573:78:@3082.4]
  wire [17:0] _T_544; // @[NV_NVDLA_CDMA_wt.scala 573:78:@3083.4]
  wire [16:0] _T_545; // @[NV_NVDLA_CDMA_wt.scala 573:78:@3084.4]
  wire [16:0] _T_546; // @[NV_NVDLA_CDMA_wt.scala 573:28:@3085.4]
  wire  _T_548; // @[NV_NVDLA_CDMA_wt.scala 574:74:@3087.4]
  wire [13:0] _GEN_46; // @[NV_NVDLA_CDMA_wt.scala 576:31:@3088.4]
  wire  _T_549; // @[NV_NVDLA_CDMA_wt.scala 579:27:@3091.4]
  wire [16:0] _GEN_47; // @[NV_NVDLA_CDMA_wt.scala 579:43:@3092.4]
  wire  _T_550; // @[NV_NVDLA_CDMA_wt.scala 582:24:@3095.4]
  wire  _T_551; // @[NV_NVDLA_CDMA_wt.scala 582:37:@3096.4]
  wire [16:0] _GEN_48; // @[NV_NVDLA_CDMA_wt.scala 582:49:@3097.4]
  reg [11:0] _T_554; // @[NV_NVDLA_CDMA_wt.scala 589:35:@3100.4]
  reg [31:0] _RAND_46;
  reg [31:0] _T_557; // @[NV_NVDLA_CDMA_wt.scala 590:40:@3101.4]
  reg [31:0] _RAND_47;
  wire [12:0] _T_568; // @[NV_NVDLA_CDMA_wt.scala 595:49:@3105.4]
  wire [11:0] _T_569; // @[NV_NVDLA_CDMA_wt.scala 595:49:@3106.4]
  wire  _T_570; // @[NV_NVDLA_CDMA_wt.scala 596:51:@3107.4]
  wire [11:0] _T_572; // @[NV_NVDLA_CDMA_wt.scala 597:33:@3108.4]
  wire  _T_575; // @[NV_NVDLA_CDMA_wt.scala 599:28:@3109.4]
  wire  _T_576; // @[NV_NVDLA_CDMA_wt.scala 598:28:@3110.4]
  wire [24:0] _T_578; // @[Cat.scala 30:58:@3111.4]
  wire [31:0] _GEN_79; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3112.4]
  wire [32:0] _T_580; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3112.4]
  wire [31:0] _T_581; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3113.4]
  wire [31:0] _T_582; // @[NV_NVDLA_CDMA_wt.scala 603:34:@3114.4]
  wire [31:0] _T_583; // @[NV_NVDLA_CDMA_wt.scala 602:34:@3115.4]
  wire  _T_584; // @[NV_NVDLA_CDMA_wt.scala 605:41:@3116.4]
  wire  _T_585; // @[NV_NVDLA_CDMA_wt.scala 605:39:@3117.4]
  wire  _T_587; // @[NV_NVDLA_CDMA_wt.scala 606:42:@3119.4]
  wire [31:0] _T_589; // @[NV_NVDLA_CDMA_wt.scala 607:38:@3120.4]
  wire  _T_590; // @[NV_NVDLA_CDMA_wt.scala 611:19:@3122.4]
  wire [31:0] _GEN_49; // @[NV_NVDLA_CDMA_wt.scala 611:36:@3123.4]
  wire [26:0] _T_592; // @[NV_NVDLA_CDMA_wt.scala 615:45:@3126.4]
  wire [25:0] _T_593; // @[NV_NVDLA_CDMA_wt.scala 615:45:@3127.4]
  wire [25:0] _T_595; // @[NV_NVDLA_CDMA_wt.scala 616:31:@3128.4]
  wire  _T_608; // @[NV_NVDLA_CDMA_wt.scala 624:19:@3139.4]
  wire [11:0] _GEN_50; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  wire  _GEN_51; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  wire [31:0] _GEN_52; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  wire  _T_609; // @[NV_NVDLA_CDMA_wt.scala 629:19:@3145.4]
  wire [25:0] _GEN_53; // @[NV_NVDLA_CDMA_wt.scala 629:38:@3146.4]
  reg  _T_612; // @[NV_NVDLA_CDMA_wt.scala 641:31:@3149.4]
  reg [31:0] _RAND_48;
  reg [14:0] _T_618; // @[NV_NVDLA_CDMA_wt.scala 643:34:@3151.4]
  reg [31:0] _RAND_49;
  reg [5:0] _T_621; // @[NV_NVDLA_CDMA_wt.scala 644:34:@3152.4]
  reg [31:0] _RAND_50;
  wire [25:0] _T_623; // @[NV_NVDLA_CDMA_wt.scala 646:35:@3153.4]
  wire  _T_628; // @[NV_NVDLA_CDMA_wt.scala 655:33:@3159.4]
  wire [5:0] _T_630; // @[NV_NVDLA_CDMA_wt.scala 656:52:@3160.4]
  wire [6:0] _T_632; // @[NV_NVDLA_CDMA_wt.scala 656:71:@3161.4]
  wire [6:0] _T_633; // @[NV_NVDLA_CDMA_wt.scala 655:32:@3162.4]
  wire [25:0] _GEN_54; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  wire [14:0] _GEN_55; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  wire [6:0] _GEN_56; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  reg  _T_638; // @[NV_NVDLA_CDMA_wt.scala 666:69:@3170.4]
  reg [31:0] _RAND_51;
  reg  _T_641; // @[NV_NVDLA_CDMA_wt.scala 666:69:@3171.4]
  reg [31:0] _RAND_52;
  reg  _T_644; // @[NV_NVDLA_CDMA_wt.scala 666:69:@3172.4]
  reg [31:0] _RAND_53;
  reg [5:0] _T_649; // @[NV_NVDLA_CDMA_wt.scala 668:72:@3174.4]
  reg [31:0] _RAND_54;
  reg [5:0] _T_652; // @[NV_NVDLA_CDMA_wt.scala 668:72:@3175.4]
  reg [31:0] _RAND_55;
  reg [5:0] _T_655; // @[NV_NVDLA_CDMA_wt.scala 668:72:@3176.4]
  reg [31:0] _RAND_56;
  reg [14:0] _T_660; // @[NV_NVDLA_CDMA_wt.scala 670:72:@3178.4]
  reg [31:0] _RAND_57;
  reg [14:0] _T_663; // @[NV_NVDLA_CDMA_wt.scala 670:72:@3179.4]
  reg [31:0] _RAND_58;
  reg [14:0] _T_666; // @[NV_NVDLA_CDMA_wt.scala 670:72:@3180.4]
  reg [31:0] _RAND_59;
  wire [14:0] _GEN_57; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3185.4]
  wire [5:0] _GEN_58; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3185.4]
  wire [14:0] _GEN_59; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3190.4]
  wire [5:0] _GEN_60; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3190.4]
  wire [14:0] _GEN_61; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3195.4]
  wire [5:0] _GEN_62; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3195.4]
  wire  _T_667; // @[NV_NVDLA_CDMA_wt.scala 692:52:@3202.4]
  wire  _T_668; // @[NV_NVDLA_CDMA_wt.scala 692:50:@3203.4]
  wire  _T_669; // @[NV_NVDLA_CDMA_wt.scala 692:68:@3204.4]
  reg  _T_672; // @[NV_NVDLA_CDMA_wt.scala 692:34:@3205.4]
  reg [31:0] _RAND_60;
  wire  _T_673; // @[NV_NVDLA_CDMA_wt.scala 693:60:@3207.4]
  reg  _T_676; // @[NV_NVDLA_CDMA_wt.scala 693:34:@3208.4]
  reg [31:0] _RAND_61;
  wire  _T_677; // @[NV_NVDLA_CDMA_wt.scala 694:51:@3210.4]
  reg  _T_680; // @[NV_NVDLA_CDMA_wt.scala 694:34:@3211.4]
  reg [31:0] _RAND_62;
  reg  _T_687; // @[NV_NVDLA_CDMA_wt.scala 707:36:@3225.4]
  reg [31:0] _RAND_63;
  wire  _T_688; // @[NV_NVDLA_CDMA_wt.scala 708:56:@3227.4]
  reg  _T_691; // @[NV_NVDLA_CDMA_wt.scala 708:36:@3228.4]
  reg [31:0] _RAND_64;
  reg  _T_694; // @[NV_NVDLA_CDMA_wt.scala 709:36:@3230.4]
  reg [31:0] _RAND_65;
  reg  _T_698; // @[NV_NVDLA_CDMA_wt.scala 710:36:@3233.4]
  reg [31:0] _RAND_66;
  wire [8:0] _T_700; // @[NV_NVDLA_CDMA_wt.scala 712:41:@3235.4 NV_NVDLA_CDMA_wt.scala 722:31:@3248.4]
  wire  _T_702; // @[NV_NVDLA_CDMA_wt.scala 713:48:@3236.4]
  NV_soDLA_DMAIF_rdreq NV_soDLA_DMAIF_rdreq ( // @[NV_NVDLA_CDMA_wt.scala 299:41:@2828.4]
    .reset(NV_NVDLA_DMAIF_rdreq_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk),
    .io_dmaif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready),
    .io_dmaif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid),
    .io_dmaif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits),
    .io_mcif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready),
    .io_mcif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid),
    .io_mcif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits),
    .io_cvif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready),
    .io_cvif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid),
    .io_cvif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits),
    .io_reg2dp_src_ram_type(NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type)
  );
  NV_soDLA_DMAIF_rdrsp NV_soDLA_DMAIF_rdrsp ( // @[NV_NVDLA_CDMA_wt.scala 311:41:@2842.4]
    .reset(NV_NVDLA_DMAIF_rdrsp_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk),
    .io_mcif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready),
    .io_mcif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid),
    .io_mcif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits),
    .io_cvif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready),
    .io_cvif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid),
    .io_cvif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits),
    .io_dmaif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready),
    .io_dmaif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid),
    .io_dmaif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits)
  );
  NV_NVDLA_fifo NV_NVDLA_fifo ( // @[NV_NVDLA_CDMA_wt.scala 323:30:@2853.4]
    .clock(NV_NVDLA_fifo_clock),
    .reset(NV_NVDLA_fifo_reset),
    .io_clk(NV_NVDLA_fifo_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_io_wr_pd),
    .io_rd_pvld(NV_NVDLA_fifo_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_io_rd_pd)
  );
  NV_NVDLA_fifo_1 NV_NVDLA_fifo_1 ( // @[NV_NVDLA_CDMA_wt.scala 392:24:@2930.4]
    .clock(NV_NVDLA_fifo_1_clock),
    .reset(NV_NVDLA_fifo_1_reset),
    .io_clk(NV_NVDLA_fifo_1_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_1_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_1_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_1_io_wr_pd),
    .io_rd_pvld(NV_NVDLA_fifo_1_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_1_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_1_io_rd_pd)
  );
  NV_COUNTER_STAGE_histogram NV_COUNTER_STAGE_histogram ( // @[NV_NVDLA_CDMA_wt.scala 698:21:@3213.4]
    .reset(NV_COUNTER_STAGE_histogram_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_io_rd_stall_inc),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_io_cnt_cur)
  );
  NV_COUNTER_STAGE_histogram_1 NV_COUNTER_STAGE_histogram_1 ( // @[NV_NVDLA_CDMA_wt.scala 716:23:@3240.4]
    .reset(NV_COUNTER_STAGE_histogram_1_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_1_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc),
    .io_rd_stall_dec(NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_1_io_cnt_cur)
  );
  assign _T_92 = 2'h0 == _T_89; // @[Conditional.scala 37:30:@2616.4]
  assign _T_135 = _T_105 != io_reg2dp_data_bank; // @[NV_NVDLA_CDMA_wt.scala 133:38:@2672.4]
  assign _T_136 = _T_112 != io_reg2dp_weight_bank; // @[NV_NVDLA_CDMA_wt.scala 133:83:@2673.4]
  assign _T_137 = _T_135 | _T_136; // @[NV_NVDLA_CDMA_wt.scala 133:63:@2674.4]
  assign _T_93 = io_reg2dp_op_en & _T_137; // @[NV_NVDLA_CDMA_wt.scala 104:31:@2618.6]
  assign _T_94 = io_reg2dp_op_en & io_reg2dp_weight_reuse; // @[NV_NVDLA_CDMA_wt.scala 105:36:@2623.8]
  assign _T_95 = _T_94 & _T_83; // @[NV_NVDLA_CDMA_wt.scala 105:61:@2624.8]
  assign _GEN_0 = io_reg2dp_op_en ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_wt.scala 106:37:@2629.10]
  assign _GEN_1 = _T_95 ? 2'h3 : _GEN_0; // @[NV_NVDLA_CDMA_wt.scala 105:85:@2625.8]
  assign _GEN_2 = _T_93 ? 2'h1 : _GEN_1; // @[NV_NVDLA_CDMA_wt.scala 104:47:@2619.6]
  assign _T_96 = 2'h1 == _T_89; // @[Conditional.scala 37:30:@2634.6]
  assign _T_157 = ~ _T_144; // @[NV_NVDLA_CDMA_wt.scala 153:41:@2692.4]
  assign _T_158 = _T_147 & _T_157; // @[NV_NVDLA_CDMA_wt.scala 153:39:@2693.4]
  assign _GEN_3 = _T_158 ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_wt.scala 109:32:@2636.8]
  assign _T_97 = 2'h2 == _T_89; // @[Conditional.scala 37:30:@2641.8]
  assign _T_133 = _T_122 == 4'h8; // @[NV_NVDLA_CDMA_wt.scala 132:50:@2669.4]
  assign _T_134 = _T_119 & _T_133; // @[NV_NVDLA_CDMA_wt.scala 132:31:@2670.4]
  assign _GEN_4 = _T_134 ? 2'h3 : 2'h0; // @[NV_NVDLA_CDMA_wt.scala 112:27:@2643.10]
  assign _GEN_7 = _T_97 ? _GEN_4 : 2'h0; // @[Conditional.scala 39:67:@2642.8]
  assign _GEN_8 = _T_96 ? _GEN_3 : _GEN_7; // @[Conditional.scala 39:67:@2635.6]
  assign _GEN_9 = _T_92 ? _GEN_2 : _GEN_8; // @[Conditional.scala 40:58:@2617.4]
  assign _T_125 = _T_122 != 4'h8; // @[NV_NVDLA_CDMA_wt.scala 130:64:@2663.4]
  assign _T_126 = _T_119 & _T_125; // @[NV_NVDLA_CDMA_wt.scala 130:45:@2664.4]
  assign _T_128 = _T_122 + 4'h1; // @[NV_NVDLA_CDMA_wt.scala 130:103:@2665.4]
  assign _T_129 = _T_122 + 4'h1; // @[NV_NVDLA_CDMA_wt.scala 130:103:@2666.4]
  assign _T_130 = _T_126 ? _T_129 : _T_122; // @[NV_NVDLA_CDMA_wt.scala 130:32:@2667.4]
  assign _T_151 = _T_89 == 2'h0; // @[NV_NVDLA_CDMA_wt.scala 146:47:@2684.4]
  assign _T_152 = io_reg2dp_op_en & _T_151; // @[NV_NVDLA_CDMA_wt.scala 146:33:@2685.4]
  assign _T_131 = _T_152 ? 4'h0 : _T_130; // @[NV_NVDLA_CDMA_wt.scala 129:32:@2668.4]
  assign _T_153 = _T_89 == 2'h2; // @[NV_NVDLA_CDMA_wt.scala 148:30:@2687.4]
  assign _T_138 = _T_152 | _T_153; // @[NV_NVDLA_CDMA_wt.scala 135:19:@2676.4]
  assign _GEN_10 = _T_138 ? _T_131 : _T_122; // @[NV_NVDLA_CDMA_wt.scala 135:32:@2677.4]
  assign _T_154 = _T_89 == 2'h1; // @[NV_NVDLA_CDMA_wt.scala 149:33:@2689.4]
  assign _T_155 = _T_150 & _T_144; // @[NV_NVDLA_CDMA_wt.scala 150:33:@2690.4]
  assign _T_156 = _GEN_9 == 2'h2; // @[NV_NVDLA_CDMA_wt.scala 151:37:@2691.4]
  assign _GEN_11 = io_status2dma_fsm_switch ? io_reg2dp_data_bank : _T_105; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  assign _GEN_12 = io_status2dma_fsm_switch ? io_reg2dp_weight_bank : _T_112; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  assign _GEN_13 = io_status2dma_fsm_switch ? io_reg2dp_skip_weight_rls : _T_83; // @[NV_NVDLA_CDMA_wt.scala 166:20:@2701.4]
  assign _T_187 = io_reg2dp_byte_per_kernel + 18'h1; // @[NV_NVDLA_CDMA_wt.scala 181:63:@2715.4]
  assign _T_192 = io_reg2dp_weight_kernel[12:6]; // @[NV_NVDLA_CDMA_wt.scala 184:43:@2720.4]
  assign _T_194 = _T_192 + 7'h1; // @[NV_NVDLA_CDMA_wt.scala 185:28:@2721.4]
  assign _T_196 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CDMA_wt.scala 186:43:@2722.4]
  assign _T_198 = io_reg2dp_weight_bank + 5'h1; // @[NV_NVDLA_CDMA_wt.scala 187:47:@2723.4]
  assign _T_199 = _T_198 + _T_196; // @[NV_NVDLA_CDMA_wt.scala 188:43:@2724.4]
  assign _GEN_15 = _T_152 ? {{4'd0}, _T_194} : _T_168; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  assign _GEN_16 = _T_152 ? _T_198 : _T_175; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  assign _GEN_17 = _T_152 ? _T_199 : _T_182; // @[NV_NVDLA_CDMA_wt.scala 192:19:@2728.4]
  assign _GEN_63 = {{25'd0}, _T_209}; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2738.4]
  assign _T_218 = _T_212 - _GEN_63; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2738.4]
  assign _T_219 = $unsigned(_T_218); // @[NV_NVDLA_CDMA_wt.scala 211:52:@2739.4]
  assign _T_220 = _T_219[28:0]; // @[NV_NVDLA_CDMA_wt.scala 211:52:@2740.4]
  assign _T_221 = io_reg2dp_weight_bytes[31:5]; // @[NV_NVDLA_CDMA_wt.scala 212:66:@2741.4]
  assign _T_222 = _T_152 ? {{2'd0}, _T_221} : _T_220; // @[NV_NVDLA_CDMA_wt.scala 212:33:@2742.4]
  assign _T_224 = io_reg2dp_weight_addr_low[2:0]; // @[NV_NVDLA_CDMA_wt.scala 213:92:@2743.4]
  assign _GEN_64 = {{1'd0}, _T_224}; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2744.4]
  assign _T_225 = 4'h8 - _GEN_64; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2744.4]
  assign _T_226 = $unsigned(_T_225); // @[NV_NVDLA_CDMA_wt.scala 213:65:@2745.4]
  assign _T_227 = _T_226[3:0]; // @[NV_NVDLA_CDMA_wt.scala 213:65:@2746.4]
  assign _T_229 = _T_152 ? _T_227 : 4'h8; // @[NV_NVDLA_CDMA_wt.scala 213:37:@2747.4]
  assign _GEN_65 = {{25'd0}, _T_229}; // @[NV_NVDLA_CDMA_wt.scala 214:52:@2748.4]
  assign _T_230 = _GEN_65 > _T_222; // @[NV_NVDLA_CDMA_wt.scala 214:52:@2748.4]
  assign _T_231 = _T_222[3:0]; // @[NV_NVDLA_CDMA_wt.scala 214:92:@2749.4]
  assign _T_232 = _T_230 ? _T_231 : _T_229; // @[NV_NVDLA_CDMA_wt.scala 214:28:@2750.4]
  assign _T_308 = ~ _T_272; // @[NV_NVDLA_CDMA_wt.scala 275:48:@2810.4]
  assign _T_313 = NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 277:30:@2815.4 NV_NVDLA_CDMA_wt.scala 309:20:@2841.4]
  assign _T_315 = NV_NVDLA_fifo_1_io_wr_prdy; // @[NV_NVDLA_CDMA_wt.scala 278:34:@2816.4 NV_NVDLA_CDMA_wt.scala 399:24:@2936.4]
  assign _T_316 = _T_313 & _T_315; // @[NV_NVDLA_CDMA_wt.scala 279:41:@2817.4]
  assign _GEN_66 = {{3'd0}, _T_289}; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2801.4]
  assign _T_296 = _GEN_66 + _T_292; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2801.4]
  assign _T_297 = _GEN_66 + _T_292; // @[NV_NVDLA_CDMA_wt.scala 269:36:@2802.4]
  assign _T_298 = _T_297 + _T_295; // @[NV_NVDLA_CDMA_wt.scala 269:53:@2803.4]
  assign _T_299 = _T_297 + _T_295; // @[NV_NVDLA_CDMA_wt.scala 269:53:@2804.4]
  assign _T_301 = {_T_175,10'h0}; // @[Cat.scala 30:58:@2805.4]
  assign _T_303 = _T_301 + 16'h4; // @[NV_NVDLA_CDMA_wt.scala 270:115:@2806.4]
  assign _T_304 = _T_299 > _T_303; // @[NV_NVDLA_CDMA_wt.scala 270:53:@2807.4]
  assign _T_305 = _T_153 & _T_304; // @[NV_NVDLA_CDMA_wt.scala 270:38:@2808.4]
  assign _T_317 = ~ _T_305; // @[NV_NVDLA_CDMA_wt.scala 280:42:@2818.4]
  assign _T_318 = _T_272 & _T_317; // @[NV_NVDLA_CDMA_wt.scala 280:40:@2819.4]
  assign _T_319 = ~ _T_284; // @[NV_NVDLA_CDMA_wt.scala 280:64:@2820.4]
  assign _T_320 = _T_318 & _T_319; // @[NV_NVDLA_CDMA_wt.scala 280:62:@2821.4]
  assign _T_321 = _T_316 & _T_320; // @[NV_NVDLA_CDMA_wt.scala 281:34:@2822.4]
  assign _T_309 = _T_308 | _T_321; // @[NV_NVDLA_CDMA_wt.scala 275:63:@2811.4]
  assign _T_310 = _T_153 & _T_309; // @[NV_NVDLA_CDMA_wt.scala 275:45:@2812.4]
  assign _T_311 = _T_152 | _T_310; // @[NV_NVDLA_CDMA_wt.scala 275:31:@2813.4]
  assign _GEN_19 = _T_311 ? _T_232 : _T_209; // @[NV_NVDLA_CDMA_wt.scala 216:27:@2751.4]
  assign _GEN_20 = _T_311 ? _T_222 : _T_212; // @[NV_NVDLA_CDMA_wt.scala 216:27:@2751.4]
  assign _T_251 = _T_212 == _GEN_63; // @[NV_NVDLA_CDMA_wt.scala 231:69:@2762.4]
  assign _T_252 = _T_215 & _T_251; // @[NV_NVDLA_CDMA_wt.scala 231:45:@2763.4]
  assign _T_253 = _T_235[58:3]; // @[NV_NVDLA_CDMA_wt.scala 232:41:@2764.4]
  assign _T_255 = _T_253 + 56'h1; // @[NV_NVDLA_CDMA_wt.scala 232:61:@2765.4]
  assign _T_256 = ~ _T_250; // @[NV_NVDLA_CDMA_wt.scala 233:29:@2766.4]
  assign _T_257 = {io_reg2dp_weight_addr_high,io_reg2dp_weight_addr_low}; // @[Cat.scala 30:58:@2767.4]
  assign _T_259 = {_T_255,3'h0}; // @[Cat.scala 30:58:@2768.4]
  assign _T_260 = _T_256 ? {{1'd0}, _T_257} : _T_259; // @[NV_NVDLA_CDMA_wt.scala 233:28:@2769.4]
  assign _T_261 = _T_209[2:0]; // @[NV_NVDLA_CDMA_wt.scala 234:43:@2770.4]
  assign _T_263 = _T_261 - 3'h1; // @[NV_NVDLA_CDMA_wt.scala 234:50:@2771.4]
  assign _T_264 = $unsigned(_T_263); // @[NV_NVDLA_CDMA_wt.scala 234:50:@2772.4]
  assign _T_267 = _T_244 ? 1'h1 : _T_247; // @[NV_NVDLA_CDMA_wt.scala 235:51:@2773.4]
  assign _T_268 = _T_152 ? 1'h0 : _T_267; // @[NV_NVDLA_CDMA_wt.scala 235:28:@2774.4]
  assign _GEN_21 = _T_311 ? _T_260 : {{1'd0}, _T_235}; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  assign _GEN_22 = _T_311 ? _T_209 : _T_238; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  assign _GEN_23 = _T_311 ? _T_264 : {{1'd0}, _T_241}; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  assign _GEN_24 = _T_311 ? _T_252 : _T_244; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  assign _GEN_25 = _T_311 ? _T_268 : _T_247; // @[NV_NVDLA_CDMA_wt.scala 237:27:@2775.4]
  assign _T_269 = _T_215 & _T_156; // @[NV_NVDLA_CDMA_wt.scala 244:48:@2782.4]
  assign _T_285 = _T_156 & _T_250; // @[NV_NVDLA_CDMA_wt.scala 253:39:@2789.4]
  assign _T_286 = _T_153 & _T_247; // @[NV_NVDLA_CDMA_wt.scala 260:39:@2795.6]
  assign _GEN_26 = _T_311 ? _T_235 : _T_275; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  assign _GEN_27 = _T_311 ? _T_238 : _T_278; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  assign _GEN_28 = _T_311 ? _T_241 : _T_281; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  assign _GEN_29 = _T_311 ? _T_286 : _T_284; // @[NV_NVDLA_CDMA_wt.scala 256:28:@2791.4]
  assign _T_337 = {12'h0,_T_281}; // @[Cat.scala 30:58:@2868.4]
  assign _T_335 = {_T_275,5'h0}; // @[Cat.scala 30:58:@2866.4]
  assign _T_333 = _T_320 & _T_315; // @[NV_NVDLA_CDMA_wt.scala 337:38:@2864.4]
  assign _T_344 = _T_342 == 4'h1; // @[NV_NVDLA_CDMA_wt.scala 348:44:@2873.6]
  assign _T_347 = _T_342 + 4'h1; // @[NV_NVDLA_CDMA_wt.scala 352:72:@2878.8]
  assign _T_348 = _T_342 + 4'h1; // @[NV_NVDLA_CDMA_wt.scala 352:72:@2879.8]
  assign _GEN_30 = _T_344 ? 4'h0 : _T_348; // @[NV_NVDLA_CDMA_wt.scala 348:76:@2874.6]
  assign _T_385 = {_T_175,9'h0}; // @[Cat.scala 30:58:@2924.4]
  assign _GEN_68 = {{2'd0}, _T_385}; // @[NV_NVDLA_CDMA_wt.scala 387:40:@2925.4]
  assign _T_386 = _T_357 < _GEN_68; // @[NV_NVDLA_CDMA_wt.scala 387:40:@2925.4]
  assign _T_411 = NV_NVDLA_fifo_io_rd_pvld & _T_386; // @[NV_NVDLA_CDMA_wt.scala 421:40:@2957.4]
  assign _T_401 = NV_NVDLA_fifo_1_io_rd_pd[5:4]; // @[NV_NVDLA_CDMA_wt.scala 416:40:@2947.4]
  assign _T_412 = _T_401 == 2'h0; // @[NV_NVDLA_CDMA_wt.scala 421:72:@2958.4]
  assign _T_413 = _T_411 & _T_412; // @[NV_NVDLA_CDMA_wt.scala 421:57:@2959.4]
  assign _GEN_31 = _T_413 ? _GEN_30 : _T_342; // @[NV_NVDLA_CDMA_wt.scala 347:31:@2872.4]
  assign _T_359 = _T_351 == 1'h0; // @[NV_NVDLA_CDMA_wt.scala 360:30:@2886.4]
  assign _T_360 = _T_413 & _T_359; // @[NV_NVDLA_CDMA_wt.scala 360:27:@2887.4]
  assign _T_364 = _T_357 + 17'h1; // @[NV_NVDLA_CDMA_wt.scala 366:52:@2891.8]
  assign _T_365 = _T_357 + 17'h1; // @[NV_NVDLA_CDMA_wt.scala 366:52:@2892.8]
  assign _GEN_32 = _T_344 ? _T_365 : _T_357; // @[NV_NVDLA_CDMA_wt.scala 365:76:@2890.6]
  assign _T_366 = _T_413 & _T_351; // @[NV_NVDLA_CDMA_wt.scala 370:32:@2897.6]
  assign _GEN_69 = {{2'd0}, _T_354}; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2903.10]
  assign _T_372 = _T_365 - _GEN_69; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2903.10]
  assign _T_373 = $unsigned(_T_372); // @[NV_NVDLA_CDMA_wt.scala 376:58:@2904.10]
  assign _T_374 = _T_373[16:0]; // @[NV_NVDLA_CDMA_wt.scala 376:58:@2905.10]
  assign _T_375 = _T_357 - _GEN_69; // @[NV_NVDLA_CDMA_wt.scala 379:52:@2909.10]
  assign _T_376 = $unsigned(_T_375); // @[NV_NVDLA_CDMA_wt.scala 379:52:@2910.10]
  assign _T_377 = _T_376[16:0]; // @[NV_NVDLA_CDMA_wt.scala 379:52:@2911.10]
  assign _GEN_33 = _T_344 ? _T_374 : _T_377; // @[NV_NVDLA_CDMA_wt.scala 375:76:@2900.8]
  assign _T_379 = _T_413 == 1'h0; // @[NV_NVDLA_CDMA_wt.scala 383:15:@2916.8]
  assign _T_380 = _T_379 & _T_351; // @[NV_NVDLA_CDMA_wt.scala 383:33:@2917.8]
  assign _GEN_34 = _T_380 ? _T_377 : _T_357; // @[NV_NVDLA_CDMA_wt.scala 383:46:@2918.8]
  assign _GEN_35 = _T_366 ? _GEN_33 : _GEN_34; // @[NV_NVDLA_CDMA_wt.scala 370:45:@2898.6]
  assign _GEN_36 = _T_360 ? _GEN_32 : _GEN_35; // @[NV_NVDLA_CDMA_wt.scala 360:43:@2888.4]
  assign _T_398 = NV_NVDLA_fifo_io_rd_pd[255:0]; // @[NV_NVDLA_CDMA_wt.scala 413:40:@2944.4]
  assign _T_399 = NV_NVDLA_fifo_io_rd_pd[256]; // @[NV_NVDLA_CDMA_wt.scala 414:40:@2945.4]
  assign _T_400 = NV_NVDLA_fifo_1_io_rd_pd[3:0]; // @[NV_NVDLA_CDMA_wt.scala 415:41:@2946.4]
  assign _GEN_72 = {{3'd0}, _T_399}; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2949.4]
  assign _T_403 = _T_397 + _GEN_72; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2949.4]
  assign _T_404 = _T_397 + _GEN_72; // @[NV_NVDLA_CDMA_wt.scala 417:49:@2950.4]
  assign _T_405 = _T_404 == _T_400; // @[NV_NVDLA_CDMA_wt.scala 419:55:@2951.4]
  assign _T_407 = _T_405 ? 4'h0 : _T_404; // @[NV_NVDLA_CDMA_wt.scala 419:33:@2952.4]
  assign _T_410 = _T_411 & _T_405; // @[NV_NVDLA_CDMA_wt.scala 420:60:@2955.4]
  assign _GEN_37 = _T_411 ? _T_407 : _T_397; // @[NV_NVDLA_CDMA_wt.scala 425:42:@2961.4]
  assign _T_437 = _T_422 + 17'h1; // @[NV_NVDLA_CDMA_wt.scala 477:45:@2978.4]
  assign _T_438 = _T_422 + 17'h1; // @[NV_NVDLA_CDMA_wt.scala 477:45:@2979.4]
  assign _T_440 = _T_422 != 17'h0; // @[NV_NVDLA_CDMA_wt.scala 478:59:@2980.4]
  assign _T_441 = ~ _T_440; // @[NV_NVDLA_CDMA_wt.scala 478:42:@2981.4]
  assign _T_442 = _T_152 & _T_441; // @[NV_NVDLA_CDMA_wt.scala 478:40:@2982.4]
  assign _T_444 = {_T_182,10'h0}; // @[Cat.scala 30:58:@2983.4]
  assign _T_445 = _T_438 == _T_444; // @[NV_NVDLA_CDMA_wt.scala 480:51:@2984.4]
  assign _T_446 = _T_155 | _T_442; // @[NV_NVDLA_CDMA_wt.scala 481:42:@2985.4]
  assign _T_447 = _T_446 | _T_445; // @[NV_NVDLA_CDMA_wt.scala 481:63:@2986.4]
  assign _T_449 = {_T_196,10'h0}; // @[Cat.scala 30:58:@2987.4]
  assign _T_451 = _T_447 ? {{1'd0}, _T_449} : _T_438; // @[NV_NVDLA_CDMA_wt.scala 481:31:@2989.4]
  assign _T_452 = _T_442 | _T_155; // @[NV_NVDLA_CDMA_wt.scala 490:29:@2996.4]
  assign _T_453 = _T_452 | _T_413; // @[NV_NVDLA_CDMA_wt.scala 490:41:@2997.4]
  assign _GEN_40 = _T_453 ? _T_451 : _T_422; // @[NV_NVDLA_CDMA_wt.scala 490:60:@2998.4]
  assign _T_458 = _T_456 + 18'h1; // @[NV_NVDLA_CDMA_wt.scala 501:49:@3002.4]
  assign _T_459 = _T_456 + 18'h1; // @[NV_NVDLA_CDMA_wt.scala 501:49:@3003.4]
  assign _T_460 = _T_456[13]; // @[NV_NVDLA_CDMA_wt.scala 502:49:@3004.4]
  assign _T_461 = ~ _T_460; // @[NV_NVDLA_CDMA_wt.scala 502:31:@3005.4]
  assign _GEN_41 = _T_461 ? _T_459 : _T_456; // @[NV_NVDLA_CDMA_wt.scala 506:30:@3008.4]
  assign _T_463 = _T_413 | _T_461; // @[NV_NVDLA_CDMA_wt.scala 510:48:@3011.4]
  assign _T_471 = _T_422[16:1]; // @[NV_NVDLA_CDMA_wt.scala 518:70:@3015.4]
  assign _T_473 = _T_456[16:1]; // @[NV_NVDLA_CDMA_wt.scala 519:118:@3016.4]
  assign _T_474 = 16'h1000 + _T_473; // @[NV_NVDLA_CDMA_wt.scala 519:99:@3017.4]
  assign _T_475 = 16'h1000 + _T_473; // @[NV_NVDLA_CDMA_wt.scala 519:99:@3018.4]
  assign _T_476 = _T_413 ? _T_471 : _T_475; // @[NV_NVDLA_CDMA_wt.scala 518:37:@3019.4]
  assign _T_477 = _T_422[0]; // @[NV_NVDLA_CDMA_wt.scala 520:73:@3021.4]
  assign _T_478 = _T_456[0]; // @[NV_NVDLA_CDMA_wt.scala 520:129:@3022.4]
  assign _T_479 = _T_413 ? _T_477 : _T_478; // @[NV_NVDLA_CDMA_wt.scala 520:40:@3023.4]
  assign _GEN_73 = {{1'd0}, _T_479}; // @[NV_NVDLA_CDMA_wt.scala 522:118:@3026.6]
  assign _T_481 = _GEN_73 == 2'h2; // @[NV_NVDLA_CDMA_wt.scala 522:118:@3026.6]
  assign _T_492 = {_T_481,_T_481}; // @[NV_NVDLA_CDMA_wt.scala 522:150:@3031.6]
  assign _GEN_42 = _T_463 ? _T_492 : _T_468; // @[NV_NVDLA_CDMA_wt.scala 521:34:@3025.4]
  assign _T_494 = _T_413 ? _T_398 : 256'h0; // @[NV_NVDLA_CDMA_wt.scala 531:36:@3035.4]
  assign _T_465 = {{1'd0}, _T_476}; // @[NV_NVDLA_CDMA_wt.scala 511:37:@3012.4 NV_NVDLA_CDMA_wt.scala 518:31:@3020.4]
  assign _GEN_43 = _T_463 ? _T_465 : _T_500; // @[Reg.scala 20:19:@3040.4]
  assign _GEN_44 = _T_463 ? _T_494 : _T_503; // @[Reg.scala 20:19:@3045.4]
  assign _GEN_45 = io_sc2cdma_wt_updt_valid ? io_sc2cdma_wt_updt_bits_entries : _T_354; // @[NV_NVDLA_CDMA_wt.scala 548:35:@3052.4]
  assign _T_514 = _T_311 & _T_250; // @[NV_NVDLA_CDMA_wt.scala 556:50:@3059.4]
  assign _T_515 = ~ _T_247; // @[NV_NVDLA_CDMA_wt.scala 556:74:@3060.4]
  assign _T_516 = _T_514 & _T_515; // @[NV_NVDLA_CDMA_wt.scala 556:72:@3061.4]
  assign _T_518 = _T_516 ? _T_238 : 4'h0; // @[NV_NVDLA_CDMA_wt.scala 556:32:@3062.4]
  assign _T_521 = _T_413 ? 3'h1 : 3'h0; // @[NV_NVDLA_CDMA_wt.scala 557:32:@3063.4]
  assign _T_624 = _T_560 - _T_615; // @[NV_NVDLA_CDMA_wt.scala 647:39:@3154.4]
  assign _T_625 = $unsigned(_T_624); // @[NV_NVDLA_CDMA_wt.scala 647:39:@3155.4]
  assign _T_626 = _T_625[25:0]; // @[NV_NVDLA_CDMA_wt.scala 647:39:@3156.4]
  assign _T_627 = _T_626[15:1]; // @[NV_NVDLA_CDMA_wt.scala 652:41:@3157.4]
  assign _T_523 = {_T_627,1'h0}; // @[Cat.scala 30:58:@3064.4]
  assign _T_605 = ~ _T_563; // @[NV_NVDLA_CDMA_wt.scala 622:26:@3136.4]
  assign _T_597 = {_T_560,8'h0}; // @[Cat.scala 30:58:@3129.4]
  assign _GEN_75 = {{2'd0}, _T_566}; // @[NV_NVDLA_CDMA_wt.scala 618:95:@3130.4]
  assign _T_598 = _T_597 >= _GEN_75; // @[NV_NVDLA_CDMA_wt.scala 618:95:@3130.4]
  assign _T_599 = _T_153 & _T_598; // @[NV_NVDLA_CDMA_wt.scala 618:35:@3131.4]
  assign _T_600 = _T_560[1:0]; // @[NV_NVDLA_CDMA_wt.scala 619:40:@3132.4]
  assign _T_602 = _T_600 != 2'h0; // @[NV_NVDLA_CDMA_wt.scala 619:70:@3133.4]
  assign _T_603 = ~ _T_602; // @[NV_NVDLA_CDMA_wt.scala 619:24:@3134.4]
  assign _T_604 = _T_599 & _T_603; // @[NV_NVDLA_CDMA_wt.scala 618:117:@3135.4]
  assign _T_607 = _T_605 ? 1'h0 : _T_604; // @[NV_NVDLA_CDMA_wt.scala 622:25:@3137.4]
  assign _T_525 = _T_607 ? {{1'd0}, _T_523} : 17'h0; // @[NV_NVDLA_CDMA_wt.scala 563:34:@3065.4]
  assign _T_527 = {_T_354,1'h0}; // @[Cat.scala 30:58:@3067.4]
  assign _T_529 = _T_351 ? {{1'd0}, _T_527} : 17'h0; // @[NV_NVDLA_CDMA_wt.scala 564:31:@3068.4]
  assign _GEN_76 = {{10'd0}, _T_518}; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3070.4]
  assign _T_530 = _T_289 + _GEN_76; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3070.4]
  assign _T_531 = _T_289 + _GEN_76; // @[NV_NVDLA_CDMA_wt.scala 571:41:@3071.4]
  assign _GEN_77 = {{11'd0}, _T_521}; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3072.4]
  assign _T_532 = _T_531 - _GEN_77; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3072.4]
  assign _T_533 = $unsigned(_T_532); // @[NV_NVDLA_CDMA_wt.scala 571:61:@3073.4]
  assign _T_534 = _T_533[13:0]; // @[NV_NVDLA_CDMA_wt.scala 571:61:@3074.4]
  assign _GEN_78 = {{14'd0}, _T_521}; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3075.4]
  assign _T_535 = _T_292 + _GEN_78; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3075.4]
  assign _T_536 = _T_292 + _GEN_78; // @[NV_NVDLA_CDMA_wt.scala 572:43:@3076.4]
  assign _T_537 = _T_536 - _T_525; // @[NV_NVDLA_CDMA_wt.scala 572:63:@3077.4]
  assign _T_538 = $unsigned(_T_537); // @[NV_NVDLA_CDMA_wt.scala 572:63:@3078.4]
  assign _T_539 = _T_538[16:0]; // @[NV_NVDLA_CDMA_wt.scala 572:63:@3079.4]
  assign _T_541 = _T_295 + _T_525; // @[NV_NVDLA_CDMA_wt.scala 573:57:@3080.4]
  assign _T_542 = _T_295 + _T_525; // @[NV_NVDLA_CDMA_wt.scala 573:57:@3081.4]
  assign _T_543 = _T_542 - _T_529; // @[NV_NVDLA_CDMA_wt.scala 573:78:@3082.4]
  assign _T_544 = $unsigned(_T_543); // @[NV_NVDLA_CDMA_wt.scala 573:78:@3083.4]
  assign _T_545 = _T_544[16:0]; // @[NV_NVDLA_CDMA_wt.scala 573:78:@3084.4]
  assign _T_546 = _T_155 ? 17'h0 : _T_545; // @[NV_NVDLA_CDMA_wt.scala 573:28:@3085.4]
  assign _T_548 = _T_514 | _T_413; // @[NV_NVDLA_CDMA_wt.scala 574:74:@3087.4]
  assign _GEN_46 = _T_548 ? _T_534 : _T_289; // @[NV_NVDLA_CDMA_wt.scala 576:31:@3088.4]
  assign _T_549 = _T_413 | _T_607; // @[NV_NVDLA_CDMA_wt.scala 579:27:@3091.4]
  assign _GEN_47 = _T_549 ? _T_539 : _T_292; // @[NV_NVDLA_CDMA_wt.scala 579:43:@3092.4]
  assign _T_550 = _T_607 | _T_351; // @[NV_NVDLA_CDMA_wt.scala 582:24:@3095.4]
  assign _T_551 = _T_550 | _T_155; // @[NV_NVDLA_CDMA_wt.scala 582:37:@3096.4]
  assign _GEN_48 = _T_551 ? _T_546 : _T_295; // @[NV_NVDLA_CDMA_wt.scala 582:49:@3097.4]
  assign _T_568 = _T_554 + 12'h1; // @[NV_NVDLA_CDMA_wt.scala 595:49:@3105.4]
  assign _T_569 = _T_554 + 12'h1; // @[NV_NVDLA_CDMA_wt.scala 595:49:@3106.4]
  assign _T_570 = _T_569 == _T_168; // @[NV_NVDLA_CDMA_wt.scala 596:51:@3107.4]
  assign _T_572 = _T_152 ? 12'h0 : _T_569; // @[NV_NVDLA_CDMA_wt.scala 597:33:@3108.4]
  assign _T_575 = _T_570 ? 1'h1 : _T_119; // @[NV_NVDLA_CDMA_wt.scala 599:28:@3109.4]
  assign _T_576 = _T_152 ? 1'h0 : _T_575; // @[NV_NVDLA_CDMA_wt.scala 598:28:@3110.4]
  assign _T_578 = {_T_189,6'h0}; // @[Cat.scala 30:58:@3111.4]
  assign _GEN_79 = {{7'd0}, _T_578}; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3112.4]
  assign _T_580 = _T_557 + _GEN_79; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3112.4]
  assign _T_581 = _T_557 + _GEN_79; // @[NV_NVDLA_CDMA_wt.scala 604:53:@3113.4]
  assign _T_582 = _T_570 ? io_reg2dp_weight_bytes : _T_581; // @[NV_NVDLA_CDMA_wt.scala 603:34:@3114.4]
  assign _T_583 = _T_152 ? 32'h0 : _T_582; // @[NV_NVDLA_CDMA_wt.scala 602:34:@3115.4]
  assign _T_584 = ~ _T_607; // @[NV_NVDLA_CDMA_wt.scala 605:41:@3116.4]
  assign _T_585 = _T_153 & _T_584; // @[NV_NVDLA_CDMA_wt.scala 605:39:@3117.4]
  assign _T_587 = _T_605 & _T_585; // @[NV_NVDLA_CDMA_wt.scala 606:42:@3119.4]
  assign _T_589 = _T_152 ? 32'h0 : _T_566; // @[NV_NVDLA_CDMA_wt.scala 607:38:@3120.4]
  assign _T_590 = _T_152 | _T_587; // @[NV_NVDLA_CDMA_wt.scala 611:19:@3122.4]
  assign _GEN_49 = _T_590 ? _T_583 : _T_566; // @[NV_NVDLA_CDMA_wt.scala 611:36:@3123.4]
  assign _T_592 = _T_560 + 26'h1; // @[NV_NVDLA_CDMA_wt.scala 615:45:@3126.4]
  assign _T_593 = _T_560 + 26'h1; // @[NV_NVDLA_CDMA_wt.scala 615:45:@3127.4]
  assign _T_595 = _T_152 ? 26'h0 : _T_593; // @[NV_NVDLA_CDMA_wt.scala 616:31:@3128.4]
  assign _T_608 = _T_152 | _T_607; // @[NV_NVDLA_CDMA_wt.scala 624:19:@3139.4]
  assign _GEN_50 = _T_608 ? _T_572 : _T_554; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  assign _GEN_51 = _T_608 ? _T_576 : _T_119; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  assign _GEN_52 = _T_608 ? _T_589 : _T_557; // @[NV_NVDLA_CDMA_wt.scala 624:35:@3140.4]
  assign _T_609 = _T_152 | _T_413; // @[NV_NVDLA_CDMA_wt.scala 629:19:@3145.4]
  assign _GEN_53 = _T_609 ? _T_595 : _T_560; // @[NV_NVDLA_CDMA_wt.scala 629:38:@3146.4]
  assign _T_623 = _T_570 ? 26'h0 : _T_560; // @[NV_NVDLA_CDMA_wt.scala 646:35:@3153.4]
  assign _T_628 = ~ _T_570; // @[NV_NVDLA_CDMA_wt.scala 655:33:@3159.4]
  assign _T_630 = io_reg2dp_weight_kernel[5:0]; // @[NV_NVDLA_CDMA_wt.scala 656:52:@3160.4]
  assign _T_632 = _T_630 + 6'h1; // @[NV_NVDLA_CDMA_wt.scala 656:71:@3161.4]
  assign _T_633 = _T_628 ? 7'h20 : _T_632; // @[NV_NVDLA_CDMA_wt.scala 655:32:@3162.4]
  assign _GEN_54 = _T_607 ? _T_623 : _T_615; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  assign _GEN_55 = _T_607 ? _T_627 : _T_618; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  assign _GEN_56 = _T_607 ? _T_633 : {{1'd0}, _T_621}; // @[NV_NVDLA_CDMA_wt.scala 659:24:@3164.4]
  assign _GEN_57 = _T_612 ? _T_618 : _T_660; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3185.4]
  assign _GEN_58 = _T_612 ? _T_621 : _T_649; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3185.4]
  assign _GEN_59 = _T_638 ? _T_660 : _T_663; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3190.4]
  assign _GEN_60 = _T_638 ? _T_649 : _T_652; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3190.4]
  assign _GEN_61 = _T_641 ? _T_663 : _T_666; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3195.4]
  assign _GEN_62 = _T_641 ? _T_652 : _T_655; // @[NV_NVDLA_CDMA_wt.scala 677:32:@3195.4]
  assign _T_667 = ~ _T_313; // @[NV_NVDLA_CDMA_wt.scala 692:52:@3202.4]
  assign _T_668 = _T_333 & _T_667; // @[NV_NVDLA_CDMA_wt.scala 692:50:@3203.4]
  assign _T_669 = _T_668 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_wt.scala 692:68:@3204.4]
  assign _T_673 = io_status2dma_fsm_switch & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_wt.scala 693:60:@3207.4]
  assign _T_677 = io_reg2dp_op_en & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_wt.scala 694:51:@3210.4]
  assign _T_688 = _T_410 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_wt.scala 708:56:@3227.4]
  assign _T_700 = NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_wt.scala 712:41:@3235.4 NV_NVDLA_CDMA_wt.scala 722:31:@3248.4]
  assign _T_702 = _T_700 != 9'h1ff; // @[NV_NVDLA_CDMA_wt.scala 713:48:@3236.4]
  assign io_cdma_wt2mcif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 305:31:@2837.4]
  assign io_cdma_wt2mcif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 305:31:@2836.4]
  assign io_mcif2cdma_wt_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 316:47:@2851.4]
  assign io_cdma_wt2cvif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 303:39:@2834.4]
  assign io_cdma_wt2cvif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 303:39:@2833.4]
  assign io_cvif2cdma_wt_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 314:55:@2848.4]
  assign io_cdma2buf_wt_wr_sel = _T_468; // @[NV_NVDLA_CDMA_wt.scala 524:35:@3034.4]
  assign io_cdma2buf_wt_wr_addr_valid = _T_497; // @[NV_NVDLA_CDMA_wt.scala 532:34:@3038.4]
  assign io_cdma2buf_wt_wr_addr_bits = _T_500; // @[NV_NVDLA_CDMA_wt.scala 533:33:@3043.4]
  assign io_cdma2buf_wt_wr_data = _T_503; // @[NV_NVDLA_CDMA_wt.scala 537:28:@3048.4]
  assign io_wt2status_state = _T_141; // @[NV_NVDLA_CDMA_wt.scala 160:24:@2699.4]
  assign io_cdma2sc_wt_updt_valid = _T_644; // @[NV_NVDLA_CDMA_wt.scala 684:30:@3199.4]
  assign io_cdma2sc_wt_updt_bits_entries = _T_666; // @[NV_NVDLA_CDMA_wt.scala 686:37:@3201.4]
  assign io_cdma2sc_wt_updt_bits_kernels = {{8'd0}, _T_655}; // @[NV_NVDLA_CDMA_wt.scala 685:37:@3200.4]
  assign io_cdma2sc_wt_pending_ack = _T_150; // @[NV_NVDLA_CDMA_wt.scala 161:31:@2700.4]
  assign io_dp2reg_wt_flush_done = _T_456[13]; // @[NV_NVDLA_CDMA_wt.scala 504:29:@3007.4]
  assign io_dp2reg_wt_rd_stall = NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_wt.scala 704:27:@3221.4]
  assign NV_NVDLA_DMAIF_rdreq_reset = reset; // @[:@2830.4]
  assign NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 300:47:@2831.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid = _T_320 & _T_315; // @[NV_NVDLA_CDMA_wt.scala 308:54:@2840.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits = {_T_337,_T_335}; // @[NV_NVDLA_CDMA_wt.scala 307:53:@2839.4]
  assign NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready = io_cdma_wt2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 305:31:@2838.4]
  assign NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready = io_cdma_wt2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_wt.scala 303:39:@2835.4]
  assign NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type = io_reg2dp_weight_ram_type; // @[NV_NVDLA_CDMA_wt.scala 301:52:@2832.4]
  assign NV_NVDLA_DMAIF_rdrsp_reset = reset; // @[:@2844.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 312:47:@2845.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid = io_mcif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 316:47:@2850.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits = io_mcif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 316:47:@2849.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid = io_cvif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_wt.scala 314:55:@2847.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits = io_cvif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 314:55:@2846.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready = NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_wt.scala 329:54:@2859.4]
  assign NV_NVDLA_fifo_clock = io_nvdla_core_clk; // @[:@2854.4]
  assign NV_NVDLA_fifo_reset = reset; // @[:@2855.4]
  assign NV_NVDLA_fifo_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 326:25:@2856.4]
  assign NV_NVDLA_fifo_io_wr_pvld = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits[0]; // @[NV_NVDLA_CDMA_wt.scala 328:29:@2858.4]
  assign NV_NVDLA_fifo_io_wr_pd = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_wt.scala 330:27:@2860.4]
  assign NV_NVDLA_fifo_io_rd_prdy = _T_357 < _GEN_68; // @[NV_NVDLA_CDMA_wt.scala 332:29:@2861.4]
  assign NV_NVDLA_fifo_1_clock = io_nvdla_core_clk; // @[:@2931.4]
  assign NV_NVDLA_fifo_1_reset = reset; // @[:@2932.4]
  assign NV_NVDLA_fifo_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 395:19:@2933.4]
  assign NV_NVDLA_fifo_1_io_wr_pvld = _T_320 & _T_313; // @[NV_NVDLA_CDMA_wt.scala 398:23:@2935.4]
  assign NV_NVDLA_fifo_1_io_wr_pd = {2'h0,_T_278}; // @[NV_NVDLA_CDMA_wt.scala 400:21:@2937.4]
  assign NV_NVDLA_fifo_1_io_rd_prdy = _T_411 & _T_405; // @[NV_NVDLA_CDMA_wt.scala 402:23:@2938.4]
  assign NV_COUNTER_STAGE_histogram_reset = reset; // @[:@3215.4]
  assign NV_COUNTER_STAGE_histogram_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 699:16:@3216.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_inc = _T_672; // @[NV_NVDLA_CDMA_wt.scala 700:25:@3217.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_clr = _T_676; // @[NV_NVDLA_CDMA_wt.scala 702:25:@3219.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_cen = _T_680; // @[NV_NVDLA_CDMA_wt.scala 703:25:@3220.4]
  assign NV_COUNTER_STAGE_histogram_1_reset = reset; // @[:@3242.4]
  assign NV_COUNTER_STAGE_histogram_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_wt.scala 717:18:@3243.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc = _T_702 & _T_687; // @[NV_NVDLA_CDMA_wt.scala 718:27:@3244.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec = _T_702 & _T_691; // @[NV_NVDLA_CDMA_wt.scala 719:27:@3245.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr = _T_694; // @[NV_NVDLA_CDMA_wt.scala 720:27:@3246.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen = _T_698; // @[NV_NVDLA_CDMA_wt.scala 721:27:@3247.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_83 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_89 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_105 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_112 = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_147 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_144 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_119 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_122 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_141 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_150 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_168 = _RAND_10[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_175 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_182 = _RAND_12[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_189 = _RAND_13[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_209 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_212 = _RAND_15[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_215 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_272 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_289 = _RAND_18[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_292 = _RAND_19[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_295 = _RAND_20[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_284 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_235 = _RAND_22[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_238 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_241 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_244 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_247 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_250 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_275 = _RAND_28[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_278 = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_281 = _RAND_30[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_342 = _RAND_31[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_357 = _RAND_32[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_351 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_354 = _RAND_34[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_397 = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_422 = _RAND_36[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_456 = _RAND_37[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_468 = _RAND_38[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_497 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_500 = _RAND_40[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {8{`RANDOM}};
  _T_503 = _RAND_41[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_560 = _RAND_42[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_615 = _RAND_43[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_563 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_566 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_554 = _RAND_46[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_557 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_612 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_618 = _RAND_49[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_621 = _RAND_50[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_638 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_641 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_644 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_649 = _RAND_54[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_652 = _RAND_55[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_655 = _RAND_56[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_660 = _RAND_57[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_663 = _RAND_58[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_666 = _RAND_59[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_672 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_676 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_680 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_687 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_691 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_694 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_698 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_83 <= 1'h0;
    end else begin
      if (io_status2dma_fsm_switch) begin
        _T_83 <= io_reg2dp_skip_weight_rls;
      end
    end
    if (reset) begin
      _T_89 <= 2'h0;
    end else begin
      if (_T_92) begin
        if (_T_93) begin
          _T_89 <= 2'h1;
        end else begin
          if (_T_95) begin
            _T_89 <= 2'h3;
          end else begin
            if (io_reg2dp_op_en) begin
              _T_89 <= 2'h2;
            end else begin
              _T_89 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_158) begin
            _T_89 <= 2'h2;
          end else begin
            _T_89 <= 2'h0;
          end
        end else begin
          if (_T_97) begin
            if (_T_134) begin
              _T_89 <= 2'h3;
            end else begin
              _T_89 <= 2'h0;
            end
          end else begin
            _T_89 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_105 <= 5'h1f;
    end else begin
      if (io_status2dma_fsm_switch) begin
        _T_105 <= io_reg2dp_data_bank;
      end
    end
    if (reset) begin
      _T_112 <= 5'h1f;
    end else begin
      if (io_status2dma_fsm_switch) begin
        _T_112 <= io_reg2dp_weight_bank;
      end
    end
    if (reset) begin
      _T_147 <= 1'h0;
    end else begin
      _T_147 <= _T_144;
    end
    if (reset) begin
      _T_144 <= 1'h0;
    end else begin
      _T_144 <= io_sc2cdma_wt_pending_req;
    end
    if (reset) begin
      _T_119 <= 1'h0;
    end else begin
      if (_T_608) begin
        if (_T_152) begin
          _T_119 <= 1'h0;
        end else begin
          if (_T_570) begin
            _T_119 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_122 <= 4'h0;
    end else begin
      if (_T_138) begin
        if (_T_152) begin
          _T_122 <= 4'h0;
        end else begin
          if (_T_126) begin
            _T_122 <= _T_129;
          end
        end
      end
    end
    if (reset) begin
      _T_141 <= 2'h0;
    end else begin
      if (_T_92) begin
        if (_T_93) begin
          _T_141 <= 2'h1;
        end else begin
          if (_T_95) begin
            _T_141 <= 2'h3;
          end else begin
            if (io_reg2dp_op_en) begin
              _T_141 <= 2'h2;
            end else begin
              _T_141 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_158) begin
            _T_141 <= 2'h2;
          end else begin
            _T_141 <= 2'h0;
          end
        end else begin
          if (_T_97) begin
            if (_T_134) begin
              _T_141 <= 2'h3;
            end else begin
              _T_141 <= 2'h0;
            end
          end else begin
            _T_141 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_150 <= 1'h0;
    end else begin
      _T_150 <= _T_154;
    end
    if (reset) begin
      _T_168 <= 12'hfff;
    end else begin
      if (_T_152) begin
        _T_168 <= {{4'd0}, _T_194};
      end
    end
    if (reset) begin
      _T_175 <= 6'h3f;
    end else begin
      if (_T_152) begin
        _T_175 <= _T_198;
      end
    end
    if (reset) begin
      _T_182 <= 7'h7f;
    end else begin
      if (_T_152) begin
        _T_182 <= _T_199;
      end
    end
    if (_T_152) begin
      _T_189 <= _T_187;
    end
    if (reset) begin
      _T_209 <= 4'h0;
    end else begin
      if (_T_311) begin
        if (_T_230) begin
          _T_209 <= _T_231;
        end else begin
          if (_T_152) begin
            _T_209 <= _T_227;
          end else begin
            _T_209 <= 4'h8;
          end
        end
      end
    end
    if (reset) begin
      _T_212 <= 29'h0;
    end else begin
      if (_T_311) begin
        if (_T_152) begin
          _T_212 <= {{2'd0}, _T_221};
        end else begin
          _T_212 <= _T_220;
        end
      end
    end
    if (reset) begin
      _T_215 <= 1'h0;
    end else begin
      _T_215 <= _T_156;
    end
    if (reset) begin
      _T_272 <= 1'h0;
    end else begin
      _T_272 <= _T_285;
    end
    if (reset) begin
      _T_284 <= 1'h1;
    end else begin
      if (_T_311) begin
        _T_284 <= _T_286;
      end
    end
    if (reset) begin
      _T_235 <= 59'h0;
    end else begin
      _T_235 <= _GEN_21[58:0];
    end
    if (reset) begin
      _T_238 <= 4'h0;
    end else begin
      if (_T_311) begin
        _T_238 <= _T_209;
      end
    end
    if (reset) begin
      _T_241 <= 3'h0;
    end else begin
      _T_241 <= _GEN_23[2:0];
    end
    if (reset) begin
      _T_244 <= 1'h0;
    end else begin
      if (_T_311) begin
        _T_244 <= _T_252;
      end
    end
    if (reset) begin
      _T_247 <= 1'h1;
    end else begin
      if (_T_311) begin
        if (_T_152) begin
          _T_247 <= 1'h0;
        end else begin
          if (_T_244) begin
            _T_247 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_250 <= 1'h0;
    end else begin
      _T_250 <= _T_269;
    end
    if (reset) begin
      _T_275 <= 59'h0;
    end else begin
      if (_T_311) begin
        _T_275 <= _T_235;
      end
    end
    if (reset) begin
      _T_278 <= 4'h0;
    end else begin
      if (_T_311) begin
        _T_278 <= _T_238;
      end
    end
    if (reset) begin
      _T_281 <= 3'h0;
    end else begin
      if (_T_311) begin
        _T_281 <= _T_241;
      end
    end
    if (reset) begin
      _T_342 <= 4'h0;
    end else begin
      if (_T_413) begin
        if (_T_344) begin
          _T_342 <= 4'h0;
        end else begin
          _T_342 <= _T_348;
        end
      end
    end
    if (reset) begin
      _T_357 <= 17'h0;
    end else begin
      if (_T_360) begin
        if (_T_344) begin
          _T_357 <= _T_365;
        end
      end else begin
        if (_T_366) begin
          if (_T_344) begin
            _T_357 <= _T_374;
          end else begin
            _T_357 <= _T_377;
          end
        end else begin
          if (_T_380) begin
            _T_357 <= _T_377;
          end
        end
      end
    end
    if (reset) begin
      _T_397 <= 4'h0;
    end else begin
      if (_T_411) begin
        if (_T_405) begin
          _T_397 <= 4'h0;
        end else begin
          _T_397 <= _T_404;
        end
      end
    end
    if (reset) begin
      _T_422 <= 17'h0;
    end else begin
      if (_T_453) begin
        if (_T_447) begin
          _T_422 <= {{1'd0}, _T_449};
        end else begin
          _T_422 <= _T_438;
        end
      end
    end
    if (reset) begin
      _T_503 <= 256'h0;
    end else begin
      if (_T_463) begin
        if (_T_413) begin
          _T_503 <= _T_398;
        end else begin
          _T_503 <= 256'h0;
        end
      end
    end
    if (reset) begin
      _T_560 <= 26'h0;
    end else begin
      if (_T_609) begin
        if (_T_152) begin
          _T_560 <= 26'h0;
        end else begin
          _T_560 <= _T_593;
        end
      end
    end
    if (reset) begin
      _T_615 <= 26'h0;
    end else begin
      if (_T_607) begin
        if (_T_570) begin
          _T_615 <= 26'h0;
        end else begin
          _T_615 <= _T_560;
        end
      end
    end
    if (reset) begin
      _T_563 <= 1'h0;
    end else begin
      _T_563 <= _T_585;
    end
    if (reset) begin
      _T_566 <= 32'h0;
    end else begin
      if (_T_590) begin
        if (_T_152) begin
          _T_566 <= 32'h0;
        end else begin
          if (_T_570) begin
            _T_566 <= io_reg2dp_weight_bytes;
          end else begin
            _T_566 <= _T_581;
          end
        end
      end
    end
    if (reset) begin
      _T_554 <= 12'h0;
    end else begin
      if (_T_608) begin
        if (_T_152) begin
          _T_554 <= 12'h0;
        end else begin
          _T_554 <= _T_569;
        end
      end
    end
    if (reset) begin
      _T_557 <= 32'h0;
    end else begin
      if (_T_608) begin
        if (_T_152) begin
          _T_557 <= 32'h0;
        end else begin
          _T_557 <= _T_566;
        end
      end
    end
    if (reset) begin
      _T_612 <= 1'h0;
    end else begin
      if (_T_605) begin
        _T_612 <= 1'h0;
      end else begin
        _T_612 <= _T_604;
      end
    end
    if (reset) begin
      _T_618 <= 15'h0;
    end else begin
      if (_T_607) begin
        _T_618 <= _T_627;
      end
    end
    if (reset) begin
      _T_621 <= 6'h0;
    end else begin
      _T_621 <= _GEN_56[5:0];
    end
    if (reset) begin
      _T_638 <= 1'h0;
    end else begin
      _T_638 <= _T_612;
    end
    if (reset) begin
      _T_641 <= 1'h0;
    end else begin
      _T_641 <= _T_638;
    end
    if (reset) begin
      _T_644 <= 1'h0;
    end else begin
      _T_644 <= _T_641;
    end
    if (reset) begin
      _T_649 <= 6'h0;
    end else begin
      if (_T_612) begin
        _T_649 <= _T_621;
      end
    end
    if (reset) begin
      _T_652 <= 6'h0;
    end else begin
      if (_T_638) begin
        _T_652 <= _T_649;
      end
    end
    if (reset) begin
      _T_655 <= 6'h0;
    end else begin
      if (_T_641) begin
        _T_655 <= _T_652;
      end
    end
    if (reset) begin
      _T_660 <= 15'h0;
    end else begin
      if (_T_612) begin
        _T_660 <= _T_618;
      end
    end
    if (reset) begin
      _T_663 <= 15'h0;
    end else begin
      if (_T_638) begin
        _T_663 <= _T_660;
      end
    end
    if (reset) begin
      _T_666 <= 15'h0;
    end else begin
      if (_T_641) begin
        _T_666 <= _T_663;
      end
    end
    if (reset) begin
      _T_672 <= 1'h0;
    end else begin
      _T_672 <= _T_669;
    end
    if (reset) begin
      _T_676 <= 1'h0;
    end else begin
      _T_676 <= _T_673;
    end
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
    if (reset) begin
      _T_687 <= 1'h0;
    end else begin
      _T_687 <= _T_669;
    end
    if (reset) begin
      _T_691 <= 1'h0;
    end else begin
      _T_691 <= _T_688;
    end
    if (reset) begin
      _T_694 <= 1'h0;
    end else begin
      _T_694 <= io_status2dma_fsm_switch;
    end
    if (reset) begin
      _T_698 <= 1'h0;
    end else begin
      _T_698 <= _T_677;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_289 <= 14'h0;
    end else begin
      if (_T_548) begin
        _T_289 <= _T_534;
      end
    end
    if (reset) begin
      _T_292 <= 17'h0;
    end else begin
      if (_T_549) begin
        _T_292 <= _T_539;
      end
    end
    if (reset) begin
      _T_295 <= 17'h0;
    end else begin
      if (_T_551) begin
        if (_T_155) begin
          _T_295 <= 17'h0;
        end else begin
          _T_295 <= _T_545;
        end
      end
    end
    if (reset) begin
      _T_351 <= 1'h0;
    end else begin
      _T_351 <= io_sc2cdma_wt_updt_valid;
    end
    if (reset) begin
      _T_354 <= 15'h0;
    end else begin
      if (io_sc2cdma_wt_updt_valid) begin
        _T_354 <= io_sc2cdma_wt_updt_bits_entries;
      end
    end
    if (reset) begin
      _T_456 <= 18'h0;
    end else begin
      if (_T_461) begin
        _T_456 <= _T_459;
      end
    end
    if (reset) begin
      _T_468 <= 2'h0;
    end else begin
      if (_T_463) begin
        _T_468 <= _T_492;
      end
    end
    if (reset) begin
      _T_497 <= 1'h0;
    end else begin
      _T_497 <= _T_463;
    end
    if (reset) begin
      _T_500 <= 17'h0;
    end else begin
      if (_T_463) begin
        _T_500 <= _T_465;
      end
    end
  end
endmodule
module NV_NVDLA_slcg( // @[:@3250.2]
  input   io_nvdla_clock_nvdla_core_clk, // @[:@3253.4]
  output  io_nvdla_core_gated_clk // @[:@3253.4]
);
  assign io_nvdla_core_gated_clk = io_nvdla_clock_nvdla_core_clk; // @[slcg.scala 23:31:@3255.4]
endmodule
module NV_NVDLA_CDMA_dc( // @[:@3869.2]
  input          reset, // @[:@3871.4]
  input          io_nvdla_core_clk, // @[:@3872.4]
  input          io_nvdla_core_ng_clk, // @[:@3872.4]
  input          io_dc_dat2mcif_rd_req_pd_ready, // @[:@3872.4]
  output         io_dc_dat2mcif_rd_req_pd_valid, // @[:@3872.4]
  output [78:0]  io_dc_dat2mcif_rd_req_pd_bits, // @[:@3872.4]
  output         io_mcif2dc_dat_rd_rsp_pd_ready, // @[:@3872.4]
  input          io_mcif2dc_dat_rd_rsp_pd_valid, // @[:@3872.4]
  input  [256:0] io_mcif2dc_dat_rd_rsp_pd_bits, // @[:@3872.4]
  input          io_dc_dat2cvif_rd_req_pd_ready, // @[:@3872.4]
  output         io_dc_dat2cvif_rd_req_pd_valid, // @[:@3872.4]
  output [78:0]  io_dc_dat2cvif_rd_req_pd_bits, // @[:@3872.4]
  output         io_cvif2dc_dat_rd_rsp_pd_ready, // @[:@3872.4]
  input          io_cvif2dc_dat_rd_rsp_pd_valid, // @[:@3872.4]
  input  [256:0] io_cvif2dc_dat_rd_rsp_pd_bits, // @[:@3872.4]
  output         io_dc2cvt_dat_wr_sel, // @[:@3872.4]
  output         io_dc2cvt_dat_wr_addr_valid, // @[:@3872.4]
  output [16:0]  io_dc2cvt_dat_wr_addr_bits, // @[:@3872.4]
  output [255:0] io_dc2cvt_dat_wr_data, // @[:@3872.4]
  output [11:0]  io_dc2cvt_dat_wr_info_pd, // @[:@3872.4]
  input          io_reg2dp_op_en, // @[:@3872.4]
  input          io_reg2dp_conv_mode, // @[:@3872.4]
  input          io_reg2dp_data_reuse, // @[:@3872.4]
  input          io_reg2dp_skip_data_rls, // @[:@3872.4]
  input          io_reg2dp_datain_format, // @[:@3872.4]
  input  [12:0]  io_reg2dp_datain_width, // @[:@3872.4]
  input  [12:0]  io_reg2dp_datain_height, // @[:@3872.4]
  input  [12:0]  io_reg2dp_datain_channel, // @[:@3872.4]
  input          io_reg2dp_datain_ram_type, // @[:@3872.4]
  input  [31:0]  io_reg2dp_datain_addr_high_0, // @[:@3872.4]
  input  [26:0]  io_reg2dp_datain_addr_low_0, // @[:@3872.4]
  input  [26:0]  io_reg2dp_line_stride, // @[:@3872.4]
  input  [26:0]  io_reg2dp_surf_stride, // @[:@3872.4]
  input  [26:0]  io_reg2dp_batch_stride, // @[:@3872.4]
  input          io_reg2dp_line_packed, // @[:@3872.4]
  input          io_reg2dp_surf_packed, // @[:@3872.4]
  input  [4:0]   io_reg2dp_batches, // @[:@3872.4]
  input  [16:0]  io_reg2dp_entries, // @[:@3872.4]
  input  [11:0]  io_reg2dp_grains, // @[:@3872.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@3872.4]
  input          io_reg2dp_dma_en, // @[:@3872.4]
  output [31:0]  io_dp2reg_dc_rd_stall, // @[:@3872.4]
  output [31:0]  io_dp2reg_dc_rd_latency, // @[:@3872.4]
  output [1:0]   io_dc2status_state, // @[:@3872.4]
  output         io_dc2status_dat_updt_valid, // @[:@3872.4]
  output [14:0]  io_dc2status_dat_updt_bits_entries, // @[:@3872.4]
  output [13:0]  io_dc2status_dat_updt_bits_slices, // @[:@3872.4]
  input          io_status2dma_fsm_switch, // @[:@3872.4]
  input  [14:0]  io_status2dma_free_entries, // @[:@3872.4]
  input  [14:0]  io_status2dma_wr_idx, // @[:@3872.4]
  output         io_dc2sbuf_p0_wr_addr_valid, // @[:@3872.4]
  output [7:0]   io_dc2sbuf_p0_wr_addr_bits, // @[:@3872.4]
  output [255:0] io_dc2sbuf_p0_wr_data, // @[:@3872.4]
  output         io_dc2sbuf_p0_rd_addr_valid, // @[:@3872.4]
  output [7:0]   io_dc2sbuf_p0_rd_addr_bits, // @[:@3872.4]
  input  [255:0] io_dc2sbuf_p0_rd_data, // @[:@3872.4]
  input          io_sc2cdma_dat_pending_req // @[:@3872.4]
);
  wire  NV_NVDLA_DMAIF_rdreq_reset; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type; // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
  wire  NV_NVDLA_DMAIF_rdrsp_reset; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
  wire  NV_NVDLA_fifo_clock; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_reset; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_io_clk; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_io_wr_pvld; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire [5:0] NV_NVDLA_fifo_io_wr_pd; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_NVDLA_fifo_io_rd_prdy; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire [5:0] NV_NVDLA_fifo_io_rd_pd; // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
  wire  NV_COUNTER_STAGE_histogram_reset; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire  NV_COUNTER_STAGE_histogram_io_clk; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_inc; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_clr; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_cen; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire [31:0] NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
  wire  NV_COUNTER_STAGE_histogram_1_reset; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_clk; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire [8:0] NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
  wire  NV_COUNTER_STAGE_histogram_2_reset; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_clk; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  wire [31:0] NV_COUNTER_STAGE_histogram_2_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
  reg  _T_85; // @[NV_NVDLA_CDMA_dc.scala 86:69:@3879.4]
  reg [31:0] _RAND_0;
  reg [1:0] _T_91; // @[NV_NVDLA_CDMA_dc.scala 89:28:@3880.4]
  reg [31:0] _RAND_1;
  wire  _T_94; // @[Conditional.scala 37:30:@3883.4]
  wire  _T_128; // @[NV_NVDLA_CDMA_dc.scala 123:38:@3938.4]
  wire  _T_129; // @[NV_NVDLA_CDMA_dc.scala 124:30:@3939.4]
  wire  _T_126; // @[NV_NVDLA_CDMA_dc.scala 122:47:@3937.4]
  wire  _T_130; // @[NV_NVDLA_CDMA_dc.scala 124:38:@3940.4]
  reg [4:0] _T_116; // @[NV_NVDLA_CDMA_dc.scala 116:65:@3927.4]
  reg [31:0] _RAND_2;
  wire  _T_123; // @[NV_NVDLA_CDMA_dc.scala 120:37:@3933.4]
  wire  _T_95; // @[NV_NVDLA_CDMA_dc.scala 94:21:@3885.6]
  wire  _T_96; // @[NV_NVDLA_CDMA_dc.scala 95:26:@3890.8]
  wire  _T_97; // @[NV_NVDLA_CDMA_dc.scala 95:49:@3891.8]
  reg  _T_119; // @[NV_NVDLA_CDMA_dc.scala 117:58:@3928.4]
  reg [31:0] _RAND_3;
  wire  _T_124; // @[NV_NVDLA_CDMA_dc.scala 121:25:@3935.4]
  wire  _T_98; // @[NV_NVDLA_CDMA_dc.scala 95:70:@3892.8]
  wire [1:0] _GEN_0; // @[NV_NVDLA_CDMA_dc.scala 96:27:@3897.10]
  wire [1:0] _GEN_1; // @[NV_NVDLA_CDMA_dc.scala 95:84:@3893.8]
  wire [1:0] _GEN_2; // @[NV_NVDLA_CDMA_dc.scala 94:37:@3886.6]
  wire  _T_99; // @[Conditional.scala 37:30:@3902.6]
  reg  _T_154; // @[NV_NVDLA_CDMA_dc.scala 150:65:@3967.4]
  reg [31:0] _RAND_4;
  reg  _T_151; // @[NV_NVDLA_CDMA_dc.scala 149:62:@3966.4]
  reg [31:0] _RAND_5;
  wire  _T_155; // @[NV_NVDLA_CDMA_dc.scala 152:41:@3968.4]
  wire  _T_156; // @[NV_NVDLA_CDMA_dc.scala 152:39:@3969.4]
  wire [1:0] _GEN_3; // @[NV_NVDLA_CDMA_dc.scala 99:32:@3904.8]
  wire  _T_100; // @[Conditional.scala 37:30:@3909.8]
  wire  _T_141; // @[NV_NVDLA_CDMA_dc.scala 139:30:@3957.4]
  wire  _T_909; // @[NV_NVDLA_CDMA_dc.scala 736:20:@4748.4]
  reg [13:0] _T_893; // @[NV_NVDLA_CDMA_dc.scala 728:32:@4735.4]
  reg [31:0] _RAND_6;
  reg [13:0] _T_201; // @[NV_NVDLA_CDMA_dc.scala 177:30:@4018.4]
  reg [31:0] _RAND_7;
  wire  _T_910; // @[NV_NVDLA_CDMA_dc.scala 736:54:@4749.4]
  wire  _T_911; // @[NV_NVDLA_CDMA_dc.scala 736:37:@4750.4]
  wire  _T_120; // @[NV_NVDLA_CDMA_dc.scala 119:30:@3929.4]
  reg [4:0] _T_108; // @[NV_NVDLA_CDMA_dc.scala 114:28:@3925.4]
  reg [31:0] _RAND_8;
  wire  _T_121; // @[NV_NVDLA_CDMA_dc.scala 119:57:@3930.4]
  wire  _T_122; // @[NV_NVDLA_CDMA_dc.scala 119:44:@3931.4]
  wire [1:0] _GEN_4; // @[NV_NVDLA_CDMA_dc.scala 102:27:@3911.10]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@3910.8]
  wire [1:0] _GEN_8; // @[Conditional.scala 39:67:@3903.6]
  wire [1:0] _GEN_9; // @[Conditional.scala 40:58:@3884.4]
  wire  _T_131; // @[NV_NVDLA_CDMA_dc.scala 126:10:@3942.4]
  wire [5:0] _T_134; // @[NV_NVDLA_CDMA_dc.scala 130:32:@3948.8]
  wire [4:0] _T_135; // @[NV_NVDLA_CDMA_dc.scala 130:32:@3949.8]
  wire [4:0] _GEN_10; // @[NV_NVDLA_CDMA_dc.scala 129:27:@3947.6]
  wire [4:0] _GEN_11; // @[NV_NVDLA_CDMA_dc.scala 126:22:@3943.4]
  wire  _T_139; // @[NV_NVDLA_CDMA_dc.scala 137:27:@3954.4]
  wire  _T_138; // @[NV_NVDLA_CDMA_dc.scala 136:26:@3953.4]
  wire  _T_143; // @[NV_NVDLA_CDMA_dc.scala 141:37:@3960.4]
  wire  _T_145; // @[NV_NVDLA_CDMA_dc.scala 142:40:@3962.4]
  reg [1:0] _T_148; // @[NV_NVDLA_CDMA_dc.scala 145:34:@3963.4]
  reg [31:0] _RAND_9;
  wire  _T_157; // @[NV_NVDLA_CDMA_dc.scala 154:26:@3971.4]
  wire  _T_158; // @[NV_NVDLA_CDMA_dc.scala 157:37:@3975.6]
  wire  _GEN_12; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  wire [4:0] _GEN_13; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  wire  _GEN_14; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  wire  _GEN_15; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  wire  _GEN_16; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  reg [15:0] _T_195; // @[NV_NVDLA_CDMA_dc.scala 175:29:@4016.4]
  reg [31:0] _RAND_10;
  reg [14:0] _T_198; // @[NV_NVDLA_CDMA_dc.scala 176:37:@4017.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_204; // @[NV_NVDLA_CDMA_dc.scala 178:29:@4019.4]
  reg [31:0] _RAND_12;
  reg [17:0] _T_207; // @[NV_NVDLA_CDMA_dc.scala 179:31:@4020.4]
  reg [31:0] _RAND_13;
  reg [12:0] _T_210; // @[NV_NVDLA_CDMA_dc.scala 180:30:@4021.4]
  reg [31:0] _RAND_14;
  reg [10:0] _T_213; // @[NV_NVDLA_CDMA_dc.scala 181:31:@4022.4]
  reg [31:0] _RAND_15;
  reg [38:0] _T_216; // @[NV_NVDLA_CDMA_dc.scala 182:29:@4023.4]
  reg [63:0] _RAND_16;
  reg [5:0] _T_219; // @[NV_NVDLA_CDMA_dc.scala 183:28:@4024.4]
  reg [31:0] _RAND_17;
  wire  _T_221; // @[NV_NVDLA_CDMA_dc.scala 185:49:@4025.4]
  wire  _T_223; // @[NV_NVDLA_CDMA_dc.scala 185:85:@4026.4]
  wire  _T_224; // @[NV_NVDLA_CDMA_dc.scala 185:58:@4027.4]
  wire  _T_225; // @[NV_NVDLA_CDMA_dc.scala 185:94:@4028.4]
  wire [7:0] _T_226; // @[NV_NVDLA_CDMA_dc.scala 186:52:@4029.4]
  wire [8:0] _T_228; // @[NV_NVDLA_CDMA_dc.scala 186:70:@4030.4]
  wire [13:0] _T_231; // @[NV_NVDLA_CDMA_dc.scala 188:49:@4031.4]
  wire [8:0] _T_233; // @[NV_NVDLA_CDMA_dc.scala 189:29:@4032.4]
  wire  _T_234; // @[NV_NVDLA_CDMA_dc.scala 190:29:@4033.4]
  wire [12:0] _T_237; // @[NV_NVDLA_CDMA_dc.scala 190:74:@4034.4]
  wire [11:0] _T_238; // @[NV_NVDLA_CDMA_dc.scala 190:74:@4035.4]
  wire [11:0] _T_239; // @[NV_NVDLA_CDMA_dc.scala 190:28:@4036.4]
  wire [26:0] _GEN_157; // @[NV_NVDLA_CDMA_dc.scala 191:38:@4037.4]
  wire [38:0] _T_240; // @[NV_NVDLA_CDMA_dc.scala 191:38:@4037.4]
  wire [13:0] _T_242; // @[NV_NVDLA_CDMA_dc.scala 198:50:@4043.8]
  wire [13:0] _GEN_23; // @[NV_NVDLA_CDMA_dc.scala 194:28:@4039.6]
  wire [12:0] _T_244; // @[NV_NVDLA_CDMA_dc.scala 200:34:@4047.6]
  wire [5:0] _T_246; // @[NV_NVDLA_CDMA_dc.scala 202:41:@4050.6]
  wire [17:0] _T_248; // @[NV_NVDLA_CDMA_dc.scala 203:43:@4052.6]
  wire [16:0] _T_249; // @[NV_NVDLA_CDMA_dc.scala 203:43:@4053.6]
  wire [5:0] _T_251; // @[NV_NVDLA_CDMA_dc.scala 207:42:@4058.6]
  wire [15:0] _GEN_24; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [14:0] _GEN_25; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [13:0] _GEN_26; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [5:0] _GEN_27; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [17:0] _GEN_28; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [12:0] _GEN_29; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [10:0] _GEN_30; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [38:0] _GEN_31; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  reg [13:0] _T_254; // @[NV_NVDLA_CDMA_dc.scala 214:36:@4061.4]
  reg [31:0] _RAND_18;
  reg [13:0] _T_257; // @[NV_NVDLA_CDMA_dc.scala 215:35:@4062.4]
  reg [31:0] _RAND_19;
  reg  _T_260; // @[NV_NVDLA_CDMA_dc.scala 216:39:@4063.4]
  reg [31:0] _RAND_20;
  reg  _T_263; // @[NV_NVDLA_CDMA_dc.scala 217:31:@4064.4]
  reg [31:0] _RAND_21;
  wire  _T_266; // @[NV_NVDLA_CDMA_dc.scala 220:21:@4066.4]
  reg  _T_298; // @[NV_NVDLA_CDMA_dc.scala 253:31:@4107.4]
  reg [31:0] _RAND_22;
  wire  _T_305; // @[NV_NVDLA_CDMA_dc.scala 258:21:@4113.4]
  reg  _T_350; // @[NV_NVDLA_CDMA_dc.scala 292:30:@4148.4]
  reg [31:0] _RAND_23;
  wire  _T_360; // @[NV_NVDLA_CDMA_dc.scala 297:23:@4158.4]
  reg  _T_320; // @[NV_NVDLA_CDMA_dc.scala 282:37:@4138.4]
  reg [31:0] _RAND_24;
  wire  _T_361; // @[NV_NVDLA_CDMA_dc.scala 297:38:@4159.4]
  wire  _T_362; // @[NV_NVDLA_CDMA_dc.scala 297:36:@4160.4]
  reg  _T_323; // @[NV_NVDLA_CDMA_dc.scala 283:37:@4139.4]
  reg [31:0] _RAND_25;
  wire  _T_363; // @[NV_NVDLA_CDMA_dc.scala 297:76:@4161.4]
  wire  _T_364; // @[NV_NVDLA_CDMA_dc.scala 297:74:@4162.4]
  wire  _T_365; // @[NV_NVDLA_CDMA_dc.scala 297:59:@4163.4]
  wire  _T_306; // @[NV_NVDLA_CDMA_dc.scala 258:35:@4114.4]
  wire  _T_267; // @[NV_NVDLA_CDMA_dc.scala 220:35:@4067.4]
  wire  _T_268; // @[NV_NVDLA_CDMA_dc.scala 221:54:@4068.4]
  wire  _T_269; // @[NV_NVDLA_CDMA_dc.scala 221:33:@4069.4]
  wire  _T_270; // @[NV_NVDLA_CDMA_dc.scala 221:71:@4070.4]
  wire [14:0] _T_271; // @[NV_NVDLA_CDMA_dc.scala 222:38:@4071.4]
  wire [14:0] _T_272; // @[NV_NVDLA_CDMA_dc.scala 222:38:@4072.4]
  wire [13:0] _T_273; // @[NV_NVDLA_CDMA_dc.scala 222:38:@4073.4]
  wire [13:0] _GEN_158; // @[NV_NVDLA_CDMA_dc.scala 223:45:@4074.4]
  wire  _T_274; // @[NV_NVDLA_CDMA_dc.scala 223:45:@4074.4]
  wire [13:0] _T_275; // @[NV_NVDLA_CDMA_dc.scala 224:31:@4075.4]
  wire [14:0] _T_277; // @[NV_NVDLA_CDMA_dc.scala 230:48:@4081.8]
  wire [13:0] _T_278; // @[NV_NVDLA_CDMA_dc.scala 230:48:@4082.8]
  wire [13:0] _GEN_33; // @[NV_NVDLA_CDMA_dc.scala 229:26:@4080.6]
  wire [13:0] _GEN_34; // @[NV_NVDLA_CDMA_dc.scala 226:19:@4076.4]
  wire [13:0] _GEN_35; // @[NV_NVDLA_CDMA_dc.scala 233:21:@4085.4]
  wire  _GEN_36; // @[NV_NVDLA_CDMA_dc.scala 233:21:@4085.4]
  wire  _GEN_37; // @[NV_NVDLA_CDMA_dc.scala 244:32:@4099.8]
  wire  _GEN_38; // @[NV_NVDLA_CDMA_dc.scala 241:48:@4095.6]
  wire  _GEN_39; // @[NV_NVDLA_CDMA_dc.scala 237:22:@4090.4]
  reg  _T_286; // @[NV_NVDLA_CDMA_dc.scala 249:32:@4103.4]
  reg [31:0] _RAND_26;
  reg [17:0] _T_289; // @[NV_NVDLA_CDMA_dc.scala 250:37:@4104.4]
  reg [31:0] _RAND_27;
  reg [13:0] _T_292; // @[NV_NVDLA_CDMA_dc.scala 251:35:@4105.4]
  reg [31:0] _RAND_28;
  reg  _T_295; // @[NV_NVDLA_CDMA_dc.scala 252:39:@4106.4]
  reg [31:0] _RAND_29;
  wire [15:0] _GEN_159; // @[NV_NVDLA_CDMA_dc.scala 256:44:@4109.4]
  wire [29:0] _T_301; // @[NV_NVDLA_CDMA_dc.scala 256:44:@4109.4]
  wire [14:0] _T_302; // @[NV_NVDLA_CDMA_dc.scala 256:57:@4110.4]
  wire [17:0] _GEN_160; // @[NV_NVDLA_CDMA_dc.scala 257:41:@4111.4]
  wire [23:0] _T_303; // @[NV_NVDLA_CDMA_dc.scala 257:41:@4111.4]
  wire [17:0] _T_304; // @[NV_NVDLA_CDMA_dc.scala 257:54:@4112.4]
  wire  _T_307; // @[NV_NVDLA_CDMA_dc.scala 259:38:@4116.4]
  wire [14:0] _GEN_40; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  wire [17:0] _GEN_41; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  wire [13:0] _GEN_42; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  wire  _GEN_43; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  wire  _GEN_44; // @[NV_NVDLA_CDMA_dc.scala 275:32:@4132.8]
  wire  _GEN_45; // @[NV_NVDLA_CDMA_dc.scala 272:27:@4128.6]
  wire  _GEN_46; // @[NV_NVDLA_CDMA_dc.scala 268:22:@4124.4]
  reg [13:0] _T_314; // @[NV_NVDLA_CDMA_dc.scala 280:34:@4136.4]
  reg [31:0] _RAND_30;
  reg [13:0] _T_317; // @[NV_NVDLA_CDMA_dc.scala 281:34:@4137.4]
  reg [31:0] _RAND_31;
  reg [17:0] _T_326; // @[NV_NVDLA_CDMA_dc.scala 284:33:@4140.4]
  reg [31:0] _RAND_32;
  reg [17:0] _T_329; // @[NV_NVDLA_CDMA_dc.scala 285:33:@4141.4]
  reg [31:0] _RAND_33;
  reg [17:0] _T_332; // @[NV_NVDLA_CDMA_dc.scala 286:33:@4142.4]
  reg [31:0] _RAND_34;
  reg [17:0] _T_335; // @[NV_NVDLA_CDMA_dc.scala 287:33:@4143.4]
  reg [31:0] _RAND_35;
  reg [17:0] _T_338; // @[NV_NVDLA_CDMA_dc.scala 288:39:@4144.4]
  reg [31:0] _RAND_36;
  reg [17:0] _T_341; // @[NV_NVDLA_CDMA_dc.scala 289:39:@4145.4]
  reg [31:0] _RAND_37;
  reg [13:0] _T_344; // @[NV_NVDLA_CDMA_dc.scala 290:33:@4146.4]
  reg [31:0] _RAND_38;
  wire [17:0] _GEN_161; // @[NV_NVDLA_CDMA_dc.scala 294:44:@4149.4]
  wire [31:0] _T_351; // @[NV_NVDLA_CDMA_dc.scala 294:44:@4149.4]
  wire [17:0] _T_352; // @[NV_NVDLA_CDMA_dc.scala 294:65:@4150.4]
  wire  _T_354; // @[NV_NVDLA_CDMA_dc.scala 295:41:@4152.4]
  wire  _T_356; // @[NV_NVDLA_CDMA_dc.scala 295:56:@4154.4]
  wire  _T_357; // @[NV_NVDLA_CDMA_dc.scala 296:41:@4155.4]
  wire  _T_359; // @[NV_NVDLA_CDMA_dc.scala 296:55:@4157.4]
  wire  _T_366; // @[NV_NVDLA_CDMA_dc.scala 298:38:@4165.4]
  wire  _T_368; // @[NV_NVDLA_CDMA_dc.scala 299:60:@4167.4]
  wire  _T_369; // @[NV_NVDLA_CDMA_dc.scala 299:58:@4168.4]
  wire  _T_371; // @[NV_NVDLA_CDMA_dc.scala 300:58:@4170.4]
  wire [13:0] _GEN_47; // @[NV_NVDLA_CDMA_dc.scala 302:27:@4171.4]
  wire [17:0] _GEN_48; // @[NV_NVDLA_CDMA_dc.scala 302:27:@4171.4]
  wire [13:0] _GEN_49; // @[NV_NVDLA_CDMA_dc.scala 306:27:@4175.4]
  wire [17:0] _GEN_50; // @[NV_NVDLA_CDMA_dc.scala 306:27:@4175.4]
  wire [17:0] _GEN_51; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  wire [17:0] _GEN_52; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  wire [13:0] _GEN_53; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  wire [17:0] _GEN_54; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  wire [17:0] _GEN_55; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  wire [13:0] _GEN_56; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  reg  _T_374; // @[NV_NVDLA_CDMA_dc.scala 322:30:@4189.4]
  reg [31:0] _RAND_39;
  wire  _T_380; // @[NV_NVDLA_CDMA_dc.scala 328:33:@4192.4]
  wire  _T_395; // @[NV_NVDLA_CDMA_dc.scala 334:28:@4203.4]
  reg [2:0] _T_423; // @[NV_NVDLA_CDMA_dc.scala 376:29:@4244.4]
  reg [31:0] _RAND_40;
  wire  _T_488; // @[NV_NVDLA_CDMA_dc.scala 423:39:@4307.4]
  reg [13:0] _T_464; // @[NV_NVDLA_CDMA_dc.scala 412:32:@4291.4]
  reg [31:0] _RAND_41;
  wire [13:0] _T_479; // @[NV_NVDLA_CDMA_dc.scala 421:22:@4299.4]
  wire  _T_480; // @[NV_NVDLA_CDMA_dc.scala 422:42:@4300.4]
  reg [13:0] _T_461; // @[NV_NVDLA_CDMA_dc.scala 411:32:@4290.4]
  reg [31:0] _RAND_42;
  wire  _T_481; // @[NV_NVDLA_CDMA_dc.scala 422:71:@4301.4]
  reg [13:0] _T_458; // @[NV_NVDLA_CDMA_dc.scala 410:32:@4289.4]
  reg [31:0] _RAND_43;
  wire  _T_482; // @[NV_NVDLA_CDMA_dc.scala 422:100:@4302.4]
  reg [13:0] _T_455; // @[NV_NVDLA_CDMA_dc.scala 409:32:@4288.4]
  reg [31:0] _RAND_44;
  wire  _T_483; // @[NV_NVDLA_CDMA_dc.scala 422:129:@4303.4]
  wire [3:0] _T_486; // @[Cat.scala 30:58:@4306.4]
  wire  _T_489; // @[NV_NVDLA_CDMA_dc.scala 423:60:@4308.4]
  wire  _T_490; // @[NV_NVDLA_CDMA_dc.scala 423:64:@4309.4]
  wire  _T_492; // @[NV_NVDLA_CDMA_dc.scala 423:64:@4310.4]
  wire  _T_493; // @[NV_NVDLA_CDMA_dc.scala 423:47:@4311.4]
  wire  _T_495; // @[NV_NVDLA_CDMA_dc.scala 424:39:@4312.4]
  wire [1:0] _T_496; // @[NV_NVDLA_CDMA_dc.scala 424:60:@4313.4]
  wire [1:0] _T_497; // @[NV_NVDLA_CDMA_dc.scala 424:67:@4314.4]
  wire  _T_499; // @[NV_NVDLA_CDMA_dc.scala 424:67:@4315.4]
  wire  _T_500; // @[NV_NVDLA_CDMA_dc.scala 424:47:@4316.4]
  wire  _T_501; // @[NV_NVDLA_CDMA_dc.scala 423:70:@4317.4]
  wire  _T_503; // @[NV_NVDLA_CDMA_dc.scala 425:39:@4318.4]
  wire [2:0] _T_504; // @[NV_NVDLA_CDMA_dc.scala 425:60:@4319.4]
  wire [2:0] _T_505; // @[NV_NVDLA_CDMA_dc.scala 425:67:@4320.4]
  wire  _T_507; // @[NV_NVDLA_CDMA_dc.scala 425:67:@4321.4]
  wire  _T_508; // @[NV_NVDLA_CDMA_dc.scala 425:47:@4322.4]
  wire  _T_509; // @[NV_NVDLA_CDMA_dc.scala 424:73:@4323.4]
  wire  _T_511; // @[NV_NVDLA_CDMA_dc.scala 426:39:@4324.4]
  wire [3:0] _T_513; // @[NV_NVDLA_CDMA_dc.scala 426:67:@4326.4]
  wire  _T_515; // @[NV_NVDLA_CDMA_dc.scala 426:67:@4327.4]
  wire  _T_516; // @[NV_NVDLA_CDMA_dc.scala 426:47:@4328.4]
  wire  _T_517; // @[NV_NVDLA_CDMA_dc.scala 425:73:@4329.4]
  wire  _T_723; // @[NV_NVDLA_CDMA_dc.scala 561:39:@4541.4]
  reg [10:0] _T_420; // @[NV_NVDLA_CDMA_dc.scala 375:29:@4243.4]
  reg [31:0] _RAND_45;
  wire [10:0] _GEN_162; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4271.4]
  wire [11:0] _T_443; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4271.4]
  wire [11:0] _T_444; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4272.4]
  wire [10:0] _T_445; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4273.4]
  wire  _T_446; // @[NV_NVDLA_CDMA_dc.scala 397:34:@4274.4]
  wire  _T_724; // @[NV_NVDLA_CDMA_dc.scala 561:56:@4542.4]
  reg [4:0] _T_411; // @[NV_NVDLA_CDMA_dc.scala 356:32:@4225.4]
  reg [31:0] _RAND_46;
  wire  _T_417; // @[NV_NVDLA_CDMA_dc.scala 372:40:@4241.4]
  wire  _T_725; // @[NV_NVDLA_CDMA_dc.scala 561:72:@4543.4]
  wire  _T_381; // @[NV_NVDLA_CDMA_dc.scala 328:46:@4193.4]
  wire  _T_383; // @[NV_NVDLA_CDMA_dc.scala 328:32:@4194.4]
  wire  _T_384; // @[NV_NVDLA_CDMA_dc.scala 327:32:@4195.4]
  wire  _T_385; // @[NV_NVDLA_CDMA_dc.scala 326:32:@4196.4]
  wire  _T_389; // @[NV_NVDLA_CDMA_dc.scala 332:45:@4198.4]
  wire  _T_391; // @[NV_NVDLA_CDMA_dc.scala 332:32:@4199.4]
  wire  _T_392; // @[NV_NVDLA_CDMA_dc.scala 331:32:@4200.4]
  wire  _T_393; // @[NV_NVDLA_CDMA_dc.scala 330:32:@4201.4]
  wire [1:0] _T_400; // @[NV_NVDLA_CDMA_dc.scala 342:40:@4211.8]
  wire  _T_401; // @[NV_NVDLA_CDMA_dc.scala 342:40:@4212.8]
  wire  _GEN_57; // @[NV_NVDLA_CDMA_dc.scala 341:28:@4210.6]
  wire [1:0] _T_403; // @[NV_NVDLA_CDMA_dc.scala 345:40:@4216.8]
  wire  _T_404; // @[NV_NVDLA_CDMA_dc.scala 345:40:@4217.8]
  wire  _GEN_58; // @[NV_NVDLA_CDMA_dc.scala 344:25:@4215.6]
  wire  _GEN_59; // @[NV_NVDLA_CDMA_dc.scala 336:22:@4205.4]
  wire  _GEN_60; // @[NV_NVDLA_CDMA_dc.scala 336:22:@4205.4]
  wire [5:0] _T_415; // @[NV_NVDLA_CDMA_dc.scala 367:48:@4235.10]
  wire [4:0] _T_416; // @[NV_NVDLA_CDMA_dc.scala 367:48:@4236.10]
  wire [4:0] _GEN_61; // @[NV_NVDLA_CDMA_dc.scala 363:35:@4231.8]
  wire [4:0] _GEN_62; // @[NV_NVDLA_CDMA_dc.scala 362:31:@4230.6]
  wire [4:0] _GEN_63; // @[NV_NVDLA_CDMA_dc.scala 358:19:@4226.4]
  wire  _T_431; // @[NV_NVDLA_CDMA_dc.scala 381:38:@4248.4]
  wire [11:0] _T_432; // @[NV_NVDLA_CDMA_dc.scala 381:84:@4249.4]
  wire [11:0] _T_433; // @[NV_NVDLA_CDMA_dc.scala 381:84:@4250.4]
  wire [10:0] _T_434; // @[NV_NVDLA_CDMA_dc.scala 381:84:@4251.4]
  wire [11:0] _T_435; // @[NV_NVDLA_CDMA_dc.scala 381:97:@4252.4]
  wire [11:0] _T_436; // @[NV_NVDLA_CDMA_dc.scala 381:97:@4253.4]
  wire [10:0] _T_437; // @[NV_NVDLA_CDMA_dc.scala 381:97:@4254.4]
  wire [10:0] _T_438; // @[NV_NVDLA_CDMA_dc.scala 381:28:@4255.4]
  wire [11:0] _T_441; // @[NV_NVDLA_CDMA_dc.scala 392:42:@4265.10]
  wire [10:0] _T_442; // @[NV_NVDLA_CDMA_dc.scala 392:42:@4266.10]
  wire [10:0] _GEN_64; // @[NV_NVDLA_CDMA_dc.scala 388:32:@4261.8]
  wire [10:0] _GEN_65; // @[NV_NVDLA_CDMA_dc.scala 387:28:@4260.6]
  wire [10:0] _GEN_66; // @[NV_NVDLA_CDMA_dc.scala 383:19:@4256.4]
  wire  _T_447; // @[NV_NVDLA_CDMA_dc.scala 398:19:@4276.4]
  wire  _T_448; // @[NV_NVDLA_CDMA_dc.scala 399:28:@4278.6]
  wire [2:0] _T_449; // @[NV_NVDLA_CDMA_dc.scala 403:40:@4283.8]
  wire [2:0] _GEN_67; // @[NV_NVDLA_CDMA_dc.scala 399:42:@4279.6]
  wire [2:0] _GEN_68; // @[NV_NVDLA_CDMA_dc.scala 398:35:@4277.4]
  reg [1:0] _T_452; // @[NV_NVDLA_CDMA_dc.scala 408:30:@4287.4]
  reg [31:0] _RAND_47;
  wire  _T_523; // @[Mux.scala 46:19:@4330.4]
  wire [13:0] _T_524; // @[Mux.scala 46:16:@4331.4]
  wire  _T_525; // @[Mux.scala 46:19:@4332.4]
  wire [13:0] _T_526; // @[Mux.scala 46:16:@4333.4]
  wire  _T_527; // @[Mux.scala 46:19:@4334.4]
  wire [13:0] _T_528; // @[Mux.scala 46:16:@4335.4]
  wire  _T_529; // @[Mux.scala 46:19:@4336.4]
  wire [13:0] _T_530; // @[Mux.scala 46:16:@4337.4]
  wire [14:0] _T_550; // @[NV_NVDLA_CDMA_dc.scala 444:32:@4352.4]
  wire [14:0] _T_551; // @[NV_NVDLA_CDMA_dc.scala 444:32:@4353.4]
  wire [13:0] _T_552; // @[NV_NVDLA_CDMA_dc.scala 444:32:@4354.4]
  wire  _T_554; // @[NV_NVDLA_CDMA_dc.scala 445:51:@4355.4]
  reg [58:0] _T_611; // @[NV_NVDLA_CDMA_dc.scala 486:32:@4419.4]
  reg [63:0] _RAND_48;
  wire [58:0] _GEN_165; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4445.4]
  wire [59:0] _T_637; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4445.4]
  wire [58:0] _T_638; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4446.4]
  wire [2:0] _T_556; // @[NV_NVDLA_CDMA_dc.scala 445:85:@4356.4]
  wire [3:0] _GEN_166; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4357.4]
  wire [4:0] _T_557; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4357.4]
  wire [4:0] _T_558; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4358.4]
  wire [3:0] _T_559; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4359.4]
  wire [3:0] _T_561; // @[NV_NVDLA_CDMA_dc.scala 445:38:@4360.4]
  wire [13:0] _GEN_167; // @[NV_NVDLA_CDMA_dc.scala 446:38:@4361.4]
  wire  _T_562; // @[NV_NVDLA_CDMA_dc.scala 446:38:@4361.4]
  wire [3:0] _T_563; // @[NV_NVDLA_CDMA_dc.scala 446:77:@4362.4]
  wire [3:0] _T_564; // @[NV_NVDLA_CDMA_dc.scala 446:24:@4363.4]
  wire [13:0] _GEN_168; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4338.4]
  wire [14:0] _T_531; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4338.4]
  wire [13:0] _T_532; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4339.4]
  wire  _T_537; // @[NV_NVDLA_CDMA_dc.scala 439:45:@4341.4]
  wire  _T_539; // @[NV_NVDLA_CDMA_dc.scala 440:45:@4342.4]
  wire  _T_541; // @[NV_NVDLA_CDMA_dc.scala 441:45:@4343.4]
  wire  _T_543; // @[Mux.scala 46:16:@4345.4]
  wire  _T_545; // @[Mux.scala 46:16:@4347.4]
  wire  _T_547; // @[Mux.scala 46:16:@4349.4]
  wire  _T_549; // @[Mux.scala 46:16:@4351.4]
  wire [4:0] _T_566; // @[NV_NVDLA_CDMA_dc.scala 447:41:@4365.4]
  wire [4:0] _T_567; // @[NV_NVDLA_CDMA_dc.scala 447:41:@4366.4]
  wire [3:0] _T_568; // @[NV_NVDLA_CDMA_dc.scala 447:41:@4367.4]
  wire  _T_570; // @[NV_NVDLA_CDMA_dc.scala 448:43:@4369.4]
  wire [13:0] _T_572; // @[NV_NVDLA_CDMA_dc.scala 448:30:@4370.4]
  wire [3:0] _T_586; // @[NV_NVDLA_CDMA_dc.scala 453:57:@4380.4]
  wire [3:0] _T_587; // @[NV_NVDLA_CDMA_dc.scala 453:57:@4381.4]
  wire [3:0] _GEN_169; // @[NV_NVDLA_CDMA_dc.scala 453:43:@4382.4]
  wire  _T_588; // @[NV_NVDLA_CDMA_dc.scala 453:43:@4382.4]
  wire  _T_591; // @[NV_NVDLA_CDMA_dc.scala 459:37:@4389.8]
  wire [2:0] _T_594; // @[NV_NVDLA_CDMA_dc.scala 463:44:@4394.10]
  wire [1:0] _T_595; // @[NV_NVDLA_CDMA_dc.scala 463:44:@4395.10]
  wire [1:0] _GEN_69; // @[NV_NVDLA_CDMA_dc.scala 459:54:@4390.8]
  reg  _T_648; // @[NV_NVDLA_CDMA_dc.scala 520:32:@4457.4]
  reg [31:0] _RAND_49;
  wire  _T_681; // @[NV_NVDLA_CDMA_dc.scala 553:37:@4496.4]
  wire  _T_671; // @[NV_NVDLA_CDMA_dc.scala 547:34:@4485.4 NV_NVDLA_CDMA_dc.scala 621:24:@4596.4]
  wire  _T_673; // @[NV_NVDLA_CDMA_dc.scala 548:30:@4486.4 NV_NVDLA_CDMA_dc.scala 581:20:@4556.4]
  wire  _T_674; // @[NV_NVDLA_CDMA_dc.scala 550:40:@4487.4]
  reg  _T_642; // @[NV_NVDLA_CDMA_dc.scala 518:31:@4455.4]
  reg [31:0] _RAND_50;
  wire  _T_675; // @[NV_NVDLA_CDMA_dc.scala 551:39:@4489.4]
  wire  _T_676; // @[NV_NVDLA_CDMA_dc.scala 551:37:@4490.4]
  wire  _T_682; // @[NV_NVDLA_CDMA_dc.scala 553:69:@4497.4]
  wire  _T_683; // @[NV_NVDLA_CDMA_dc.scala 553:53:@4498.4]
  wire [1:0] _GEN_70; // @[NV_NVDLA_CDMA_dc.scala 458:29:@4388.6]
  wire [1:0] _GEN_71; // @[NV_NVDLA_CDMA_dc.scala 454:22:@4384.4]
  wire  _T_686; // @[NV_NVDLA_CDMA_dc.scala 554:89:@4501.4]
  wire  _T_689; // @[NV_NVDLA_CDMA_dc.scala 554:98:@4504.4]
  wire  _T_690; // @[NV_NVDLA_CDMA_dc.scala 554:116:@4505.4]
  wire  _T_691; // @[NV_NVDLA_CDMA_dc.scala 554:73:@4506.4]
  wire  _T_692; // @[NV_NVDLA_CDMA_dc.scala 554:55:@4507.4]
  wire  _T_596; // @[NV_NVDLA_CDMA_dc.scala 469:19:@4400.4]
  wire [13:0] _GEN_72; // @[NV_NVDLA_CDMA_dc.scala 469:38:@4401.4]
  wire  _T_695; // @[NV_NVDLA_CDMA_dc.scala 555:89:@4510.4]
  wire  _T_697; // @[NV_NVDLA_CDMA_dc.scala 555:100:@4512.4]
  wire  _T_698; // @[NV_NVDLA_CDMA_dc.scala 555:98:@4513.4]
  wire  _T_699; // @[NV_NVDLA_CDMA_dc.scala 555:116:@4514.4]
  wire  _T_700; // @[NV_NVDLA_CDMA_dc.scala 555:73:@4515.4]
  wire  _T_701; // @[NV_NVDLA_CDMA_dc.scala 555:55:@4516.4]
  wire  _T_597; // @[NV_NVDLA_CDMA_dc.scala 472:19:@4404.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CDMA_dc.scala 472:38:@4405.4]
  wire  _T_704; // @[NV_NVDLA_CDMA_dc.scala 556:89:@4519.4]
  wire  _T_706; // @[NV_NVDLA_CDMA_dc.scala 556:100:@4521.4]
  wire  _T_707; // @[NV_NVDLA_CDMA_dc.scala 556:98:@4522.4]
  wire  _T_708; // @[NV_NVDLA_CDMA_dc.scala 556:116:@4523.4]
  wire  _T_709; // @[NV_NVDLA_CDMA_dc.scala 556:73:@4524.4]
  wire  _T_710; // @[NV_NVDLA_CDMA_dc.scala 556:55:@4525.4]
  wire  _T_598; // @[NV_NVDLA_CDMA_dc.scala 475:19:@4408.4]
  wire [13:0] _GEN_74; // @[NV_NVDLA_CDMA_dc.scala 475:38:@4409.4]
  wire  _T_713; // @[NV_NVDLA_CDMA_dc.scala 557:89:@4528.4]
  wire  _T_715; // @[NV_NVDLA_CDMA_dc.scala 557:100:@4530.4]
  wire  _T_716; // @[NV_NVDLA_CDMA_dc.scala 557:98:@4531.4]
  wire  _T_717; // @[NV_NVDLA_CDMA_dc.scala 557:116:@4532.4]
  wire  _T_718; // @[NV_NVDLA_CDMA_dc.scala 557:73:@4533.4]
  wire  _T_719; // @[NV_NVDLA_CDMA_dc.scala 557:55:@4534.4]
  wire  _T_599; // @[NV_NVDLA_CDMA_dc.scala 478:19:@4412.4]
  wire [13:0] _GEN_75; // @[NV_NVDLA_CDMA_dc.scala 478:38:@4413.4]
  reg [58:0] _T_602; // @[NV_NVDLA_CDMA_dc.scala 483:38:@4416.4]
  reg [63:0] _RAND_51;
  reg [58:0] _T_605; // @[NV_NVDLA_CDMA_dc.scala 484:38:@4417.4]
  reg [63:0] _RAND_52;
  reg [58:0] _T_608; // @[NV_NVDLA_CDMA_dc.scala 485:35:@4418.4]
  reg [63:0] _RAND_53;
  wire [58:0] _T_612; // @[Cat.scala 30:58:@4420.4]
  wire [58:0] _GEN_170; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4421.4]
  wire [59:0] _T_613; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4421.4]
  wire [58:0] _T_614; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4422.4]
  wire [58:0] _GEN_171; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4423.4]
  wire [59:0] _T_615; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4423.4]
  wire [58:0] _T_616; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4424.4]
  wire [27:0] _GEN_172; // @[NV_NVDLA_CDMA_dc.scala 491:54:@4425.4]
  wire [27:0] _T_617; // @[NV_NVDLA_CDMA_dc.scala 491:54:@4425.4]
  wire [58:0] _GEN_173; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4426.4]
  wire [59:0] _T_618; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4426.4]
  wire [58:0] _T_619; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4427.4]
  wire [58:0] _GEN_174; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4428.4]
  wire [59:0] _T_620; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4428.4]
  wire [58:0] _T_621; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4429.4]
  wire [58:0] _T_622; // @[NV_NVDLA_CDMA_dc.scala 494:36:@4430.4]
  wire [58:0] _T_623; // @[NV_NVDLA_CDMA_dc.scala 496:36:@4431.4]
  wire [58:0] _T_624; // @[NV_NVDLA_CDMA_dc.scala 495:36:@4432.4]
  wire  _T_625; // @[NV_NVDLA_CDMA_dc.scala 499:48:@4433.4]
  wire [58:0] _T_626; // @[NV_NVDLA_CDMA_dc.scala 500:33:@4434.4]
  wire [58:0] _T_627; // @[NV_NVDLA_CDMA_dc.scala 499:33:@4435.4]
  wire [58:0] _T_628; // @[NV_NVDLA_CDMA_dc.scala 498:33:@4436.4]
  wire  _T_629; // @[NV_NVDLA_CDMA_dc.scala 503:46:@4437.4]
  wire  _T_630; // @[NV_NVDLA_CDMA_dc.scala 503:62:@4438.4]
  wire [58:0] _T_632; // @[NV_NVDLA_CDMA_dc.scala 506:30:@4440.4]
  wire [58:0] _T_633; // @[NV_NVDLA_CDMA_dc.scala 505:30:@4441.4]
  wire [58:0] _T_634; // @[NV_NVDLA_CDMA_dc.scala 504:30:@4442.4]
  wire [58:0] _T_635; // @[NV_NVDLA_CDMA_dc.scala 503:30:@4443.4]
  wire [58:0] _T_636; // @[NV_NVDLA_CDMA_dc.scala 502:30:@4444.4]
  wire  _T_639; // @[NV_NVDLA_CDMA_dc.scala 510:27:@4448.4]
  wire [58:0] _GEN_76; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  wire [58:0] _GEN_77; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  wire [58:0] _GEN_78; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  wire [58:0] _GEN_79; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  reg [58:0] _T_645; // @[NV_NVDLA_CDMA_dc.scala 519:30:@4456.4]
  reg [63:0] _RAND_54;
  reg [3:0] _T_651; // @[NV_NVDLA_CDMA_dc.scala 521:30:@4458.4]
  reg [31:0] _RAND_55;
  reg [2:0] _T_654; // @[NV_NVDLA_CDMA_dc.scala 522:34:@4459.4]
  reg [31:0] _RAND_56;
  reg [1:0] _T_657; // @[NV_NVDLA_CDMA_dc.scala 523:32:@4460.4]
  reg [31:0] _RAND_57;
  wire  _T_662; // @[NV_NVDLA_CDMA_dc.scala 527:35:@4463.4]
  wire  _T_663; // @[NV_NVDLA_CDMA_dc.scala 527:51:@4464.4]
  wire  _T_664; // @[NV_NVDLA_CDMA_dc.scala 527:69:@4465.4]
  wire  _T_665; // @[NV_NVDLA_CDMA_dc.scala 527:67:@4466.4]
  wire  _GEN_80; // @[NV_NVDLA_CDMA_dc.scala 535:28:@4476.8]
  wire  _GEN_81; // @[NV_NVDLA_CDMA_dc.scala 532:28:@4472.6]
  wire  _GEN_82; // @[NV_NVDLA_CDMA_dc.scala 529:22:@4468.4]
  wire  _T_679; // @[NV_NVDLA_CDMA_dc.scala 552:49:@4493.4]
  wire  _T_680; // @[NV_NVDLA_CDMA_dc.scala 552:65:@4494.4]
  wire [58:0] _GEN_83; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  wire [3:0] _GEN_84; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  wire [3:0] _GEN_85; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  wire [1:0] _GEN_86; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  reg  _T_738; // @[NV_NVDLA_CDMA_dc.scala 602:30:@4575.4]
  reg [31:0] _RAND_58;
  wire [15:0] _T_745; // @[Cat.scala 30:58:@4583.4]
  wire [14:0] _T_731; // @[NV_NVDLA_CDMA_dc.scala 572:31:@4547.4 NV_NVDLA_CDMA_dc.scala 607:21:@4584.4]
  wire [63:0] _T_742; // @[Cat.scala 30:58:@4580.4]
  wire  _T_740; // @[NV_NVDLA_CDMA_dc.scala 604:42:@4578.4]
  wire  _T_746; // @[NV_NVDLA_CDMA_dc.scala 609:23:@4585.4]
  reg [3:0] _T_753; // @[NV_NVDLA_CDMA_dc.scala 632:35:@4599.4]
  reg [31:0] _RAND_59;
  wire  _T_755; // @[NV_NVDLA_CDMA_dc.scala 635:40:@4601.4]
  wire [3:0] _T_756; // @[NV_NVDLA_CDMA_dc.scala 636:41:@4602.4]
  wire [1:0] _T_757; // @[NV_NVDLA_CDMA_dc.scala 637:43:@4603.4]
  wire [1:0] _GEN_175; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4605.4]
  wire [2:0] _T_760; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4605.4]
  wire [1:0] _T_761; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4606.4]
  wire [3:0] _GEN_176; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4607.4]
  wire [4:0] _T_762; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4607.4]
  wire [3:0] _T_763; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4608.4]
  wire  _T_764; // @[NV_NVDLA_CDMA_dc.scala 643:55:@4609.4]
  wire [3:0] _T_766; // @[NV_NVDLA_CDMA_dc.scala 643:33:@4610.4]
  wire  _T_768; // @[NV_NVDLA_CDMA_dc.scala 644:43:@4612.4]
  wire  _T_770; // @[NV_NVDLA_CDMA_dc.scala 644:58:@4614.4]
  wire [3:0] _GEN_87; // @[NV_NVDLA_CDMA_dc.scala 646:40:@4618.4]
  reg [5:0] _T_775; // @[NV_NVDLA_CDMA_dc.scala 652:37:@4621.4]
  reg [31:0] _RAND_60;
  reg [5:0] _T_778; // @[NV_NVDLA_CDMA_dc.scala 653:37:@4622.4]
  reg [31:0] _RAND_61;
  reg [5:0] _T_781; // @[NV_NVDLA_CDMA_dc.scala 654:37:@4623.4]
  reg [31:0] _RAND_62;
  reg [5:0] _T_784; // @[NV_NVDLA_CDMA_dc.scala 655:37:@4624.4]
  reg [31:0] _RAND_63;
  wire  _T_786; // @[NV_NVDLA_CDMA_dc.scala 657:57:@4625.4]
  wire  _T_787; // @[NV_NVDLA_CDMA_dc.scala 657:39:@4626.4]
  wire  _T_789; // @[NV_NVDLA_CDMA_dc.scala 658:57:@4627.4]
  wire  _T_790; // @[NV_NVDLA_CDMA_dc.scala 658:39:@4628.4]
  wire  _T_792; // @[NV_NVDLA_CDMA_dc.scala 659:57:@4629.4]
  wire  _T_793; // @[NV_NVDLA_CDMA_dc.scala 659:39:@4630.4]
  wire  _T_795; // @[NV_NVDLA_CDMA_dc.scala 660:57:@4631.4]
  wire  _T_796; // @[NV_NVDLA_CDMA_dc.scala 660:39:@4632.4]
  wire  _T_799; // @[NV_NVDLA_CDMA_dc.scala 661:64:@4635.4]
  wire  _T_800; // @[NV_NVDLA_CDMA_dc.scala 661:77:@4636.4]
  wire  _T_804; // @[NV_NVDLA_CDMA_dc.scala 662:77:@4640.4]
  wire  _T_808; // @[NV_NVDLA_CDMA_dc.scala 663:77:@4644.4]
  wire  _T_812; // @[NV_NVDLA_CDMA_dc.scala 664:77:@4648.4]
  wire [5:0] _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4654.8]
  wire [6:0] _T_814; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4654.8]
  wire [5:0] _T_815; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4655.8]
  wire [5:0] _GEN_88; // @[NV_NVDLA_CDMA_dc.scala 670:37:@4653.6]
  wire [6:0] _T_816; // @[NV_NVDLA_CDMA_dc.scala 674:54:@4659.8]
  wire [5:0] _T_817; // @[NV_NVDLA_CDMA_dc.scala 674:54:@4660.8]
  wire [5:0] _GEN_89; // @[NV_NVDLA_CDMA_dc.scala 673:37:@4658.6]
  wire [6:0] _T_818; // @[NV_NVDLA_CDMA_dc.scala 677:54:@4664.8]
  wire [5:0] _T_819; // @[NV_NVDLA_CDMA_dc.scala 677:54:@4665.8]
  wire [5:0] _GEN_90; // @[NV_NVDLA_CDMA_dc.scala 676:37:@4663.6]
  wire [6:0] _T_820; // @[NV_NVDLA_CDMA_dc.scala 680:54:@4669.8]
  wire [5:0] _T_821; // @[NV_NVDLA_CDMA_dc.scala 680:54:@4670.8]
  wire [5:0] _GEN_91; // @[NV_NVDLA_CDMA_dc.scala 679:37:@4668.6]
  wire [5:0] _GEN_92; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  wire [5:0] _GEN_93; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  wire [5:0] _GEN_94; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  wire [5:0] _GEN_95; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  wire  _T_823; // @[NV_NVDLA_CDMA_dc.scala 685:66:@4674.4]
  wire [4:0] _T_824; // @[NV_NVDLA_CDMA_dc.scala 685:89:@4675.4]
  wire [7:0] _T_826; // @[Cat.scala 30:58:@4677.4]
  wire  _T_828; // @[NV_NVDLA_CDMA_dc.scala 686:66:@4678.4]
  wire [4:0] _T_829; // @[NV_NVDLA_CDMA_dc.scala 686:89:@4679.4]
  wire [7:0] _T_831; // @[Cat.scala 30:58:@4681.4]
  wire  _T_833; // @[NV_NVDLA_CDMA_dc.scala 687:66:@4682.4]
  wire [4:0] _T_834; // @[NV_NVDLA_CDMA_dc.scala 687:89:@4683.4]
  wire [7:0] _T_836; // @[Cat.scala 30:58:@4685.4]
  wire  _T_838; // @[NV_NVDLA_CDMA_dc.scala 688:66:@4686.4]
  wire [4:0] _T_839; // @[NV_NVDLA_CDMA_dc.scala 688:89:@4687.4]
  wire [7:0] _T_841; // @[Cat.scala 30:58:@4689.4]
  wire  _T_842; // @[NV_NVDLA_CDMA_dc.scala 694:31:@4690.4]
  wire  _T_844; // @[NV_NVDLA_CDMA_dc.scala 694:48:@4692.4]
  wire [7:0] _T_848; // @[Bitwise.scala 72:12:@4694.4]
  wire [7:0] _GEN_181; // @[NV_NVDLA_CDMA_dc.scala 695:41:@4695.4]
  wire [7:0] _T_849; // @[NV_NVDLA_CDMA_dc.scala 695:41:@4695.4]
  wire [7:0] _T_850; // @[NV_NVDLA_CDMA_dc.scala 695:55:@4696.4]
  wire [7:0] _GEN_182; // @[NV_NVDLA_CDMA_dc.scala 696:41:@4699.4]
  wire [7:0] _T_855; // @[NV_NVDLA_CDMA_dc.scala 696:41:@4699.4]
  wire [7:0] _T_856; // @[NV_NVDLA_CDMA_dc.scala 696:55:@4700.4]
  wire [7:0] _T_857; // @[NV_NVDLA_CDMA_dc.scala 695:71:@4701.4]
  wire [7:0] _GEN_183; // @[NV_NVDLA_CDMA_dc.scala 697:41:@4704.4]
  wire [7:0] _T_862; // @[NV_NVDLA_CDMA_dc.scala 697:41:@4704.4]
  wire [7:0] _T_863; // @[NV_NVDLA_CDMA_dc.scala 697:55:@4705.4]
  wire [7:0] _T_864; // @[NV_NVDLA_CDMA_dc.scala 696:71:@4706.4]
  wire [7:0] _GEN_184; // @[NV_NVDLA_CDMA_dc.scala 698:41:@4709.4]
  wire [7:0] _T_869; // @[NV_NVDLA_CDMA_dc.scala 698:41:@4709.4]
  wire [7:0] _T_870; // @[NV_NVDLA_CDMA_dc.scala 698:55:@4710.4]
  reg [4:0] _T_879; // @[NV_NVDLA_CDMA_dc.scala 710:26:@4718.4]
  reg [31:0] _RAND_64;
  wire [1:0] _T_881; // @[NV_NVDLA_CDMA_dc.scala 712:26:@4719.4]
  wire  _T_1007; // @[NV_NVDLA_CDMA_dc.scala 861:10:@4884.4]
  wire  _T_1008; // @[NV_NVDLA_CDMA_dc.scala 861:23:@4885.4]
  wire [2:0] _GEN_116; // @[NV_NVDLA_CDMA_dc.scala 861:36:@4886.4]
  wire [2:0] _T_883; // @[NV_NVDLA_CDMA_dc.scala 713:26:@4720.4]
  wire  _T_1006; // @[NV_NVDLA_CDMA_dc.scala 859:28:@4883.4]
  wire  _GEN_115; // @[NV_NVDLA_CDMA_dc.scala 861:36:@4886.4]
  reg  _T_1017; // @[NV_NVDLA_CDMA_dc.scala 874:32:@4895.4]
  reg [31:0] _RAND_65;
  wire  _T_1018; // @[NV_NVDLA_CDMA_dc.scala 876:43:@4896.4]
  wire  _T_1019; // @[NV_NVDLA_CDMA_dc.scala 876:41:@4897.4]
  wire  _T_885; // @[NV_NVDLA_CDMA_dc.scala 719:37:@4725.6]
  wire [4:0] _GEN_185; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4727.8]
  wire [5:0] _T_886; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4727.8]
  wire [4:0] _T_887; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4728.8]
  wire [4:0] _GEN_186; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4729.8]
  wire [5:0] _T_888; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4729.8]
  wire [5:0] _T_889; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4730.8]
  wire [4:0] _T_890; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4731.8]
  wire [4:0] _GEN_96; // @[NV_NVDLA_CDMA_dc.scala 719:62:@4726.6]
  wire [4:0] _GEN_97; // @[NV_NVDLA_CDMA_dc.scala 715:19:@4721.4]
  reg [12:0] _T_896; // @[NV_NVDLA_CDMA_dc.scala 729:32:@4736.4]
  reg [31:0] _RAND_66;
  wire [13:0] _GEN_187; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4738.4]
  wire [14:0] _T_899; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4738.4]
  wire [13:0] _T_900; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4739.4]
  wire [14:0] _T_901; // @[NV_NVDLA_CDMA_dc.scala 733:69:@4740.4]
  wire [14:0] _T_902; // @[NV_NVDLA_CDMA_dc.scala 733:69:@4741.4]
  wire [13:0] _T_903; // @[NV_NVDLA_CDMA_dc.scala 733:69:@4742.4]
  wire [13:0] _T_904; // @[NV_NVDLA_CDMA_dc.scala 733:31:@4743.4]
  wire [13:0] _GEN_188; // @[NV_NVDLA_CDMA_dc.scala 734:48:@4744.4]
  wire  _T_905; // @[NV_NVDLA_CDMA_dc.scala 734:48:@4744.4]
  wire [12:0] _T_906; // @[NV_NVDLA_CDMA_dc.scala 734:96:@4745.4]
  wire [12:0] _T_907; // @[NV_NVDLA_CDMA_dc.scala 734:30:@4746.4]
  wire  _T_908; // @[NV_NVDLA_CDMA_dc.scala 735:47:@4747.4]
  reg [15:0] _T_973; // @[NV_NVDLA_CDMA_dc.scala 816:28:@4840.4]
  reg [31:0] _RAND_67;
  wire [15:0] _GEN_189; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4859.4]
  wire [16:0] _T_985; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4859.4]
  wire [16:0] _T_986; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4860.4]
  wire [15:0] _T_987; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4861.4]
  wire  _T_988; // @[NV_NVDLA_CDMA_dc.scala 835:32:@4862.4]
  wire  _T_1001; // @[NV_NVDLA_CDMA_dc.scala 850:34:@4875.4]
  reg [11:0] _T_956; // @[NV_NVDLA_CDMA_dc.scala 797:28:@4818.4]
  reg [31:0] _RAND_68;
  wire [13:0] _T_967; // @[NV_NVDLA_CDMA_dc.scala 813:49:@4835.4]
  wire [13:0] _T_968; // @[NV_NVDLA_CDMA_dc.scala 813:49:@4836.4]
  wire [12:0] _T_969; // @[NV_NVDLA_CDMA_dc.scala 813:49:@4837.4]
  wire [12:0] _GEN_190; // @[NV_NVDLA_CDMA_dc.scala 813:32:@4838.4]
  wire  _T_970; // @[NV_NVDLA_CDMA_dc.scala 813:32:@4838.4]
  wire  _T_1002; // @[NV_NVDLA_CDMA_dc.scala 851:35:@4877.4]
  reg [10:0] _T_927; // @[NV_NVDLA_CDMA_dc.scala 768:29:@4781.4]
  reg [31:0] _RAND_69;
  reg [2:0] _T_930; // @[NV_NVDLA_CDMA_dc.scala 769:29:@4782.4]
  reg [31:0] _RAND_70;
  wire [10:0] _GEN_191; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4795.4]
  wire [11:0] _T_945; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4795.4]
  wire [11:0] _T_946; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4796.4]
  wire [10:0] _T_947; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4797.4]
  wire  _T_948; // @[NV_NVDLA_CDMA_dc.scala 778:33:@4798.4]
  wire  _T_1003; // @[NV_NVDLA_CDMA_dc.scala 852:39:@4879.4]
  reg [4:0] _T_916; // @[NV_NVDLA_CDMA_dc.scala 751:32:@4764.4]
  reg [31:0] _RAND_71;
  wire  _T_917; // @[NV_NVDLA_CDMA_dc.scala 752:43:@4765.4]
  wire  _T_1004; // @[NV_NVDLA_CDMA_dc.scala 853:42:@4881.4]
  wire [13:0] _GEN_98; // @[NV_NVDLA_CDMA_dc.scala 742:31:@4756.6]
  wire  _T_913; // @[NV_NVDLA_CDMA_dc.scala 745:23:@4759.6]
  wire [12:0] _GEN_99; // @[NV_NVDLA_CDMA_dc.scala 745:42:@4760.6]
  wire [13:0] _GEN_100; // @[NV_NVDLA_CDMA_dc.scala 738:19:@4752.4]
  wire [12:0] _GEN_101; // @[NV_NVDLA_CDMA_dc.scala 738:19:@4752.4]
  wire [5:0] _T_923; // @[NV_NVDLA_CDMA_dc.scala 763:44:@4776.10]
  wire [4:0] _T_924; // @[NV_NVDLA_CDMA_dc.scala 763:44:@4777.10]
  wire [4:0] _GEN_102; // @[NV_NVDLA_CDMA_dc.scala 759:31:@4772.8]
  wire [4:0] _GEN_103; // @[NV_NVDLA_CDMA_dc.scala 758:32:@4771.6]
  wire [4:0] _GEN_104; // @[NV_NVDLA_CDMA_dc.scala 755:19:@4767.4]
  wire [11:0] _T_935; // @[NV_NVDLA_CDMA_dc.scala 774:37:@4785.4]
  wire [10:0] _T_936; // @[NV_NVDLA_CDMA_dc.scala 774:37:@4786.4]
  wire  _T_937; // @[NV_NVDLA_CDMA_dc.scala 775:38:@4787.4]
  wire [11:0] _T_938; // @[NV_NVDLA_CDMA_dc.scala 775:84:@4788.4]
  wire [11:0] _T_939; // @[NV_NVDLA_CDMA_dc.scala 775:84:@4789.4]
  wire [10:0] _T_940; // @[NV_NVDLA_CDMA_dc.scala 775:84:@4790.4]
  wire [10:0] _T_941; // @[NV_NVDLA_CDMA_dc.scala 775:28:@4791.4]
  wire  _T_942; // @[NV_NVDLA_CDMA_dc.scala 776:42:@4792.4]
  wire [2:0] _T_943; // @[NV_NVDLA_CDMA_dc.scala 776:83:@4793.4]
  wire [2:0] _T_944; // @[NV_NVDLA_CDMA_dc.scala 776:27:@4794.4]
  wire [10:0] _GEN_105; // @[NV_NVDLA_CDMA_dc.scala 784:28:@4805.8]
  wire [10:0] _GEN_106; // @[NV_NVDLA_CDMA_dc.scala 783:29:@4804.6]
  wire [10:0] _GEN_107; // @[NV_NVDLA_CDMA_dc.scala 780:19:@4800.4]
  wire  _T_953; // @[NV_NVDLA_CDMA_dc.scala 792:19:@4814.4]
  wire [2:0] _GEN_108; // @[NV_NVDLA_CDMA_dc.scala 792:35:@4815.4]
  wire [12:0] _T_964; // @[NV_NVDLA_CDMA_dc.scala 809:36:@4830.10]
  wire [11:0] _T_965; // @[NV_NVDLA_CDMA_dc.scala 809:36:@4831.10]
  wire [11:0] _GEN_109; // @[NV_NVDLA_CDMA_dc.scala 805:27:@4826.8]
  wire [11:0] _GEN_110; // @[NV_NVDLA_CDMA_dc.scala 804:28:@4825.6]
  wire [11:0] _GEN_111; // @[NV_NVDLA_CDMA_dc.scala 801:19:@4821.4]
  wire [15:0] _GEN_194; // @[NV_NVDLA_CDMA_dc.scala 820:34:@4844.4]
  wire  _T_980; // @[NV_NVDLA_CDMA_dc.scala 820:34:@4844.4]
  wire [16:0] _T_983; // @[NV_NVDLA_CDMA_dc.scala 830:36:@4854.10]
  wire [15:0] _T_984; // @[NV_NVDLA_CDMA_dc.scala 830:36:@4855.10]
  wire [15:0] _GEN_112; // @[NV_NVDLA_CDMA_dc.scala 826:27:@4850.8]
  wire [15:0] _GEN_113; // @[NV_NVDLA_CDMA_dc.scala 825:28:@4849.6]
  wire [15:0] _GEN_114; // @[NV_NVDLA_CDMA_dc.scala 822:19:@4845.4]
  wire  _T_992; // @[NV_NVDLA_CDMA_dc.scala 839:39:@4865.4]
  wire  _T_993; // @[NV_NVDLA_CDMA_dc.scala 839:26:@4866.4]
  wire  _T_994; // @[NV_NVDLA_CDMA_dc.scala 839:48:@4867.4]
  wire  _T_995; // @[NV_NVDLA_CDMA_dc.scala 841:55:@4868.4]
  wire  _T_997; // @[NV_NVDLA_CDMA_dc.scala 840:40:@4870.4]
  reg [5:0] _T_1014; // @[NV_NVDLA_CDMA_dc.scala 873:37:@4894.4]
  reg [31:0] _RAND_72;
  wire  _T_1023; // @[NV_NVDLA_CDMA_dc.scala 882:29:@4903.8]
  wire  _GEN_117; // @[NV_NVDLA_CDMA_dc.scala 882:36:@4904.8]
  wire  _GEN_118; // @[NV_NVDLA_CDMA_dc.scala 881:24:@4902.6]
  wire [5:0] _GEN_196; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4915.8]
  wire [6:0] _T_1026; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4915.8]
  wire [5:0] _T_1027; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4916.8]
  wire [5:0] _GEN_119; // @[NV_NVDLA_CDMA_dc.scala 892:37:@4914.6]
  wire [5:0] _GEN_120; // @[NV_NVDLA_CDMA_dc.scala 878:19:@4899.4]
  wire  _GEN_121; // @[NV_NVDLA_CDMA_dc.scala 878:19:@4899.4]
  wire  _T_1029; // @[NV_NVDLA_CDMA_dc.scala 897:66:@4920.4]
  wire [4:0] _T_1030; // @[NV_NVDLA_CDMA_dc.scala 897:89:@4921.4]
  wire [7:0] _T_1032; // @[Cat.scala 30:58:@4923.4]
  wire  _T_1034; // @[NV_NVDLA_CDMA_dc.scala 901:22:@4925.4]
  wire  _T_1037; // @[NV_NVDLA_CDMA_dc.scala 905:37:@4931.6]
  wire  _T_1038; // @[NV_NVDLA_CDMA_dc.scala 905:49:@4932.6]
  wire  _GEN_122; // @[NV_NVDLA_CDMA_dc.scala 901:33:@4926.4]
  reg  _T_1041; // @[NV_NVDLA_CDMA_dc.scala 909:43:@4935.4]
  reg [31:0] _RAND_73;
  reg [7:0] _T_1044; // @[Reg.scala 19:20:@4938.4]
  reg [31:0] _RAND_74;
  wire [7:0] _GEN_123; // @[Reg.scala 20:19:@4939.4]
  reg [17:0] _T_1047; // @[NV_NVDLA_CDMA_dc.scala 915:32:@4943.4]
  reg [31:0] _RAND_75;
  reg [17:0] _T_1050; // @[NV_NVDLA_CDMA_dc.scala 916:35:@4944.4]
  reg [31:0] _RAND_76;
  reg [17:0] _T_1053; // @[NV_NVDLA_CDMA_dc.scala 917:31:@4945.4]
  reg [31:0] _RAND_77;
  wire  _T_1064; // @[NV_NVDLA_CDMA_dc.scala 922:86:@4952.4]
  wire  _T_1077; // @[NV_NVDLA_CDMA_dc.scala 933:71:@4965.4]
  wire  _T_1078; // @[NV_NVDLA_CDMA_dc.scala 933:60:@4966.4]
  wire  _T_1079; // @[NV_NVDLA_CDMA_dc.scala 933:58:@4967.4]
  wire  _T_1065; // @[NV_NVDLA_CDMA_dc.scala 922:75:@4953.4]
  wire  _T_1068; // @[NV_NVDLA_CDMA_dc.scala 922:91:@4956.4]
  wire [17:0] _GEN_197; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4958.4]
  wire [18:0] _T_1071; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4958.4]
  wire [17:0] _T_1072; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4959.4]
  wire [17:0] _T_1073; // @[NV_NVDLA_CDMA_dc.scala 931:34:@4960.4]
  wire  _T_1080; // @[NV_NVDLA_CDMA_dc.scala 936:40:@4969.4]
  wire [18:0] _T_1082; // @[NV_NVDLA_CDMA_dc.scala 936:96:@4970.4]
  wire [17:0] _T_1083; // @[NV_NVDLA_CDMA_dc.scala 936:96:@4971.4]
  wire [17:0] _T_1084; // @[NV_NVDLA_CDMA_dc.scala 936:30:@4972.4]
  wire [17:0] _T_1074; // @[NV_NVDLA_CDMA_dc.scala 930:34:@4961.4]
  wire [17:0] _T_1075; // @[NV_NVDLA_CDMA_dc.scala 929:31:@4962.4]
  wire [18:0] _T_1086; // @[NV_NVDLA_CDMA_dc.scala 939:61:@4974.4]
  wire [17:0] _T_1087; // @[NV_NVDLA_CDMA_dc.scala 939:61:@4975.4]
  wire [18:0] _T_1088; // @[NV_NVDLA_CDMA_dc.scala 940:39:@4976.4]
  wire [17:0] _T_1089; // @[NV_NVDLA_CDMA_dc.scala 940:39:@4977.4]
  wire [17:0] _T_1090; // @[NV_NVDLA_CDMA_dc.scala 939:29:@4978.4]
  wire [17:0] _T_1091; // @[NV_NVDLA_CDMA_dc.scala 938:29:@4979.4]
  wire [17:0] _T_1092; // @[NV_NVDLA_CDMA_dc.scala 937:29:@4980.4]
  reg [14:0] _T_1095; // @[NV_NVDLA_CDMA_dc.scala 941:27:@4981.4]
  reg [31:0] _RAND_78;
  reg [17:0] _T_1098; // @[NV_NVDLA_CDMA_dc.scala 942:35:@4982.4]
  reg [31:0] _RAND_79;
  reg  _T_1101; // @[NV_NVDLA_CDMA_dc.scala 943:29:@4983.4]
  reg [31:0] _RAND_80;
  wire [14:0] _T_1103; // @[NV_NVDLA_CDMA_dc.scala 946:56:@4985.4]
  wire [14:0] _T_1104; // @[NV_NVDLA_CDMA_dc.scala 947:37:@4986.4]
  wire [14:0] _T_1105; // @[NV_NVDLA_CDMA_dc.scala 946:31:@4987.4]
  wire [18:0] _T_1107; // @[NV_NVDLA_CDMA_dc.scala 948:53:@4989.4]
  wire [17:0] _T_1108; // @[NV_NVDLA_CDMA_dc.scala 948:53:@4990.4]
  wire [17:0] _GEN_198; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4991.4]
  wire [18:0] _T_1109; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4991.4]
  wire [17:0] _T_1110; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4992.4]
  wire [17:0] _GEN_199; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4993.4]
  wire [18:0] _T_1111; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4993.4]
  wire [17:0] _T_1112; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4994.4]
  wire [14:0] _T_1114; // @[Cat.scala 30:58:@4995.4]
  wire [17:0] _GEN_200; // @[NV_NVDLA_CDMA_dc.scala 949:41:@4996.4]
  wire  _T_1115; // @[NV_NVDLA_CDMA_dc.scala 949:41:@4996.4]
  wire  _T_1116; // @[NV_NVDLA_CDMA_dc.scala 950:26:@4997.4]
  wire [14:0] _T_1117; // @[NV_NVDLA_CDMA_dc.scala 950:57:@4998.4]
  wire [18:0] _T_1120; // @[NV_NVDLA_CDMA_dc.scala 951:35:@5000.4]
  wire [18:0] _T_1121; // @[NV_NVDLA_CDMA_dc.scala 951:35:@5001.4]
  wire [17:0] _T_1122; // @[NV_NVDLA_CDMA_dc.scala 951:35:@5002.4]
  wire [17:0] _T_1123; // @[NV_NVDLA_CDMA_dc.scala 950:25:@5003.4]
  wire [14:0] _GEN_124; // @[NV_NVDLA_CDMA_dc.scala 954:27:@5005.4]
  wire [17:0] _GEN_125; // @[NV_NVDLA_CDMA_dc.scala 954:27:@5005.4]
  wire  _T_1127; // @[NV_NVDLA_CDMA_dc.scala 958:19:@5009.4]
  wire [17:0] _GEN_126; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  wire [17:0] _GEN_127; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  wire [17:0] _GEN_128; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  wire [17:0] _T_1193; // @[NV_NVDLA_CDMA_dc.scala 1001:21:@5106.4]
  wire [18:0] _T_1128; // @[NV_NVDLA_CDMA_dc.scala 964:46:@5016.6]
  wire [17:0] _T_1129; // @[NV_NVDLA_CDMA_dc.scala 964:46:@5017.6]
  wire [17:0] _GEN_129; // @[NV_NVDLA_CDMA_dc.scala 963:27:@5015.4]
  reg [16:0] _T_1132; // @[NV_NVDLA_CDMA_dc.scala 968:33:@5021.4]
  reg [31:0] _RAND_81;
  wire [17:0] _GEN_130; // @[NV_NVDLA_CDMA_dc.scala 969:23:@5022.4]
  reg  _T_1135; // @[Reg.scala 19:20:@5025.4]
  reg [31:0] _RAND_82;
  wire  _GEN_131; // @[Reg.scala 20:19:@5026.4]
  wire [11:0] _T_1150; // @[Cat.scala 30:58:@5036.4]
  reg  _T_1153; // @[Reg.scala 19:20:@5037.4]
  reg [31:0] _RAND_83;
  wire  _GEN_132; // @[Reg.scala 20:19:@5038.4]
  reg  _T_1155; // @[Reg.scala 19:20:@5041.4]
  reg [31:0] _RAND_84;
  wire  _GEN_133; // @[Reg.scala 20:19:@5042.4]
  reg  _T_1157; // @[Reg.scala 19:20:@5045.4]
  reg [31:0] _RAND_85;
  wire  _GEN_134; // @[Reg.scala 20:19:@5046.4]
  reg  _T_1161; // @[Reg.scala 19:20:@5050.4]
  reg [31:0] _RAND_86;
  reg  _T_1163; // @[Reg.scala 19:20:@5054.4]
  reg [31:0] _RAND_87;
  reg  _T_1165; // @[Reg.scala 19:20:@5058.4]
  reg [31:0] _RAND_88;
  reg [16:0] _T_1168; // @[Reg.scala 19:20:@5063.4]
  reg [31:0] _RAND_89;
  wire [16:0] _GEN_138; // @[Reg.scala 20:19:@5064.4]
  reg [16:0] _T_1170; // @[Reg.scala 19:20:@5067.4]
  reg [31:0] _RAND_90;
  wire [16:0] _GEN_139; // @[Reg.scala 20:19:@5068.4]
  reg [16:0] _T_1172; // @[Reg.scala 19:20:@5071.4]
  reg [31:0] _RAND_91;
  wire [16:0] _GEN_140; // @[Reg.scala 20:19:@5072.4]
  reg [255:0] _T_1175; // @[Reg.scala 19:20:@5076.4]
  reg [255:0] _RAND_92;
  wire [255:0] _GEN_141; // @[Reg.scala 20:19:@5077.4]
  reg [255:0] _T_1177; // @[Reg.scala 19:20:@5080.4]
  reg [255:0] _RAND_93;
  wire [255:0] _GEN_142; // @[Reg.scala 20:19:@5081.4]
  reg [255:0] _T_1179; // @[Reg.scala 19:20:@5084.4]
  reg [255:0] _RAND_94;
  wire [255:0] _GEN_143; // @[Reg.scala 20:19:@5085.4]
  reg [11:0] _T_1182; // @[Reg.scala 19:20:@5089.4]
  reg [31:0] _RAND_95;
  wire [11:0] _GEN_144; // @[Reg.scala 20:19:@5090.4]
  reg [11:0] _T_1184; // @[Reg.scala 19:20:@5093.4]
  reg [31:0] _RAND_96;
  wire [11:0] _GEN_145; // @[Reg.scala 20:19:@5094.4]
  reg [11:0] _T_1186; // @[Reg.scala 19:20:@5097.4]
  reg [31:0] _RAND_97;
  wire [11:0] _GEN_146; // @[Reg.scala 20:19:@5098.4]
  reg [14:0] _T_1189; // @[NV_NVDLA_CDMA_dc.scala 998:33:@5102.4]
  reg [31:0] _RAND_98;
  wire [14:0] _T_1190; // @[NV_NVDLA_CDMA_dc.scala 1000:52:@5103.4]
  wire [14:0] _T_1191; // @[NV_NVDLA_CDMA_dc.scala 1000:75:@5104.4]
  wire [14:0] _T_1192; // @[NV_NVDLA_CDMA_dc.scala 1000:24:@5105.4]
  wire  _T_1194; // @[NV_NVDLA_CDMA_dc.scala 1002:35:@5108.4]
  wire [14:0] _T_1196; // @[NV_NVDLA_CDMA_dc.scala 1002:33:@5109.4]
  wire  _T_1197; // @[NV_NVDLA_CDMA_dc.scala 1003:35:@5110.4]
  wire [14:0] _T_1199; // @[NV_NVDLA_CDMA_dc.scala 1003:33:@5111.4]
  wire  _T_1200; // @[NV_NVDLA_CDMA_dc.scala 1005:27:@5112.4]
  wire [15:0] _T_1201; // @[NV_NVDLA_CDMA_dc.scala 1006:42:@5114.6]
  wire [14:0] _T_1202; // @[NV_NVDLA_CDMA_dc.scala 1006:42:@5115.6]
  wire [15:0] _T_1203; // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5116.6]
  wire [15:0] _T_1204; // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5117.6]
  wire [14:0] _T_1205; // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5118.6]
  wire [14:0] _GEN_147; // @[NV_NVDLA_CDMA_dc.scala 1005:57:@5113.4]
  wire [15:0] _T_1206; // @[NV_NVDLA_CDMA_dc.scala 1010:43:@5121.4]
  wire [15:0] _GEN_202; // @[NV_NVDLA_CDMA_dc.scala 1011:51:@5122.4]
  wire  _T_1207; // @[NV_NVDLA_CDMA_dc.scala 1011:51:@5122.4]
  wire [13:0] _T_1208; // @[NV_NVDLA_CDMA_dc.scala 1012:24:@5123.4]
  wire  _T_1210; // @[NV_NVDLA_CDMA_dc.scala 1014:41:@5125.4]
  wire  _T_1211; // @[NV_NVDLA_CDMA_dc.scala 1014:39:@5126.4]
  wire  _T_1212; // @[NV_NVDLA_CDMA_dc.scala 1014:56:@5127.4]
  wire  _T_1214; // @[NV_NVDLA_CDMA_dc.scala 1014:25:@5128.4]
  reg  _T_1218; // @[Reg.scala 19:20:@5130.4]
  reg [31:0] _RAND_99;
  reg  _T_1220; // @[Reg.scala 19:20:@5134.4]
  reg [31:0] _RAND_100;
  reg  _T_1222; // @[Reg.scala 19:20:@5138.4]
  reg [31:0] _RAND_101;
  reg [14:0] _T_1225; // @[Reg.scala 19:20:@5143.4]
  reg [31:0] _RAND_102;
  wire [17:0] _GEN_151; // @[Reg.scala 20:19:@5144.4]
  reg [14:0] _T_1227; // @[Reg.scala 19:20:@5147.4]
  reg [31:0] _RAND_103;
  wire [14:0] _GEN_152; // @[Reg.scala 20:19:@5148.4]
  reg [14:0] _T_1229; // @[Reg.scala 19:20:@5151.4]
  reg [31:0] _RAND_104;
  wire [14:0] _GEN_153; // @[Reg.scala 20:19:@5152.4]
  reg [13:0] _T_1232; // @[Reg.scala 19:20:@5156.4]
  reg [31:0] _RAND_105;
  wire [13:0] _GEN_154; // @[Reg.scala 20:19:@5157.4]
  reg [13:0] _T_1234; // @[Reg.scala 19:20:@5160.4]
  reg [31:0] _RAND_106;
  wire [13:0] _GEN_155; // @[Reg.scala 20:19:@5161.4]
  reg [13:0] _T_1236; // @[Reg.scala 19:20:@5164.4]
  reg [31:0] _RAND_107;
  wire [13:0] _GEN_156; // @[Reg.scala 20:19:@5165.4]
  wire  _T_1237; // @[NV_NVDLA_CDMA_dc.scala 1025:52:@5169.4]
  wire  _T_1238; // @[NV_NVDLA_CDMA_dc.scala 1025:50:@5170.4]
  wire  _T_1239; // @[NV_NVDLA_CDMA_dc.scala 1025:68:@5171.4]
  reg  _T_1242; // @[NV_NVDLA_CDMA_dc.scala 1025:34:@5172.4]
  reg [31:0] _RAND_108;
  wire  _T_1243; // @[NV_NVDLA_CDMA_dc.scala 1026:60:@5174.4]
  reg  _T_1246; // @[NV_NVDLA_CDMA_dc.scala 1026:34:@5175.4]
  reg [31:0] _RAND_109;
  wire  _T_1247; // @[NV_NVDLA_CDMA_dc.scala 1027:51:@5177.4]
  reg  _T_1250; // @[NV_NVDLA_CDMA_dc.scala 1027:34:@5178.4]
  reg [31:0] _RAND_110;
  reg  _T_1257; // @[NV_NVDLA_CDMA_dc.scala 1040:36:@5192.4]
  reg [31:0] _RAND_111;
  wire  _T_1258; // @[NV_NVDLA_CDMA_dc.scala 1041:56:@5194.4]
  reg  _T_1261; // @[NV_NVDLA_CDMA_dc.scala 1041:36:@5195.4]
  reg [31:0] _RAND_112;
  reg  _T_1264; // @[NV_NVDLA_CDMA_dc.scala 1042:36:@5197.4]
  reg [31:0] _RAND_113;
  reg  _T_1268; // @[NV_NVDLA_CDMA_dc.scala 1043:36:@5200.4]
  reg [31:0] _RAND_114;
  wire [8:0] _T_1270; // @[NV_NVDLA_CDMA_dc.scala 1045:41:@5202.4 NV_NVDLA_CDMA_dc.scala 1055:31:@5215.4]
  wire  _T_1272; // @[NV_NVDLA_CDMA_dc.scala 1046:48:@5203.4]
  wire [31:0] _T_1277; // @[NV_NVDLA_CDMA_dc.scala 1058:47:@5216.4]
  wire  _T_1279; // @[NV_NVDLA_CDMA_dc.scala 1058:47:@5217.4]
  wire  _T_1280; // @[NV_NVDLA_CDMA_dc.scala 1058:22:@5218.4]
  wire  _T_1282; // @[NV_NVDLA_CDMA_dc.scala 1058:82:@5219.4]
  NV_soDLA_DMAIF_rdreq NV_soDLA_DMAIF_rdreq ( // @[NV_NVDLA_CDMA_dc.scala 576:41:@4550.4]
    .reset(NV_NVDLA_DMAIF_rdreq_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk),
    .io_dmaif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready),
    .io_dmaif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid),
    .io_dmaif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits),
    .io_mcif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready),
    .io_mcif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid),
    .io_mcif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits),
    .io_cvif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready),
    .io_cvif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid),
    .io_cvif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits),
    .io_reg2dp_src_ram_type(NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type)
  );
  NV_soDLA_DMAIF_rdrsp NV_soDLA_DMAIF_rdrsp ( // @[NV_NVDLA_CDMA_dc.scala 590:41:@4564.4]
    .reset(NV_NVDLA_DMAIF_rdrsp_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk),
    .io_mcif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready),
    .io_mcif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid),
    .io_mcif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits),
    .io_cvif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready),
    .io_cvif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid),
    .io_cvif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits),
    .io_dmaif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready),
    .io_dmaif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid),
    .io_dmaif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits)
  );
  NV_NVDLA_fifo_1 NV_NVDLA_fifo ( // @[NV_NVDLA_CDMA_dc.scala 615:24:@4590.4]
    .clock(NV_NVDLA_fifo_clock),
    .reset(NV_NVDLA_fifo_reset),
    .io_clk(NV_NVDLA_fifo_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_io_wr_pd),
    .io_rd_pvld(NV_NVDLA_fifo_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_io_rd_pd)
  );
  NV_COUNTER_STAGE_histogram NV_COUNTER_STAGE_histogram ( // @[NV_NVDLA_CDMA_dc.scala 1031:21:@5180.4]
    .reset(NV_COUNTER_STAGE_histogram_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_io_rd_stall_inc),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_io_cnt_cur)
  );
  NV_COUNTER_STAGE_histogram_1 NV_COUNTER_STAGE_histogram_1 ( // @[NV_NVDLA_CDMA_dc.scala 1049:23:@5207.4]
    .reset(NV_COUNTER_STAGE_histogram_1_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_1_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc),
    .io_rd_stall_dec(NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_1_io_cnt_cur)
  );
  NV_COUNTER_STAGE_histogram NV_COUNTER_STAGE_histogram_2 ( // @[NV_NVDLA_CDMA_dc.scala 1061:23:@5221.4]
    .reset(NV_COUNTER_STAGE_histogram_2_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_2_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_2_io_cnt_cur)
  );
  assign _T_94 = 2'h0 == _T_91; // @[Conditional.scala 37:30:@3883.4]
  assign _T_128 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CDMA_dc.scala 123:38:@3938.4]
  assign _T_129 = io_reg2dp_op_en & _T_128; // @[NV_NVDLA_CDMA_dc.scala 124:30:@3939.4]
  assign _T_126 = io_reg2dp_datain_format == 1'h0; // @[NV_NVDLA_CDMA_dc.scala 122:47:@3937.4]
  assign _T_130 = _T_129 & _T_126; // @[NV_NVDLA_CDMA_dc.scala 124:38:@3940.4]
  assign _T_123 = _T_116 != io_reg2dp_data_bank; // @[NV_NVDLA_CDMA_dc.scala 120:37:@3933.4]
  assign _T_95 = _T_130 & _T_123; // @[NV_NVDLA_CDMA_dc.scala 94:21:@3885.6]
  assign _T_96 = _T_130 & io_reg2dp_data_reuse; // @[NV_NVDLA_CDMA_dc.scala 95:26:@3890.8]
  assign _T_97 = _T_96 & _T_85; // @[NV_NVDLA_CDMA_dc.scala 95:49:@3891.8]
  assign _T_124 = _T_130 & _T_119; // @[NV_NVDLA_CDMA_dc.scala 121:25:@3935.4]
  assign _T_98 = _T_97 & _T_124; // @[NV_NVDLA_CDMA_dc.scala 95:70:@3892.8]
  assign _GEN_0 = _T_130 ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_dc.scala 96:27:@3897.10]
  assign _GEN_1 = _T_98 ? 2'h3 : _GEN_0; // @[NV_NVDLA_CDMA_dc.scala 95:84:@3893.8]
  assign _GEN_2 = _T_95 ? 2'h1 : _GEN_1; // @[NV_NVDLA_CDMA_dc.scala 94:37:@3886.6]
  assign _T_99 = 2'h1 == _T_91; // @[Conditional.scala 37:30:@3902.6]
  assign _T_155 = ~ _T_151; // @[NV_NVDLA_CDMA_dc.scala 152:41:@3968.4]
  assign _T_156 = _T_154 & _T_155; // @[NV_NVDLA_CDMA_dc.scala 152:39:@3969.4]
  assign _GEN_3 = _T_156 ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_dc.scala 99:32:@3904.8]
  assign _T_100 = 2'h2 == _T_91; // @[Conditional.scala 37:30:@3909.8]
  assign _T_141 = _T_91 == 2'h2; // @[NV_NVDLA_CDMA_dc.scala 139:30:@3957.4]
  assign _T_909 = ~ io_reg2dp_op_en; // @[NV_NVDLA_CDMA_dc.scala 736:20:@4748.4]
  assign _T_910 = _T_893 == _T_201; // @[NV_NVDLA_CDMA_dc.scala 736:54:@4749.4]
  assign _T_911 = _T_909 | _T_910; // @[NV_NVDLA_CDMA_dc.scala 736:37:@4750.4]
  assign _T_120 = _T_141 & _T_911; // @[NV_NVDLA_CDMA_dc.scala 119:30:@3929.4]
  assign _T_121 = _T_108 == 5'h9; // @[NV_NVDLA_CDMA_dc.scala 119:57:@3930.4]
  assign _T_122 = _T_120 & _T_121; // @[NV_NVDLA_CDMA_dc.scala 119:44:@3931.4]
  assign _GEN_4 = _T_122 ? 2'h3 : 2'h0; // @[NV_NVDLA_CDMA_dc.scala 102:27:@3911.10]
  assign _GEN_7 = _T_100 ? _GEN_4 : 2'h0; // @[Conditional.scala 39:67:@3910.8]
  assign _GEN_8 = _T_99 ? _GEN_3 : _GEN_7; // @[Conditional.scala 39:67:@3903.6]
  assign _GEN_9 = _T_94 ? _GEN_2 : _GEN_8; // @[Conditional.scala 40:58:@3884.4]
  assign _T_131 = ~ _T_141; // @[NV_NVDLA_CDMA_dc.scala 126:10:@3942.4]
  assign _T_134 = _T_108 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 130:32:@3948.8]
  assign _T_135 = _T_108 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 130:32:@3949.8]
  assign _GEN_10 = _T_911 ? _T_135 : _T_108; // @[NV_NVDLA_CDMA_dc.scala 129:27:@3947.6]
  assign _GEN_11 = _T_131 ? 5'h0 : _GEN_10; // @[NV_NVDLA_CDMA_dc.scala 126:22:@3943.4]
  assign _T_139 = _T_91 == 2'h0; // @[NV_NVDLA_CDMA_dc.scala 137:27:@3954.4]
  assign _T_138 = _T_130 & _T_139; // @[NV_NVDLA_CDMA_dc.scala 136:26:@3953.4]
  assign _T_143 = _GEN_9 == 2'h2; // @[NV_NVDLA_CDMA_dc.scala 141:37:@3960.4]
  assign _T_145 = _T_131 & _T_143; // @[NV_NVDLA_CDMA_dc.scala 142:40:@3962.4]
  assign _T_157 = io_reg2dp_op_en & _T_139; // @[NV_NVDLA_CDMA_dc.scala 154:26:@3971.4]
  assign _T_158 = _T_130 & io_reg2dp_skip_data_rls; // @[NV_NVDLA_CDMA_dc.scala 157:37:@3975.6]
  assign _GEN_12 = _T_157 ? _T_130 : _T_119; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  assign _GEN_13 = _T_157 ? io_reg2dp_data_bank : _T_116; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  assign _GEN_14 = _T_157 ? _T_158 : _T_85; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  assign _GEN_15 = _T_157 ? io_sc2cdma_dat_pending_req : _T_151; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  assign _GEN_16 = _T_157 ? _T_151 : _T_154; // @[NV_NVDLA_CDMA_dc.scala 154:36:@3972.4]
  assign _T_221 = io_reg2dp_datain_width == 13'h0; // @[NV_NVDLA_CDMA_dc.scala 185:49:@4025.4]
  assign _T_223 = io_reg2dp_datain_height == 13'h0; // @[NV_NVDLA_CDMA_dc.scala 185:85:@4026.4]
  assign _T_224 = _T_221 & _T_223; // @[NV_NVDLA_CDMA_dc.scala 185:58:@4027.4]
  assign _T_225 = _T_224 & io_reg2dp_surf_packed; // @[NV_NVDLA_CDMA_dc.scala 185:94:@4028.4]
  assign _T_226 = io_reg2dp_datain_channel[12:5]; // @[NV_NVDLA_CDMA_dc.scala 186:52:@4029.4]
  assign _T_228 = _T_226 + 8'h1; // @[NV_NVDLA_CDMA_dc.scala 186:70:@4030.4]
  assign _T_231 = io_reg2dp_datain_height + 13'h1; // @[NV_NVDLA_CDMA_dc.scala 188:49:@4031.4]
  assign _T_233 = _T_225 ? 9'h1 : _T_228; // @[NV_NVDLA_CDMA_dc.scala 189:29:@4032.4]
  assign _T_234 = ~ io_reg2dp_line_packed; // @[NV_NVDLA_CDMA_dc.scala 190:29:@4033.4]
  assign _T_237 = io_reg2dp_grains + 12'h1; // @[NV_NVDLA_CDMA_dc.scala 190:74:@4034.4]
  assign _T_238 = io_reg2dp_grains + 12'h1; // @[NV_NVDLA_CDMA_dc.scala 190:74:@4035.4]
  assign _T_239 = _T_234 ? 12'h1 : _T_238; // @[NV_NVDLA_CDMA_dc.scala 190:28:@4036.4]
  assign _GEN_157 = {{15'd0}, _T_239}; // @[NV_NVDLA_CDMA_dc.scala 191:38:@4037.4]
  assign _T_240 = _GEN_157 * io_reg2dp_line_stride; // @[NV_NVDLA_CDMA_dc.scala 191:38:@4037.4]
  assign _T_242 = io_reg2dp_datain_width + 13'h1; // @[NV_NVDLA_CDMA_dc.scala 198:50:@4043.8]
  assign _GEN_23 = _T_225 ? {{5'd0}, _T_228} : _T_242; // @[NV_NVDLA_CDMA_dc.scala 194:28:@4039.6]
  assign _T_244 = _T_225 ? {{5'd0}, _T_226} : io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_dc.scala 200:34:@4047.6]
  assign _T_246 = io_reg2dp_batches + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 202:41:@4050.6]
  assign _T_248 = io_reg2dp_entries + 17'h1; // @[NV_NVDLA_CDMA_dc.scala 203:43:@4052.6]
  assign _T_249 = io_reg2dp_entries + 17'h1; // @[NV_NVDLA_CDMA_dc.scala 203:43:@4053.6]
  assign _T_251 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 207:42:@4058.6]
  assign _GEN_24 = _T_138 ? {{2'd0}, _GEN_23} : _T_195; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_25 = _T_138 ? {{2'd0}, _T_244} : _T_198; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_26 = _T_138 ? _T_231 : _T_201; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_27 = _T_138 ? _T_246 : _T_204; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_28 = _T_138 ? {{1'd0}, _T_249} : _T_207; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_29 = _T_138 ? {{1'd0}, _T_239} : _T_210; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_30 = _T_138 ? {{2'd0}, _T_233} : _T_213; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_31 = _T_138 ? _T_240 : _T_216; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _GEN_32 = _T_138 ? _T_251 : _T_219; // @[NV_NVDLA_CDMA_dc.scala 193:19:@4038.4]
  assign _T_266 = ~ _T_263; // @[NV_NVDLA_CDMA_dc.scala 220:21:@4066.4]
  assign _T_305 = ~ _T_298; // @[NV_NVDLA_CDMA_dc.scala 258:21:@4113.4]
  assign _T_360 = ~ _T_350; // @[NV_NVDLA_CDMA_dc.scala 297:23:@4158.4]
  assign _T_361 = ~ _T_320; // @[NV_NVDLA_CDMA_dc.scala 297:38:@4159.4]
  assign _T_362 = _T_360 & _T_361; // @[NV_NVDLA_CDMA_dc.scala 297:36:@4160.4]
  assign _T_363 = ~ _T_323; // @[NV_NVDLA_CDMA_dc.scala 297:76:@4161.4]
  assign _T_364 = _T_350 & _T_363; // @[NV_NVDLA_CDMA_dc.scala 297:74:@4162.4]
  assign _T_365 = _T_362 | _T_364; // @[NV_NVDLA_CDMA_dc.scala 297:59:@4163.4]
  assign _T_306 = _T_305 | _T_365; // @[NV_NVDLA_CDMA_dc.scala 258:35:@4114.4]
  assign _T_267 = _T_266 | _T_306; // @[NV_NVDLA_CDMA_dc.scala 220:35:@4067.4]
  assign _T_268 = _T_254 != _T_201; // @[NV_NVDLA_CDMA_dc.scala 221:54:@4068.4]
  assign _T_269 = _T_141 & _T_268; // @[NV_NVDLA_CDMA_dc.scala 221:33:@4069.4]
  assign _T_270 = _T_269 & _T_267; // @[NV_NVDLA_CDMA_dc.scala 221:71:@4070.4]
  assign _T_271 = _T_201 - _T_254; // @[NV_NVDLA_CDMA_dc.scala 222:38:@4071.4]
  assign _T_272 = $unsigned(_T_271); // @[NV_NVDLA_CDMA_dc.scala 222:38:@4072.4]
  assign _T_273 = _T_272[13:0]; // @[NV_NVDLA_CDMA_dc.scala 222:38:@4073.4]
  assign _GEN_158 = {{1'd0}, _T_210}; // @[NV_NVDLA_CDMA_dc.scala 223:45:@4074.4]
  assign _T_274 = _T_273 <= _GEN_158; // @[NV_NVDLA_CDMA_dc.scala 223:45:@4074.4]
  assign _T_275 = _T_274 ? _T_273 : {{1'd0}, _T_210}; // @[NV_NVDLA_CDMA_dc.scala 224:31:@4075.4]
  assign _T_277 = _T_254 + _T_275; // @[NV_NVDLA_CDMA_dc.scala 230:48:@4081.8]
  assign _T_278 = _T_254 + _T_275; // @[NV_NVDLA_CDMA_dc.scala 230:48:@4082.8]
  assign _GEN_33 = _T_270 ? _T_278 : _T_254; // @[NV_NVDLA_CDMA_dc.scala 229:26:@4080.6]
  assign _GEN_34 = _T_138 ? 14'h0 : _GEN_33; // @[NV_NVDLA_CDMA_dc.scala 226:19:@4076.4]
  assign _GEN_35 = _T_270 ? _T_275 : _T_257; // @[NV_NVDLA_CDMA_dc.scala 233:21:@4085.4]
  assign _GEN_36 = _T_270 ? _T_274 : _T_260; // @[NV_NVDLA_CDMA_dc.scala 233:21:@4085.4]
  assign _GEN_37 = _T_306 ? 1'h0 : _T_263; // @[NV_NVDLA_CDMA_dc.scala 244:32:@4099.8]
  assign _GEN_38 = _T_268 ? 1'h1 : _GEN_37; // @[NV_NVDLA_CDMA_dc.scala 241:48:@4095.6]
  assign _GEN_39 = _T_131 ? 1'h0 : _GEN_38; // @[NV_NVDLA_CDMA_dc.scala 237:22:@4090.4]
  assign _GEN_159 = {{2'd0}, _T_257}; // @[NV_NVDLA_CDMA_dc.scala 256:44:@4109.4]
  assign _T_301 = _GEN_159 * _T_195; // @[NV_NVDLA_CDMA_dc.scala 256:44:@4109.4]
  assign _T_302 = _T_301[14:0]; // @[NV_NVDLA_CDMA_dc.scala 256:57:@4110.4]
  assign _GEN_160 = {{12'd0}, _T_204}; // @[NV_NVDLA_CDMA_dc.scala 257:41:@4111.4]
  assign _T_303 = _T_207 * _GEN_160; // @[NV_NVDLA_CDMA_dc.scala 257:41:@4111.4]
  assign _T_304 = _T_303[17:0]; // @[NV_NVDLA_CDMA_dc.scala 257:54:@4112.4]
  assign _T_307 = _T_263 & _T_306; // @[NV_NVDLA_CDMA_dc.scala 259:38:@4116.4]
  assign _GEN_40 = _T_307 ? _T_302 : {{14'd0}, _T_286}; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  assign _GEN_41 = _T_307 ? _T_304 : _T_289; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  assign _GEN_42 = _T_307 ? _T_257 : _T_292; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  assign _GEN_43 = _T_307 ? _T_260 : _T_295; // @[NV_NVDLA_CDMA_dc.scala 261:24:@4117.4]
  assign _GEN_44 = _T_365 ? 1'h0 : _T_298; // @[NV_NVDLA_CDMA_dc.scala 275:32:@4132.8]
  assign _GEN_45 = _T_263 ? 1'h1 : _GEN_44; // @[NV_NVDLA_CDMA_dc.scala 272:27:@4128.6]
  assign _GEN_46 = _T_131 ? 1'h0 : _GEN_45; // @[NV_NVDLA_CDMA_dc.scala 268:22:@4124.4]
  assign _GEN_161 = {{4'd0}, _T_292}; // @[NV_NVDLA_CDMA_dc.scala 294:44:@4149.4]
  assign _T_351 = _GEN_161 * _T_289; // @[NV_NVDLA_CDMA_dc.scala 294:44:@4149.4]
  assign _T_352 = _T_351[17:0]; // @[NV_NVDLA_CDMA_dc.scala 294:65:@4150.4]
  assign _T_354 = _T_298 & _T_360; // @[NV_NVDLA_CDMA_dc.scala 295:41:@4152.4]
  assign _T_356 = _T_354 & _T_361; // @[NV_NVDLA_CDMA_dc.scala 295:56:@4154.4]
  assign _T_357 = _T_298 & _T_350; // @[NV_NVDLA_CDMA_dc.scala 296:41:@4155.4]
  assign _T_359 = _T_357 & _T_363; // @[NV_NVDLA_CDMA_dc.scala 296:55:@4157.4]
  assign _T_366 = _T_298 & _T_365; // @[NV_NVDLA_CDMA_dc.scala 298:38:@4165.4]
  assign _T_368 = ~ _T_295; // @[NV_NVDLA_CDMA_dc.scala 299:60:@4167.4]
  assign _T_369 = _T_366 & _T_368; // @[NV_NVDLA_CDMA_dc.scala 299:58:@4168.4]
  assign _T_371 = _T_366 & _T_295; // @[NV_NVDLA_CDMA_dc.scala 300:58:@4170.4]
  assign _GEN_47 = _T_356 ? {{13'd0}, _T_286} : _T_314; // @[NV_NVDLA_CDMA_dc.scala 302:27:@4171.4]
  assign _GEN_48 = _T_356 ? _T_352 : _T_326; // @[NV_NVDLA_CDMA_dc.scala 302:27:@4171.4]
  assign _GEN_49 = _T_359 ? {{13'd0}, _T_286} : _T_317; // @[NV_NVDLA_CDMA_dc.scala 306:27:@4175.4]
  assign _GEN_50 = _T_359 ? _T_352 : _T_329; // @[NV_NVDLA_CDMA_dc.scala 306:27:@4175.4]
  assign _GEN_51 = _T_369 ? _T_352 : _T_332; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  assign _GEN_52 = _T_369 ? _T_289 : _T_338; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  assign _GEN_53 = _T_369 ? _T_292 : _T_344; // @[NV_NVDLA_CDMA_dc.scala 310:29:@4179.4]
  assign _GEN_54 = _T_371 ? _T_352 : _T_335; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  assign _GEN_55 = _T_371 ? _T_289 : _T_341; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  assign _GEN_56 = _T_371 ? _T_292 : _GEN_42; // @[NV_NVDLA_CDMA_dc.scala 315:29:@4184.4]
  assign _T_380 = ~ _T_374; // @[NV_NVDLA_CDMA_dc.scala 328:33:@4192.4]
  assign _T_395 = _T_380 ? _T_320 : _T_323; // @[NV_NVDLA_CDMA_dc.scala 334:28:@4203.4]
  assign _T_488 = _T_423 == 3'h1; // @[NV_NVDLA_CDMA_dc.scala 423:39:@4307.4]
  assign _T_479 = _T_374 ? _T_317 : _T_314; // @[NV_NVDLA_CDMA_dc.scala 421:22:@4299.4]
  assign _T_480 = _T_464 == _T_479; // @[NV_NVDLA_CDMA_dc.scala 422:42:@4300.4]
  assign _T_481 = _T_461 == _T_479; // @[NV_NVDLA_CDMA_dc.scala 422:71:@4301.4]
  assign _T_482 = _T_458 == _T_479; // @[NV_NVDLA_CDMA_dc.scala 422:100:@4302.4]
  assign _T_483 = _T_455 == _T_479; // @[NV_NVDLA_CDMA_dc.scala 422:129:@4303.4]
  assign _T_486 = {_T_480,_T_481,_T_482,_T_483}; // @[Cat.scala 30:58:@4306.4]
  assign _T_489 = _T_486[0]; // @[NV_NVDLA_CDMA_dc.scala 423:60:@4308.4]
  assign _T_490 = ~ _T_489; // @[NV_NVDLA_CDMA_dc.scala 423:64:@4309.4]
  assign _T_492 = _T_490 == 1'h0; // @[NV_NVDLA_CDMA_dc.scala 423:64:@4310.4]
  assign _T_493 = _T_488 & _T_492; // @[NV_NVDLA_CDMA_dc.scala 423:47:@4311.4]
  assign _T_495 = _T_423 == 3'h2; // @[NV_NVDLA_CDMA_dc.scala 424:39:@4312.4]
  assign _T_496 = _T_486[1:0]; // @[NV_NVDLA_CDMA_dc.scala 424:60:@4313.4]
  assign _T_497 = ~ _T_496; // @[NV_NVDLA_CDMA_dc.scala 424:67:@4314.4]
  assign _T_499 = _T_497 == 2'h0; // @[NV_NVDLA_CDMA_dc.scala 424:67:@4315.4]
  assign _T_500 = _T_495 & _T_499; // @[NV_NVDLA_CDMA_dc.scala 424:47:@4316.4]
  assign _T_501 = _T_493 | _T_500; // @[NV_NVDLA_CDMA_dc.scala 423:70:@4317.4]
  assign _T_503 = _T_423 == 3'h3; // @[NV_NVDLA_CDMA_dc.scala 425:39:@4318.4]
  assign _T_504 = _T_486[2:0]; // @[NV_NVDLA_CDMA_dc.scala 425:60:@4319.4]
  assign _T_505 = ~ _T_504; // @[NV_NVDLA_CDMA_dc.scala 425:67:@4320.4]
  assign _T_507 = _T_505 == 3'h0; // @[NV_NVDLA_CDMA_dc.scala 425:67:@4321.4]
  assign _T_508 = _T_503 & _T_507; // @[NV_NVDLA_CDMA_dc.scala 425:47:@4322.4]
  assign _T_509 = _T_501 | _T_508; // @[NV_NVDLA_CDMA_dc.scala 424:73:@4323.4]
  assign _T_511 = _T_423 == 3'h4; // @[NV_NVDLA_CDMA_dc.scala 426:39:@4324.4]
  assign _T_513 = ~ _T_486; // @[NV_NVDLA_CDMA_dc.scala 426:67:@4326.4]
  assign _T_515 = _T_513 == 4'h0; // @[NV_NVDLA_CDMA_dc.scala 426:67:@4327.4]
  assign _T_516 = _T_511 & _T_515; // @[NV_NVDLA_CDMA_dc.scala 426:47:@4328.4]
  assign _T_517 = _T_509 | _T_516; // @[NV_NVDLA_CDMA_dc.scala 425:73:@4329.4]
  assign _T_723 = _T_395 & _T_517; // @[NV_NVDLA_CDMA_dc.scala 561:39:@4541.4]
  assign _GEN_162 = {{8'd0}, _T_423}; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4271.4]
  assign _T_443 = _T_213 - _GEN_162; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4271.4]
  assign _T_444 = $unsigned(_T_443); // @[NV_NVDLA_CDMA_dc.scala 396:41:@4272.4]
  assign _T_445 = _T_444[10:0]; // @[NV_NVDLA_CDMA_dc.scala 396:41:@4273.4]
  assign _T_446 = _T_420 == _T_445; // @[NV_NVDLA_CDMA_dc.scala 397:34:@4274.4]
  assign _T_724 = _T_723 & _T_446; // @[NV_NVDLA_CDMA_dc.scala 561:56:@4542.4]
  assign _T_417 = _T_411 == io_reg2dp_batches; // @[NV_NVDLA_CDMA_dc.scala 372:40:@4241.4]
  assign _T_725 = _T_724 & _T_417; // @[NV_NVDLA_CDMA_dc.scala 561:72:@4543.4]
  assign _T_381 = _T_380 & _T_725; // @[NV_NVDLA_CDMA_dc.scala 328:46:@4193.4]
  assign _T_383 = _T_381 ? 1'h0 : _T_320; // @[NV_NVDLA_CDMA_dc.scala 328:32:@4194.4]
  assign _T_384 = _T_356 ? 1'h1 : _T_383; // @[NV_NVDLA_CDMA_dc.scala 327:32:@4195.4]
  assign _T_385 = _T_131 ? 1'h0 : _T_384; // @[NV_NVDLA_CDMA_dc.scala 326:32:@4196.4]
  assign _T_389 = _T_374 & _T_725; // @[NV_NVDLA_CDMA_dc.scala 332:45:@4198.4]
  assign _T_391 = _T_389 ? 1'h0 : _T_323; // @[NV_NVDLA_CDMA_dc.scala 332:32:@4199.4]
  assign _T_392 = _T_359 ? 1'h1 : _T_391; // @[NV_NVDLA_CDMA_dc.scala 331:32:@4200.4]
  assign _T_393 = _T_131 ? 1'h0 : _T_392; // @[NV_NVDLA_CDMA_dc.scala 330:32:@4201.4]
  assign _T_400 = _T_350 + 1'h1; // @[NV_NVDLA_CDMA_dc.scala 342:40:@4211.8]
  assign _T_401 = _T_350 + 1'h1; // @[NV_NVDLA_CDMA_dc.scala 342:40:@4212.8]
  assign _GEN_57 = _T_366 ? _T_401 : _T_350; // @[NV_NVDLA_CDMA_dc.scala 341:28:@4210.6]
  assign _T_403 = _T_374 + 1'h1; // @[NV_NVDLA_CDMA_dc.scala 345:40:@4216.8]
  assign _T_404 = _T_374 + 1'h1; // @[NV_NVDLA_CDMA_dc.scala 345:40:@4217.8]
  assign _GEN_58 = _T_725 ? _T_404 : _T_374; // @[NV_NVDLA_CDMA_dc.scala 344:25:@4215.6]
  assign _GEN_59 = _T_131 ? 1'h0 : _GEN_57; // @[NV_NVDLA_CDMA_dc.scala 336:22:@4205.4]
  assign _GEN_60 = _T_131 ? 1'h0 : _GEN_58; // @[NV_NVDLA_CDMA_dc.scala 336:22:@4205.4]
  assign _T_415 = _T_411 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 367:48:@4235.10]
  assign _T_416 = _T_411 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 367:48:@4236.10]
  assign _GEN_61 = _T_417 ? 5'h0 : _T_416; // @[NV_NVDLA_CDMA_dc.scala 363:35:@4231.8]
  assign _GEN_62 = _T_724 ? _GEN_61 : _T_411; // @[NV_NVDLA_CDMA_dc.scala 362:31:@4230.6]
  assign _GEN_63 = _T_138 ? 5'h0 : _GEN_62; // @[NV_NVDLA_CDMA_dc.scala 358:19:@4226.4]
  assign _T_431 = _T_138 | _T_446; // @[NV_NVDLA_CDMA_dc.scala 381:38:@4248.4]
  assign _T_432 = _T_213 - _T_420; // @[NV_NVDLA_CDMA_dc.scala 381:84:@4249.4]
  assign _T_433 = $unsigned(_T_432); // @[NV_NVDLA_CDMA_dc.scala 381:84:@4250.4]
  assign _T_434 = _T_433[10:0]; // @[NV_NVDLA_CDMA_dc.scala 381:84:@4251.4]
  assign _T_435 = _T_434 - _GEN_162; // @[NV_NVDLA_CDMA_dc.scala 381:97:@4252.4]
  assign _T_436 = $unsigned(_T_435); // @[NV_NVDLA_CDMA_dc.scala 381:97:@4253.4]
  assign _T_437 = _T_436[10:0]; // @[NV_NVDLA_CDMA_dc.scala 381:97:@4254.4]
  assign _T_438 = _T_431 ? {{2'd0}, _T_233} : _T_437; // @[NV_NVDLA_CDMA_dc.scala 381:28:@4255.4]
  assign _T_441 = _T_420 + _GEN_162; // @[NV_NVDLA_CDMA_dc.scala 392:42:@4265.10]
  assign _T_442 = _T_420 + _GEN_162; // @[NV_NVDLA_CDMA_dc.scala 392:42:@4266.10]
  assign _GEN_64 = _T_446 ? 11'h0 : _T_442; // @[NV_NVDLA_CDMA_dc.scala 388:32:@4261.8]
  assign _GEN_65 = _T_723 ? _GEN_64 : _T_420; // @[NV_NVDLA_CDMA_dc.scala 387:28:@4260.6]
  assign _GEN_66 = _T_138 ? 11'h0 : _GEN_65; // @[NV_NVDLA_CDMA_dc.scala 383:19:@4256.4]
  assign _T_447 = _T_138 | _T_723; // @[NV_NVDLA_CDMA_dc.scala 398:19:@4276.4]
  assign _T_448 = _T_438 > 11'h1; // @[NV_NVDLA_CDMA_dc.scala 399:28:@4278.6]
  assign _T_449 = _T_438[2:0]; // @[NV_NVDLA_CDMA_dc.scala 403:40:@4283.8]
  assign _GEN_67 = _T_448 ? 3'h1 : _T_449; // @[NV_NVDLA_CDMA_dc.scala 399:42:@4279.6]
  assign _GEN_68 = _T_447 ? _GEN_67 : _T_423; // @[NV_NVDLA_CDMA_dc.scala 398:35:@4277.4]
  assign _T_523 = 2'h3 == _T_452; // @[Mux.scala 46:19:@4330.4]
  assign _T_524 = _T_523 ? _T_464 : 14'h0; // @[Mux.scala 46:16:@4331.4]
  assign _T_525 = 2'h2 == _T_452; // @[Mux.scala 46:19:@4332.4]
  assign _T_526 = _T_525 ? _T_461 : _T_524; // @[Mux.scala 46:16:@4333.4]
  assign _T_527 = 2'h1 == _T_452; // @[Mux.scala 46:19:@4334.4]
  assign _T_528 = _T_527 ? _T_458 : _T_526; // @[Mux.scala 46:16:@4335.4]
  assign _T_529 = 2'h0 == _T_452; // @[Mux.scala 46:19:@4336.4]
  assign _T_530 = _T_529 ? _T_455 : _T_528; // @[Mux.scala 46:16:@4337.4]
  assign _T_550 = _T_479 - _T_530; // @[NV_NVDLA_CDMA_dc.scala 444:32:@4352.4]
  assign _T_551 = $unsigned(_T_550); // @[NV_NVDLA_CDMA_dc.scala 444:32:@4353.4]
  assign _T_552 = _T_551[13:0]; // @[NV_NVDLA_CDMA_dc.scala 444:32:@4354.4]
  assign _T_554 = _T_530 == 14'h0; // @[NV_NVDLA_CDMA_dc.scala 445:51:@4355.4]
  assign _GEN_165 = {{45'd0}, _T_530}; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4445.4]
  assign _T_637 = _T_611 + _GEN_165; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4445.4]
  assign _T_638 = _T_611 + _GEN_165; // @[NV_NVDLA_CDMA_dc.scala 508:30:@4446.4]
  assign _T_556 = _T_638[2:0]; // @[NV_NVDLA_CDMA_dc.scala 445:85:@4356.4]
  assign _GEN_166 = {{1'd0}, _T_556}; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4357.4]
  assign _T_557 = 4'h8 - _GEN_166; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4357.4]
  assign _T_558 = $unsigned(_T_557); // @[NV_NVDLA_CDMA_dc.scala 445:76:@4358.4]
  assign _T_559 = _T_558[3:0]; // @[NV_NVDLA_CDMA_dc.scala 445:76:@4359.4]
  assign _T_561 = _T_554 ? _T_559 : 4'h8; // @[NV_NVDLA_CDMA_dc.scala 445:38:@4360.4]
  assign _GEN_167 = {{10'd0}, _T_561}; // @[NV_NVDLA_CDMA_dc.scala 446:38:@4361.4]
  assign _T_562 = _T_552 < _GEN_167; // @[NV_NVDLA_CDMA_dc.scala 446:38:@4361.4]
  assign _T_563 = _T_552[3:0]; // @[NV_NVDLA_CDMA_dc.scala 446:77:@4362.4]
  assign _T_564 = _T_562 ? _T_563 : _T_561; // @[NV_NVDLA_CDMA_dc.scala 446:24:@4363.4]
  assign _GEN_168 = {{10'd0}, _T_564}; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4338.4]
  assign _T_531 = _T_530 + _GEN_168; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4338.4]
  assign _T_532 = _T_530 + _GEN_168; // @[NV_NVDLA_CDMA_dc.scala 434:39:@4339.4]
  assign _T_537 = _T_486[1]; // @[NV_NVDLA_CDMA_dc.scala 439:45:@4341.4]
  assign _T_539 = _T_486[2]; // @[NV_NVDLA_CDMA_dc.scala 440:45:@4342.4]
  assign _T_541 = _T_486[3]; // @[NV_NVDLA_CDMA_dc.scala 441:45:@4343.4]
  assign _T_543 = _T_523 ? _T_541 : 1'h0; // @[Mux.scala 46:16:@4345.4]
  assign _T_545 = _T_525 ? _T_539 : _T_543; // @[Mux.scala 46:16:@4347.4]
  assign _T_547 = _T_527 ? _T_537 : _T_545; // @[Mux.scala 46:16:@4349.4]
  assign _T_549 = _T_529 ? _T_489 : _T_547; // @[Mux.scala 46:16:@4351.4]
  assign _T_566 = _T_564 - 4'h1; // @[NV_NVDLA_CDMA_dc.scala 447:41:@4365.4]
  assign _T_567 = $unsigned(_T_566); // @[NV_NVDLA_CDMA_dc.scala 447:41:@4366.4]
  assign _T_568 = _T_567[3:0]; // @[NV_NVDLA_CDMA_dc.scala 447:41:@4367.4]
  assign _T_570 = _T_131 | _T_517; // @[NV_NVDLA_CDMA_dc.scala 448:43:@4369.4]
  assign _T_572 = _T_570 ? 14'h0 : _T_532; // @[NV_NVDLA_CDMA_dc.scala 448:30:@4370.4]
  assign _T_586 = _T_423 - 3'h1; // @[NV_NVDLA_CDMA_dc.scala 453:57:@4380.4]
  assign _T_587 = $unsigned(_T_586); // @[NV_NVDLA_CDMA_dc.scala 453:57:@4381.4]
  assign _GEN_169 = {{2'd0}, _T_452}; // @[NV_NVDLA_CDMA_dc.scala 453:43:@4382.4]
  assign _T_588 = _GEN_169 == _T_587; // @[NV_NVDLA_CDMA_dc.scala 453:43:@4382.4]
  assign _T_591 = _T_588 | _T_517; // @[NV_NVDLA_CDMA_dc.scala 459:37:@4389.8]
  assign _T_594 = _T_452 + 2'h1; // @[NV_NVDLA_CDMA_dc.scala 463:44:@4394.10]
  assign _T_595 = _T_452 + 2'h1; // @[NV_NVDLA_CDMA_dc.scala 463:44:@4395.10]
  assign _GEN_69 = _T_591 ? 2'h0 : _T_595; // @[NV_NVDLA_CDMA_dc.scala 459:54:@4390.8]
  assign _T_681 = _T_395 & _T_648; // @[NV_NVDLA_CDMA_dc.scala 553:37:@4496.4]
  assign _T_671 = NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_dc.scala 547:34:@4485.4 NV_NVDLA_CDMA_dc.scala 621:24:@4596.4]
  assign _T_673 = NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 548:30:@4486.4 NV_NVDLA_CDMA_dc.scala 581:20:@4556.4]
  assign _T_674 = _T_671 & _T_673; // @[NV_NVDLA_CDMA_dc.scala 550:40:@4487.4]
  assign _T_675 = ~ _T_642; // @[NV_NVDLA_CDMA_dc.scala 551:39:@4489.4]
  assign _T_676 = _T_674 | _T_675; // @[NV_NVDLA_CDMA_dc.scala 551:37:@4490.4]
  assign _T_682 = _T_549 | _T_676; // @[NV_NVDLA_CDMA_dc.scala 553:69:@4497.4]
  assign _T_683 = _T_681 & _T_682; // @[NV_NVDLA_CDMA_dc.scala 553:53:@4498.4]
  assign _GEN_70 = _T_683 ? _GEN_69 : _T_452; // @[NV_NVDLA_CDMA_dc.scala 458:29:@4388.6]
  assign _GEN_71 = _T_131 ? 2'h0 : _GEN_70; // @[NV_NVDLA_CDMA_dc.scala 454:22:@4384.4]
  assign _T_686 = _T_452 == 2'h0; // @[NV_NVDLA_CDMA_dc.scala 554:89:@4501.4]
  assign _T_689 = _T_686 & _T_490; // @[NV_NVDLA_CDMA_dc.scala 554:98:@4504.4]
  assign _T_690 = _T_689 & _T_676; // @[NV_NVDLA_CDMA_dc.scala 554:116:@4505.4]
  assign _T_691 = _T_517 | _T_690; // @[NV_NVDLA_CDMA_dc.scala 554:73:@4506.4]
  assign _T_692 = _T_681 & _T_691; // @[NV_NVDLA_CDMA_dc.scala 554:55:@4507.4]
  assign _T_596 = _T_138 | _T_692; // @[NV_NVDLA_CDMA_dc.scala 469:19:@4400.4]
  assign _GEN_72 = _T_596 ? _T_572 : _T_455; // @[NV_NVDLA_CDMA_dc.scala 469:38:@4401.4]
  assign _T_695 = _T_452 == 2'h1; // @[NV_NVDLA_CDMA_dc.scala 555:89:@4510.4]
  assign _T_697 = ~ _T_537; // @[NV_NVDLA_CDMA_dc.scala 555:100:@4512.4]
  assign _T_698 = _T_695 & _T_697; // @[NV_NVDLA_CDMA_dc.scala 555:98:@4513.4]
  assign _T_699 = _T_698 & _T_676; // @[NV_NVDLA_CDMA_dc.scala 555:116:@4514.4]
  assign _T_700 = _T_517 | _T_699; // @[NV_NVDLA_CDMA_dc.scala 555:73:@4515.4]
  assign _T_701 = _T_681 & _T_700; // @[NV_NVDLA_CDMA_dc.scala 555:55:@4516.4]
  assign _T_597 = _T_138 | _T_701; // @[NV_NVDLA_CDMA_dc.scala 472:19:@4404.4]
  assign _GEN_73 = _T_597 ? _T_572 : _T_458; // @[NV_NVDLA_CDMA_dc.scala 472:38:@4405.4]
  assign _T_704 = _T_452 == 2'h2; // @[NV_NVDLA_CDMA_dc.scala 556:89:@4519.4]
  assign _T_706 = ~ _T_539; // @[NV_NVDLA_CDMA_dc.scala 556:100:@4521.4]
  assign _T_707 = _T_704 & _T_706; // @[NV_NVDLA_CDMA_dc.scala 556:98:@4522.4]
  assign _T_708 = _T_707 & _T_676; // @[NV_NVDLA_CDMA_dc.scala 556:116:@4523.4]
  assign _T_709 = _T_517 | _T_708; // @[NV_NVDLA_CDMA_dc.scala 556:73:@4524.4]
  assign _T_710 = _T_681 & _T_709; // @[NV_NVDLA_CDMA_dc.scala 556:55:@4525.4]
  assign _T_598 = _T_138 | _T_710; // @[NV_NVDLA_CDMA_dc.scala 475:19:@4408.4]
  assign _GEN_74 = _T_598 ? _T_572 : _T_461; // @[NV_NVDLA_CDMA_dc.scala 475:38:@4409.4]
  assign _T_713 = _T_452 == 2'h3; // @[NV_NVDLA_CDMA_dc.scala 557:89:@4528.4]
  assign _T_715 = ~ _T_541; // @[NV_NVDLA_CDMA_dc.scala 557:100:@4530.4]
  assign _T_716 = _T_713 & _T_715; // @[NV_NVDLA_CDMA_dc.scala 557:98:@4531.4]
  assign _T_717 = _T_716 & _T_676; // @[NV_NVDLA_CDMA_dc.scala 557:116:@4532.4]
  assign _T_718 = _T_517 | _T_717; // @[NV_NVDLA_CDMA_dc.scala 557:73:@4533.4]
  assign _T_719 = _T_681 & _T_718; // @[NV_NVDLA_CDMA_dc.scala 557:55:@4534.4]
  assign _T_599 = _T_138 | _T_719; // @[NV_NVDLA_CDMA_dc.scala 478:19:@4412.4]
  assign _GEN_75 = _T_599 ? _T_572 : _T_464; // @[NV_NVDLA_CDMA_dc.scala 478:38:@4413.4]
  assign _T_612 = {io_reg2dp_datain_addr_high_0,io_reg2dp_datain_addr_low_0}; // @[Cat.scala 30:58:@4420.4]
  assign _GEN_170 = {{20'd0}, _T_216}; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4421.4]
  assign _T_613 = _T_602 + _GEN_170; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4421.4]
  assign _T_614 = _T_602 + _GEN_170; // @[NV_NVDLA_CDMA_dc.scala 489:55:@4422.4]
  assign _GEN_171 = {{32'd0}, io_reg2dp_batch_stride}; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4423.4]
  assign _T_615 = _T_605 + _GEN_171; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4423.4]
  assign _T_616 = _T_605 + _GEN_171; // @[NV_NVDLA_CDMA_dc.scala 490:55:@4424.4]
  assign _GEN_172 = {{1'd0}, io_reg2dp_surf_stride}; // @[NV_NVDLA_CDMA_dc.scala 491:54:@4425.4]
  assign _T_617 = _GEN_172 << 1; // @[NV_NVDLA_CDMA_dc.scala 491:54:@4425.4]
  assign _GEN_173 = {{31'd0}, _T_617}; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4426.4]
  assign _T_618 = _T_608 + _GEN_173; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4426.4]
  assign _T_619 = _T_608 + _GEN_173; // @[NV_NVDLA_CDMA_dc.scala 492:49:@4427.4]
  assign _GEN_174 = {{32'd0}, io_reg2dp_surf_stride}; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4428.4]
  assign _T_620 = _T_611 + _GEN_174; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4428.4]
  assign _T_621 = _T_611 + _GEN_174; // @[NV_NVDLA_CDMA_dc.scala 493:43:@4429.4]
  assign _T_622 = _T_145 ? _T_612 : _T_614; // @[NV_NVDLA_CDMA_dc.scala 494:36:@4430.4]
  assign _T_623 = _T_417 ? _T_614 : _T_616; // @[NV_NVDLA_CDMA_dc.scala 496:36:@4431.4]
  assign _T_624 = _T_145 ? _T_612 : _T_623; // @[NV_NVDLA_CDMA_dc.scala 495:36:@4432.4]
  assign _T_625 = _T_446 & _T_417; // @[NV_NVDLA_CDMA_dc.scala 499:48:@4433.4]
  assign _T_626 = _T_446 ? _T_616 : _T_619; // @[NV_NVDLA_CDMA_dc.scala 500:33:@4434.4]
  assign _T_627 = _T_625 ? _T_614 : _T_626; // @[NV_NVDLA_CDMA_dc.scala 499:33:@4435.4]
  assign _T_628 = _T_145 ? _T_612 : _T_627; // @[NV_NVDLA_CDMA_dc.scala 498:33:@4436.4]
  assign _T_629 = _T_517 & _T_446; // @[NV_NVDLA_CDMA_dc.scala 503:46:@4437.4]
  assign _T_630 = _T_629 & _T_417; // @[NV_NVDLA_CDMA_dc.scala 503:62:@4438.4]
  assign _T_632 = _T_588 ? _T_608 : _T_621; // @[NV_NVDLA_CDMA_dc.scala 506:30:@4440.4]
  assign _T_633 = _T_517 ? _T_619 : _T_632; // @[NV_NVDLA_CDMA_dc.scala 505:30:@4441.4]
  assign _T_634 = _T_629 ? _T_616 : _T_633; // @[NV_NVDLA_CDMA_dc.scala 504:30:@4442.4]
  assign _T_635 = _T_630 ? _T_614 : _T_634; // @[NV_NVDLA_CDMA_dc.scala 503:30:@4443.4]
  assign _T_636 = _T_145 ? _T_612 : _T_635; // @[NV_NVDLA_CDMA_dc.scala 502:30:@4444.4]
  assign _T_639 = _T_145 | _T_725; // @[NV_NVDLA_CDMA_dc.scala 510:27:@4448.4]
  assign _GEN_76 = _T_639 ? _T_622 : _T_602; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  assign _GEN_77 = _T_639 ? _T_624 : _T_605; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  assign _GEN_78 = _T_639 ? _T_628 : _T_608; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  assign _GEN_79 = _T_639 ? _T_636 : _T_611; // @[NV_NVDLA_CDMA_dc.scala 510:46:@4449.4]
  assign _T_662 = _T_141 & _T_395; // @[NV_NVDLA_CDMA_dc.scala 527:35:@4463.4]
  assign _T_663 = _T_662 & _T_648; // @[NV_NVDLA_CDMA_dc.scala 527:51:@4464.4]
  assign _T_664 = ~ _T_549; // @[NV_NVDLA_CDMA_dc.scala 527:69:@4465.4]
  assign _T_665 = _T_663 & _T_664; // @[NV_NVDLA_CDMA_dc.scala 527:67:@4466.4]
  assign _GEN_80 = _T_674 ? 1'h0 : _T_642; // @[NV_NVDLA_CDMA_dc.scala 535:28:@4476.8]
  assign _GEN_81 = _T_665 ? 1'h1 : _GEN_80; // @[NV_NVDLA_CDMA_dc.scala 532:28:@4472.6]
  assign _GEN_82 = _T_131 ? 1'h0 : _GEN_81; // @[NV_NVDLA_CDMA_dc.scala 529:22:@4468.4]
  assign _T_679 = _T_681 & _T_664; // @[NV_NVDLA_CDMA_dc.scala 552:49:@4493.4]
  assign _T_680 = _T_679 & _T_676; // @[NV_NVDLA_CDMA_dc.scala 552:65:@4494.4]
  assign _GEN_83 = _T_680 ? _T_638 : _T_645; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  assign _GEN_84 = _T_680 ? _T_564 : _T_651; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  assign _GEN_85 = _T_680 ? _T_568 : {{1'd0}, _T_654}; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  assign _GEN_86 = _T_680 ? _T_452 : _T_657; // @[NV_NVDLA_CDMA_dc.scala 539:21:@4479.4]
  assign _T_745 = {13'h0,_T_654}; // @[Cat.scala 30:58:@4583.4]
  assign _T_731 = _T_745[14:0]; // @[NV_NVDLA_CDMA_dc.scala 572:31:@4547.4 NV_NVDLA_CDMA_dc.scala 607:21:@4584.4]
  assign _T_742 = {_T_645,5'h0}; // @[Cat.scala 30:58:@4580.4]
  assign _T_740 = _T_671 & _T_642; // @[NV_NVDLA_CDMA_dc.scala 604:42:@4578.4]
  assign _T_746 = ~ _T_738; // @[NV_NVDLA_CDMA_dc.scala 609:23:@4585.4]
  assign _T_755 = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits[256]; // @[NV_NVDLA_CDMA_dc.scala 635:40:@4601.4]
  assign _T_756 = NV_NVDLA_fifo_io_rd_pd[3:0]; // @[NV_NVDLA_CDMA_dc.scala 636:41:@4602.4]
  assign _T_757 = NV_NVDLA_fifo_io_rd_pd[5:4]; // @[NV_NVDLA_CDMA_dc.scala 637:43:@4603.4]
  assign _GEN_175 = {{1'd0}, _T_755}; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4605.4]
  assign _T_760 = _GEN_175 + 2'h2; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4605.4]
  assign _T_761 = _GEN_175 + 2'h2; // @[NV_NVDLA_CDMA_dc.scala 639:53:@4606.4]
  assign _GEN_176 = {{2'd0}, _T_761}; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4607.4]
  assign _T_762 = _T_753 + _GEN_176; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4607.4]
  assign _T_763 = _T_753 + _GEN_176; // @[NV_NVDLA_CDMA_dc.scala 641:49:@4608.4]
  assign _T_764 = _T_763 == _T_756; // @[NV_NVDLA_CDMA_dc.scala 643:55:@4609.4]
  assign _T_766 = _T_764 ? 4'h0 : _T_763; // @[NV_NVDLA_CDMA_dc.scala 643:33:@4610.4]
  assign _T_768 = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid & _T_746; // @[NV_NVDLA_CDMA_dc.scala 644:43:@4612.4]
  assign _T_770 = _T_768 & _T_764; // @[NV_NVDLA_CDMA_dc.scala 644:58:@4614.4]
  assign _GEN_87 = _T_768 ? _T_766 : _T_753; // @[NV_NVDLA_CDMA_dc.scala 646:40:@4618.4]
  assign _T_786 = _T_757 == 2'h0; // @[NV_NVDLA_CDMA_dc.scala 657:57:@4625.4]
  assign _T_787 = NV_NVDLA_fifo_io_rd_pvld & _T_786; // @[NV_NVDLA_CDMA_dc.scala 657:39:@4626.4]
  assign _T_789 = _T_757 == 2'h1; // @[NV_NVDLA_CDMA_dc.scala 658:57:@4627.4]
  assign _T_790 = NV_NVDLA_fifo_io_rd_pvld & _T_789; // @[NV_NVDLA_CDMA_dc.scala 658:39:@4628.4]
  assign _T_792 = _T_757 == 2'h2; // @[NV_NVDLA_CDMA_dc.scala 659:57:@4629.4]
  assign _T_793 = NV_NVDLA_fifo_io_rd_pvld & _T_792; // @[NV_NVDLA_CDMA_dc.scala 659:39:@4630.4]
  assign _T_795 = _T_757 == 2'h3; // @[NV_NVDLA_CDMA_dc.scala 660:57:@4631.4]
  assign _T_796 = NV_NVDLA_fifo_io_rd_pvld & _T_795; // @[NV_NVDLA_CDMA_dc.scala 660:39:@4632.4]
  assign _T_799 = _T_768 & _T_141; // @[NV_NVDLA_CDMA_dc.scala 661:64:@4635.4]
  assign _T_800 = _T_799 & _T_787; // @[NV_NVDLA_CDMA_dc.scala 661:77:@4636.4]
  assign _T_804 = _T_799 & _T_790; // @[NV_NVDLA_CDMA_dc.scala 662:77:@4640.4]
  assign _T_808 = _T_799 & _T_793; // @[NV_NVDLA_CDMA_dc.scala 663:77:@4644.4]
  assign _T_812 = _T_799 & _T_796; // @[NV_NVDLA_CDMA_dc.scala 664:77:@4648.4]
  assign _GEN_177 = {{4'd0}, _T_761}; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4654.8]
  assign _T_814 = _T_775 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4654.8]
  assign _T_815 = _T_775 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 671:54:@4655.8]
  assign _GEN_88 = _T_800 ? _T_815 : _T_775; // @[NV_NVDLA_CDMA_dc.scala 670:37:@4653.6]
  assign _T_816 = _T_778 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 674:54:@4659.8]
  assign _T_817 = _T_778 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 674:54:@4660.8]
  assign _GEN_89 = _T_804 ? _T_817 : _T_778; // @[NV_NVDLA_CDMA_dc.scala 673:37:@4658.6]
  assign _T_818 = _T_781 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 677:54:@4664.8]
  assign _T_819 = _T_781 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 677:54:@4665.8]
  assign _GEN_90 = _T_808 ? _T_819 : _T_781; // @[NV_NVDLA_CDMA_dc.scala 676:37:@4663.6]
  assign _T_820 = _T_784 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 680:54:@4669.8]
  assign _T_821 = _T_784 + _GEN_177; // @[NV_NVDLA_CDMA_dc.scala 680:54:@4670.8]
  assign _GEN_91 = _T_812 ? _T_821 : _T_784; // @[NV_NVDLA_CDMA_dc.scala 679:37:@4668.6]
  assign _GEN_92 = _T_138 ? 6'h0 : _GEN_88; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  assign _GEN_93 = _T_138 ? _T_778 : _GEN_89; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  assign _GEN_94 = _T_138 ? _T_781 : _GEN_90; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  assign _GEN_95 = _T_138 ? _T_784 : _GEN_91; // @[NV_NVDLA_CDMA_dc.scala 666:19:@4649.4]
  assign _T_823 = _T_775[0]; // @[NV_NVDLA_CDMA_dc.scala 685:66:@4674.4]
  assign _T_824 = _T_775[5:1]; // @[NV_NVDLA_CDMA_dc.scala 685:89:@4675.4]
  assign _T_826 = {2'h0,_T_823,_T_824}; // @[Cat.scala 30:58:@4677.4]
  assign _T_828 = _T_778[0]; // @[NV_NVDLA_CDMA_dc.scala 686:66:@4678.4]
  assign _T_829 = _T_778[5:1]; // @[NV_NVDLA_CDMA_dc.scala 686:89:@4679.4]
  assign _T_831 = {2'h0,_T_828,_T_829}; // @[Cat.scala 30:58:@4681.4]
  assign _T_833 = _T_781[0]; // @[NV_NVDLA_CDMA_dc.scala 687:66:@4682.4]
  assign _T_834 = _T_781[5:1]; // @[NV_NVDLA_CDMA_dc.scala 687:89:@4683.4]
  assign _T_836 = {2'h0,_T_833,_T_834}; // @[Cat.scala 30:58:@4685.4]
  assign _T_838 = _T_784[0]; // @[NV_NVDLA_CDMA_dc.scala 688:66:@4686.4]
  assign _T_839 = _T_784[5:1]; // @[NV_NVDLA_CDMA_dc.scala 688:89:@4687.4]
  assign _T_841 = {2'h0,_T_838,_T_839}; // @[Cat.scala 30:58:@4689.4]
  assign _T_842 = _T_141 & NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 694:31:@4690.4]
  assign _T_844 = _T_842 & _T_746; // @[NV_NVDLA_CDMA_dc.scala 694:48:@4692.4]
  assign _T_848 = _T_844 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@4694.4]
  assign _GEN_181 = {{7'd0}, _T_787}; // @[NV_NVDLA_CDMA_dc.scala 695:41:@4695.4]
  assign _T_849 = _T_848 & _GEN_181; // @[NV_NVDLA_CDMA_dc.scala 695:41:@4695.4]
  assign _T_850 = _T_849 & _T_826; // @[NV_NVDLA_CDMA_dc.scala 695:55:@4696.4]
  assign _GEN_182 = {{7'd0}, _T_790}; // @[NV_NVDLA_CDMA_dc.scala 696:41:@4699.4]
  assign _T_855 = _T_848 & _GEN_182; // @[NV_NVDLA_CDMA_dc.scala 696:41:@4699.4]
  assign _T_856 = _T_855 & _T_831; // @[NV_NVDLA_CDMA_dc.scala 696:55:@4700.4]
  assign _T_857 = _T_850 | _T_856; // @[NV_NVDLA_CDMA_dc.scala 695:71:@4701.4]
  assign _GEN_183 = {{7'd0}, _T_793}; // @[NV_NVDLA_CDMA_dc.scala 697:41:@4704.4]
  assign _T_862 = _T_848 & _GEN_183; // @[NV_NVDLA_CDMA_dc.scala 697:41:@4704.4]
  assign _T_863 = _T_862 & _T_836; // @[NV_NVDLA_CDMA_dc.scala 697:55:@4705.4]
  assign _T_864 = _T_857 | _T_863; // @[NV_NVDLA_CDMA_dc.scala 696:71:@4706.4]
  assign _GEN_184 = {{7'd0}, _T_796}; // @[NV_NVDLA_CDMA_dc.scala 698:41:@4709.4]
  assign _T_869 = _T_848 & _GEN_184; // @[NV_NVDLA_CDMA_dc.scala 698:41:@4709.4]
  assign _T_870 = _T_869 & _T_841; // @[NV_NVDLA_CDMA_dc.scala 698:55:@4710.4]
  assign _T_881 = _T_800 ? _T_761 : 2'h0; // @[NV_NVDLA_CDMA_dc.scala 712:26:@4719.4]
  assign _T_1007 = ~ _T_911; // @[NV_NVDLA_CDMA_dc.scala 861:10:@4884.4]
  assign _T_1008 = _T_1007 & _T_141; // @[NV_NVDLA_CDMA_dc.scala 861:23:@4885.4]
  assign _GEN_116 = _T_1008 ? 3'h1 : 3'h0; // @[NV_NVDLA_CDMA_dc.scala 861:36:@4886.4]
  assign _T_883 = _T_800 ? _GEN_116 : 3'h0; // @[NV_NVDLA_CDMA_dc.scala 713:26:@4720.4]
  assign _T_1006 = _T_879 != 5'h0; // @[NV_NVDLA_CDMA_dc.scala 859:28:@4883.4]
  assign _GEN_115 = _T_1008 ? _T_1006 : 1'h0; // @[NV_NVDLA_CDMA_dc.scala 861:36:@4886.4]
  assign _T_1018 = ~ _T_1017; // @[NV_NVDLA_CDMA_dc.scala 876:43:@4896.4]
  assign _T_1019 = _GEN_115 & _T_1018; // @[NV_NVDLA_CDMA_dc.scala 876:41:@4897.4]
  assign _T_885 = _T_800 | _T_1019; // @[NV_NVDLA_CDMA_dc.scala 719:37:@4725.6]
  assign _GEN_185 = {{3'd0}, _T_881}; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4727.8]
  assign _T_886 = _T_879 + _GEN_185; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4727.8]
  assign _T_887 = _T_879 + _GEN_185; // @[NV_NVDLA_CDMA_dc.scala 720:32:@4728.8]
  assign _GEN_186 = {{2'd0}, _T_883}; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4729.8]
  assign _T_888 = _T_887 - _GEN_186; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4729.8]
  assign _T_889 = $unsigned(_T_888); // @[NV_NVDLA_CDMA_dc.scala 720:46:@4730.8]
  assign _T_890 = _T_889[4:0]; // @[NV_NVDLA_CDMA_dc.scala 720:46:@4731.8]
  assign _GEN_96 = _T_885 ? _T_890 : _T_879; // @[NV_NVDLA_CDMA_dc.scala 719:62:@4726.6]
  assign _GEN_97 = _T_138 ? 5'h0 : _GEN_96; // @[NV_NVDLA_CDMA_dc.scala 715:19:@4721.4]
  assign _GEN_187 = {{1'd0}, _T_896}; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4738.4]
  assign _T_899 = _T_893 + _GEN_187; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4738.4]
  assign _T_900 = _T_893 + _GEN_187; // @[NV_NVDLA_CDMA_dc.scala 732:44:@4739.4]
  assign _T_901 = _T_201 - _T_900; // @[NV_NVDLA_CDMA_dc.scala 733:69:@4740.4]
  assign _T_902 = $unsigned(_T_901); // @[NV_NVDLA_CDMA_dc.scala 733:69:@4741.4]
  assign _T_903 = _T_902[13:0]; // @[NV_NVDLA_CDMA_dc.scala 733:69:@4742.4]
  assign _T_904 = _T_138 ? _T_231 : _T_903; // @[NV_NVDLA_CDMA_dc.scala 733:31:@4743.4]
  assign _GEN_188 = {{2'd0}, _T_239}; // @[NV_NVDLA_CDMA_dc.scala 734:48:@4744.4]
  assign _T_905 = _T_904 > _GEN_188; // @[NV_NVDLA_CDMA_dc.scala 734:48:@4744.4]
  assign _T_906 = _T_904[12:0]; // @[NV_NVDLA_CDMA_dc.scala 734:96:@4745.4]
  assign _T_907 = _T_905 ? {{1'd0}, _T_239} : _T_906; // @[NV_NVDLA_CDMA_dc.scala 734:30:@4746.4]
  assign _T_908 = _T_900 == _T_201; // @[NV_NVDLA_CDMA_dc.scala 735:47:@4747.4]
  assign _GEN_189 = {{13'd0}, _GEN_116}; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4859.4]
  assign _T_985 = _T_195 - _GEN_189; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4859.4]
  assign _T_986 = $unsigned(_T_985); // @[NV_NVDLA_CDMA_dc.scala 834:32:@4860.4]
  assign _T_987 = _T_986[15:0]; // @[NV_NVDLA_CDMA_dc.scala 834:32:@4861.4]
  assign _T_988 = _T_973 == _T_987; // @[NV_NVDLA_CDMA_dc.scala 835:32:@4862.4]
  assign _T_1001 = _GEN_115 & _T_988; // @[NV_NVDLA_CDMA_dc.scala 850:34:@4875.4]
  assign _T_967 = _T_896 - 13'h1; // @[NV_NVDLA_CDMA_dc.scala 813:49:@4835.4]
  assign _T_968 = $unsigned(_T_967); // @[NV_NVDLA_CDMA_dc.scala 813:49:@4836.4]
  assign _T_969 = _T_968[12:0]; // @[NV_NVDLA_CDMA_dc.scala 813:49:@4837.4]
  assign _GEN_190 = {{1'd0}, _T_956}; // @[NV_NVDLA_CDMA_dc.scala 813:32:@4838.4]
  assign _T_970 = _GEN_190 == _T_969; // @[NV_NVDLA_CDMA_dc.scala 813:32:@4838.4]
  assign _T_1002 = _T_1001 & _T_970; // @[NV_NVDLA_CDMA_dc.scala 851:35:@4877.4]
  assign _GEN_191 = {{8'd0}, _T_930}; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4795.4]
  assign _T_945 = _T_213 - _GEN_191; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4795.4]
  assign _T_946 = $unsigned(_T_945); // @[NV_NVDLA_CDMA_dc.scala 777:43:@4796.4]
  assign _T_947 = _T_946[10:0]; // @[NV_NVDLA_CDMA_dc.scala 777:43:@4797.4]
  assign _T_948 = _T_927 == _T_947; // @[NV_NVDLA_CDMA_dc.scala 778:33:@4798.4]
  assign _T_1003 = _T_1002 & _T_948; // @[NV_NVDLA_CDMA_dc.scala 852:39:@4879.4]
  assign _T_917 = _T_916 == io_reg2dp_batches; // @[NV_NVDLA_CDMA_dc.scala 752:43:@4765.4]
  assign _T_1004 = _T_1003 & _T_917; // @[NV_NVDLA_CDMA_dc.scala 853:42:@4881.4]
  assign _GEN_98 = _T_1004 ? _T_900 : _T_893; // @[NV_NVDLA_CDMA_dc.scala 742:31:@4756.6]
  assign _T_913 = _T_138 | _T_1004; // @[NV_NVDLA_CDMA_dc.scala 745:23:@4759.6]
  assign _GEN_99 = _T_913 ? _T_907 : _T_896; // @[NV_NVDLA_CDMA_dc.scala 745:42:@4760.6]
  assign _GEN_100 = _T_138 ? 14'h0 : _GEN_98; // @[NV_NVDLA_CDMA_dc.scala 738:19:@4752.4]
  assign _GEN_101 = _T_138 ? _T_896 : _GEN_99; // @[NV_NVDLA_CDMA_dc.scala 738:19:@4752.4]
  assign _T_923 = _T_916 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 763:44:@4776.10]
  assign _T_924 = _T_916 + 5'h1; // @[NV_NVDLA_CDMA_dc.scala 763:44:@4777.10]
  assign _GEN_102 = _T_917 ? 5'h0 : _T_924; // @[NV_NVDLA_CDMA_dc.scala 759:31:@4772.8]
  assign _GEN_103 = _T_1003 ? _GEN_102 : _T_916; // @[NV_NVDLA_CDMA_dc.scala 758:32:@4771.6]
  assign _GEN_104 = _T_138 ? 5'h0 : _GEN_103; // @[NV_NVDLA_CDMA_dc.scala 755:19:@4767.4]
  assign _T_935 = _T_927 + _GEN_191; // @[NV_NVDLA_CDMA_dc.scala 774:37:@4785.4]
  assign _T_936 = _T_927 + _GEN_191; // @[NV_NVDLA_CDMA_dc.scala 774:37:@4786.4]
  assign _T_937 = _T_138 | _T_948; // @[NV_NVDLA_CDMA_dc.scala 775:38:@4787.4]
  assign _T_938 = _T_213 - _T_936; // @[NV_NVDLA_CDMA_dc.scala 775:84:@4788.4]
  assign _T_939 = $unsigned(_T_938); // @[NV_NVDLA_CDMA_dc.scala 775:84:@4789.4]
  assign _T_940 = _T_939[10:0]; // @[NV_NVDLA_CDMA_dc.scala 775:84:@4790.4]
  assign _T_941 = _T_937 ? {{2'd0}, _T_233} : _T_940; // @[NV_NVDLA_CDMA_dc.scala 775:28:@4791.4]
  assign _T_942 = _T_941 > 11'h1; // @[NV_NVDLA_CDMA_dc.scala 776:42:@4792.4]
  assign _T_943 = _T_941[2:0]; // @[NV_NVDLA_CDMA_dc.scala 776:83:@4793.4]
  assign _T_944 = _T_942 ? 3'h1 : _T_943; // @[NV_NVDLA_CDMA_dc.scala 776:27:@4794.4]
  assign _GEN_105 = _T_948 ? 11'h0 : _T_936; // @[NV_NVDLA_CDMA_dc.scala 784:28:@4805.8]
  assign _GEN_106 = _T_1002 ? _GEN_105 : _T_927; // @[NV_NVDLA_CDMA_dc.scala 783:29:@4804.6]
  assign _GEN_107 = _T_138 ? 11'h0 : _GEN_106; // @[NV_NVDLA_CDMA_dc.scala 780:19:@4800.4]
  assign _T_953 = _T_138 | _T_1002; // @[NV_NVDLA_CDMA_dc.scala 792:19:@4814.4]
  assign _GEN_108 = _T_953 ? _T_944 : _T_930; // @[NV_NVDLA_CDMA_dc.scala 792:35:@4815.4]
  assign _T_964 = _T_956 + 12'h1; // @[NV_NVDLA_CDMA_dc.scala 809:36:@4830.10]
  assign _T_965 = _T_956 + 12'h1; // @[NV_NVDLA_CDMA_dc.scala 809:36:@4831.10]
  assign _GEN_109 = _T_970 ? 12'h0 : _T_965; // @[NV_NVDLA_CDMA_dc.scala 805:27:@4826.8]
  assign _GEN_110 = _T_1001 ? _GEN_109 : _T_956; // @[NV_NVDLA_CDMA_dc.scala 804:28:@4825.6]
  assign _GEN_111 = _T_138 ? 12'h0 : _GEN_110; // @[NV_NVDLA_CDMA_dc.scala 801:19:@4821.4]
  assign _GEN_194 = {{1'd0}, _T_198}; // @[NV_NVDLA_CDMA_dc.scala 820:34:@4844.4]
  assign _T_980 = _T_973 == _GEN_194; // @[NV_NVDLA_CDMA_dc.scala 820:34:@4844.4]
  assign _T_983 = _T_973 + _GEN_189; // @[NV_NVDLA_CDMA_dc.scala 830:36:@4854.10]
  assign _T_984 = _T_973 + _GEN_189; // @[NV_NVDLA_CDMA_dc.scala 830:36:@4855.10]
  assign _GEN_112 = _T_988 ? 16'h0 : _T_984; // @[NV_NVDLA_CDMA_dc.scala 826:27:@4850.8]
  assign _GEN_113 = _GEN_115 ? _GEN_112 : _T_973; // @[NV_NVDLA_CDMA_dc.scala 825:28:@4849.6]
  assign _GEN_114 = _T_138 ? 16'h0 : _GEN_113; // @[NV_NVDLA_CDMA_dc.scala 822:19:@4845.4]
  assign _T_992 = _T_930 == 3'h1; // @[NV_NVDLA_CDMA_dc.scala 839:39:@4865.4]
  assign _T_993 = ~ _T_992; // @[NV_NVDLA_CDMA_dc.scala 839:26:@4866.4]
  assign _T_994 = _T_993 | _T_980; // @[NV_NVDLA_CDMA_dc.scala 839:48:@4867.4]
  assign _T_995 = _T_927[1]; // @[NV_NVDLA_CDMA_dc.scala 841:55:@4868.4]
  assign _T_997 = _T_994 | _T_995; // @[NV_NVDLA_CDMA_dc.scala 840:40:@4870.4]
  assign _T_1023 = _T_930 <= 3'h2; // @[NV_NVDLA_CDMA_dc.scala 882:29:@4903.8]
  assign _GEN_117 = _T_1023 ? 1'h0 : _T_1018; // @[NV_NVDLA_CDMA_dc.scala 882:36:@4904.8]
  assign _GEN_118 = _GEN_115 ? _GEN_117 : 1'h0; // @[NV_NVDLA_CDMA_dc.scala 881:24:@4902.6]
  assign _GEN_196 = {{3'd0}, _GEN_116}; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4915.8]
  assign _T_1026 = _T_1014 + _GEN_196; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4915.8]
  assign _T_1027 = _T_1014 + _GEN_196; // @[NV_NVDLA_CDMA_dc.scala 893:54:@4916.8]
  assign _GEN_119 = _T_1019 ? _T_1027 : _T_1014; // @[NV_NVDLA_CDMA_dc.scala 892:37:@4914.6]
  assign _GEN_120 = _T_138 ? 6'h0 : _GEN_119; // @[NV_NVDLA_CDMA_dc.scala 878:19:@4899.4]
  assign _GEN_121 = _T_138 ? _GEN_118 : _T_1017; // @[NV_NVDLA_CDMA_dc.scala 878:19:@4899.4]
  assign _T_1029 = _T_1014[0]; // @[NV_NVDLA_CDMA_dc.scala 897:66:@4920.4]
  assign _T_1030 = _T_1014[5:1]; // @[NV_NVDLA_CDMA_dc.scala 897:89:@4921.4]
  assign _T_1032 = {2'h0,_T_1029,_T_1030}; // @[Cat.scala 30:58:@4923.4]
  assign _T_1034 = _T_131 | _T_138; // @[NV_NVDLA_CDMA_dc.scala 901:22:@4925.4]
  assign _T_1037 = _T_746 & _GEN_115; // @[NV_NVDLA_CDMA_dc.scala 905:37:@4931.6]
  assign _T_1038 = _T_1037 & _T_997; // @[NV_NVDLA_CDMA_dc.scala 905:49:@4932.6]
  assign _GEN_122 = _T_1034 ? 1'h0 : _T_1038; // @[NV_NVDLA_CDMA_dc.scala 901:33:@4926.4]
  assign _GEN_123 = _GEN_115 ? _T_1032 : _T_1044; // @[Reg.scala 20:19:@4939.4]
  assign _T_1064 = _T_973[0]; // @[NV_NVDLA_CDMA_dc.scala 922:86:@4952.4]
  assign _T_1077 = _T_927[0]; // @[NV_NVDLA_CDMA_dc.scala 933:71:@4965.4]
  assign _T_1078 = ~ _T_1077; // @[NV_NVDLA_CDMA_dc.scala 933:60:@4966.4]
  assign _T_1079 = _T_948 & _T_1078; // @[NV_NVDLA_CDMA_dc.scala 933:58:@4967.4]
  assign _T_1065 = _T_1079 & _T_1064; // @[NV_NVDLA_CDMA_dc.scala 922:75:@4953.4]
  assign _T_1068 = _T_1065 | _T_1077; // @[NV_NVDLA_CDMA_dc.scala 922:91:@4956.4]
  assign _GEN_197 = {{2'd0}, _T_195}; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4958.4]
  assign _T_1071 = _T_1047 + _GEN_197; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4958.4]
  assign _T_1072 = _T_1047 + _GEN_197; // @[NV_NVDLA_CDMA_dc.scala 931:64:@4959.4]
  assign _T_1073 = _T_1077 ? _T_1072 : _T_1047; // @[NV_NVDLA_CDMA_dc.scala 931:34:@4960.4]
  assign _T_1080 = _T_138 | _T_917; // @[NV_NVDLA_CDMA_dc.scala 936:40:@4969.4]
  assign _T_1082 = _T_1050 + _T_207; // @[NV_NVDLA_CDMA_dc.scala 936:96:@4970.4]
  assign _T_1083 = _T_1050 + _T_207; // @[NV_NVDLA_CDMA_dc.scala 936:96:@4971.4]
  assign _T_1084 = _T_1080 ? 18'h0 : _T_1083; // @[NV_NVDLA_CDMA_dc.scala 936:30:@4972.4]
  assign _T_1074 = _T_948 ? _T_1084 : _T_1073; // @[NV_NVDLA_CDMA_dc.scala 930:34:@4961.4]
  assign _T_1075 = _T_138 ? 18'h0 : _T_1074; // @[NV_NVDLA_CDMA_dc.scala 929:31:@4962.4]
  assign _T_1086 = _T_1053 + _T_341; // @[NV_NVDLA_CDMA_dc.scala 939:61:@4974.4]
  assign _T_1087 = _T_1053 + _T_341; // @[NV_NVDLA_CDMA_dc.scala 939:61:@4975.4]
  assign _T_1088 = _T_1053 + _T_338; // @[NV_NVDLA_CDMA_dc.scala 940:39:@4976.4]
  assign _T_1089 = _T_1053 + _T_338; // @[NV_NVDLA_CDMA_dc.scala 940:39:@4977.4]
  assign _T_1090 = _T_908 ? _T_1087 : _T_1089; // @[NV_NVDLA_CDMA_dc.scala 939:29:@4978.4]
  assign _T_1091 = _T_970 ? _T_1075 : _T_1090; // @[NV_NVDLA_CDMA_dc.scala 938:29:@4979.4]
  assign _T_1092 = _T_138 ? 18'h0 : _T_1091; // @[NV_NVDLA_CDMA_dc.scala 937:29:@4980.4]
  assign _T_1103 = _T_973[15:1]; // @[NV_NVDLA_CDMA_dc.scala 946:56:@4985.4]
  assign _T_1104 = _T_973[14:0]; // @[NV_NVDLA_CDMA_dc.scala 947:37:@4986.4]
  assign _T_1105 = _T_1079 ? _T_1103 : _T_1104; // @[NV_NVDLA_CDMA_dc.scala 946:31:@4987.4]
  assign _T_1107 = _T_1098 + _T_1053; // @[NV_NVDLA_CDMA_dc.scala 948:53:@4989.4]
  assign _T_1108 = _T_1098 + _T_1053; // @[NV_NVDLA_CDMA_dc.scala 948:53:@4990.4]
  assign _GEN_198 = {{3'd0}, _T_1095}; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4991.4]
  assign _T_1109 = _GEN_198 + _T_1108; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4991.4]
  assign _T_1110 = _GEN_198 + _T_1108; // @[NV_NVDLA_CDMA_dc.scala 948:33:@4992.4]
  assign _GEN_199 = {{3'd0}, _T_1105}; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4993.4]
  assign _T_1111 = _T_1110 + _GEN_199; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4993.4]
  assign _T_1112 = _T_1110 + _GEN_199; // @[NV_NVDLA_CDMA_dc.scala 948:69:@4994.4]
  assign _T_1114 = {_T_219,9'h0}; // @[Cat.scala 30:58:@4995.4]
  assign _GEN_200 = {{3'd0}, _T_1114}; // @[NV_NVDLA_CDMA_dc.scala 949:41:@4996.4]
  assign _T_1115 = _T_1112 >= _GEN_200; // @[NV_NVDLA_CDMA_dc.scala 949:41:@4996.4]
  assign _T_1116 = ~ _T_1115; // @[NV_NVDLA_CDMA_dc.scala 950:26:@4997.4]
  assign _T_1117 = _T_1112[14:0]; // @[NV_NVDLA_CDMA_dc.scala 950:57:@4998.4]
  assign _T_1120 = _T_1112 - _GEN_200; // @[NV_NVDLA_CDMA_dc.scala 951:35:@5000.4]
  assign _T_1121 = $unsigned(_T_1120); // @[NV_NVDLA_CDMA_dc.scala 951:35:@5001.4]
  assign _T_1122 = _T_1121[17:0]; // @[NV_NVDLA_CDMA_dc.scala 951:35:@5002.4]
  assign _T_1123 = _T_1116 ? {{3'd0}, _T_1117} : _T_1122; // @[NV_NVDLA_CDMA_dc.scala 950:25:@5003.4]
  assign _GEN_124 = _T_145 ? io_status2dma_wr_idx : _T_1095; // @[NV_NVDLA_CDMA_dc.scala 954:27:@5005.4]
  assign _GEN_125 = _T_145 ? 18'h0 : _T_1098; // @[NV_NVDLA_CDMA_dc.scala 954:27:@5005.4]
  assign _T_1127 = _T_138 | _T_1003; // @[NV_NVDLA_CDMA_dc.scala 958:19:@5009.4]
  assign _GEN_126 = _T_1127 ? _T_1084 : _T_1050; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  assign _GEN_127 = _T_1127 ? _T_1075 : _T_1047; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  assign _GEN_128 = _T_1127 ? _T_1092 : _T_1053; // @[NV_NVDLA_CDMA_dc.scala 958:38:@5010.4]
  assign _T_1193 = _T_908 ? _T_335 : _T_332; // @[NV_NVDLA_CDMA_dc.scala 1001:21:@5106.4]
  assign _T_1128 = _T_1098 + _T_1193; // @[NV_NVDLA_CDMA_dc.scala 964:46:@5016.6]
  assign _T_1129 = _T_1098 + _T_1193; // @[NV_NVDLA_CDMA_dc.scala 964:46:@5017.6]
  assign _GEN_129 = _T_1004 ? _T_1129 : _GEN_125; // @[NV_NVDLA_CDMA_dc.scala 963:27:@5015.4]
  assign _GEN_130 = _GEN_115 ? _T_1123 : {{1'd0}, _T_1132}; // @[NV_NVDLA_CDMA_dc.scala 969:23:@5022.4]
  assign _GEN_131 = _GEN_115 ? _T_1068 : _T_1135; // @[Reg.scala 20:19:@5026.4]
  assign _T_1150 = {6'h0,2'h0,3'h0,_GEN_115}; // @[Cat.scala 30:58:@5036.4]
  assign _GEN_132 = _T_1101 ? _T_1135 : _T_1153; // @[Reg.scala 20:19:@5038.4]
  assign _GEN_133 = _T_1101 ? _T_1153 : _T_1155; // @[Reg.scala 20:19:@5042.4]
  assign _GEN_134 = _T_1101 ? _T_1155 : _T_1157; // @[Reg.scala 20:19:@5046.4]
  assign _GEN_138 = _T_1101 ? _T_1132 : _T_1168; // @[Reg.scala 20:19:@5064.4]
  assign _GEN_139 = _T_1101 ? _T_1168 : _T_1170; // @[Reg.scala 20:19:@5068.4]
  assign _GEN_140 = _T_1101 ? _T_1170 : _T_1172; // @[Reg.scala 20:19:@5072.4]
  assign _GEN_141 = _T_1101 ? io_dc2sbuf_p0_rd_data : _T_1175; // @[Reg.scala 20:19:@5077.4]
  assign _GEN_142 = _T_1101 ? _T_1175 : _T_1177; // @[Reg.scala 20:19:@5081.4]
  assign _GEN_143 = _T_1101 ? _T_1177 : _T_1179; // @[Reg.scala 20:19:@5085.4]
  assign _GEN_144 = _T_1101 ? _T_1150 : _T_1182; // @[Reg.scala 20:19:@5090.4]
  assign _GEN_145 = _T_1101 ? _T_1182 : _T_1184; // @[Reg.scala 20:19:@5094.4]
  assign _GEN_146 = _T_1101 ? _T_1184 : _T_1186; // @[Reg.scala 20:19:@5098.4]
  assign _T_1190 = _T_329[14:0]; // @[NV_NVDLA_CDMA_dc.scala 1000:52:@5103.4]
  assign _T_1191 = _T_326[14:0]; // @[NV_NVDLA_CDMA_dc.scala 1000:75:@5104.4]
  assign _T_1192 = _T_374 ? _T_1190 : _T_1191; // @[NV_NVDLA_CDMA_dc.scala 1000:24:@5105.4]
  assign _T_1194 = ~ _T_725; // @[NV_NVDLA_CDMA_dc.scala 1002:35:@5108.4]
  assign _T_1196 = _T_1194 ? 15'h0 : _T_1192; // @[NV_NVDLA_CDMA_dc.scala 1002:33:@5109.4]
  assign _T_1197 = ~ io_dc2status_dat_updt_valid; // @[NV_NVDLA_CDMA_dc.scala 1003:35:@5110.4]
  assign _T_1199 = _T_1197 ? 15'h0 : io_dc2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_dc.scala 1003:33:@5111.4]
  assign _T_1200 = _T_725 | io_dc2status_dat_updt_valid; // @[NV_NVDLA_CDMA_dc.scala 1005:27:@5112.4]
  assign _T_1201 = _T_1189 + _T_1196; // @[NV_NVDLA_CDMA_dc.scala 1006:42:@5114.6]
  assign _T_1202 = _T_1189 + _T_1196; // @[NV_NVDLA_CDMA_dc.scala 1006:42:@5115.6]
  assign _T_1203 = _T_1202 - _T_1199; // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5116.6]
  assign _T_1204 = $unsigned(_T_1203); // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5117.6]
  assign _T_1205 = _T_1204[14:0]; // @[NV_NVDLA_CDMA_dc.scala 1006:63:@5118.6]
  assign _GEN_147 = _T_1200 ? _T_1205 : _T_1189; // @[NV_NVDLA_CDMA_dc.scala 1005:57:@5113.4]
  assign _T_1206 = _T_1189 + _T_1192; // @[NV_NVDLA_CDMA_dc.scala 1010:43:@5121.4]
  assign _GEN_202 = {{1'd0}, io_status2dma_free_entries}; // @[NV_NVDLA_CDMA_dc.scala 1011:51:@5122.4]
  assign _T_1207 = _T_1206 <= _GEN_202; // @[NV_NVDLA_CDMA_dc.scala 1011:51:@5122.4]
  assign _T_1208 = _T_908 ? 14'h0 : _T_344; // @[NV_NVDLA_CDMA_dc.scala 1012:24:@5123.4]
  assign _T_1210 = ~ _T_395; // @[NV_NVDLA_CDMA_dc.scala 1014:41:@5125.4]
  assign _T_1211 = _T_131 | _T_1210; // @[NV_NVDLA_CDMA_dc.scala 1014:39:@5126.4]
  assign _T_1212 = _T_1211 | _T_725; // @[NV_NVDLA_CDMA_dc.scala 1014:56:@5127.4]
  assign _T_1214 = _T_1212 ? 1'h0 : _T_1207; // @[NV_NVDLA_CDMA_dc.scala 1014:25:@5128.4]
  assign _GEN_151 = _T_1004 ? _T_1193 : {{3'd0}, _T_1225}; // @[Reg.scala 20:19:@5144.4]
  assign _GEN_152 = _T_1004 ? _T_1225 : _T_1227; // @[Reg.scala 20:19:@5148.4]
  assign _GEN_153 = _T_1004 ? _T_1227 : _T_1229; // @[Reg.scala 20:19:@5152.4]
  assign _GEN_154 = _T_1004 ? _T_1208 : _T_1232; // @[Reg.scala 20:19:@5157.4]
  assign _GEN_155 = _T_1004 ? _T_1232 : _T_1234; // @[Reg.scala 20:19:@5161.4]
  assign _GEN_156 = _T_1004 ? _T_1234 : _T_1236; // @[Reg.scala 20:19:@5165.4]
  assign _T_1237 = ~ _T_673; // @[NV_NVDLA_CDMA_dc.scala 1025:52:@5169.4]
  assign _T_1238 = _T_740 & _T_1237; // @[NV_NVDLA_CDMA_dc.scala 1025:50:@5170.4]
  assign _T_1239 = _T_1238 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_dc.scala 1025:68:@5171.4]
  assign _T_1243 = io_status2dma_fsm_switch & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_dc.scala 1026:60:@5174.4]
  assign _T_1247 = io_reg2dp_op_en & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_dc.scala 1027:51:@5177.4]
  assign _T_1258 = _T_770 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_dc.scala 1041:56:@5194.4]
  assign _T_1270 = NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1045:41:@5202.4 NV_NVDLA_CDMA_dc.scala 1055:31:@5215.4]
  assign _T_1272 = _T_1270 != 9'h1ff; // @[NV_NVDLA_CDMA_dc.scala 1046:48:@5203.4]
  assign _T_1277 = ~ io_dp2reg_dc_rd_latency; // @[NV_NVDLA_CDMA_dc.scala 1058:47:@5216.4]
  assign _T_1279 = _T_1277 == 32'h0; // @[NV_NVDLA_CDMA_dc.scala 1058:47:@5217.4]
  assign _T_1280 = ~ _T_1279; // @[NV_NVDLA_CDMA_dc.scala 1058:22:@5218.4]
  assign _T_1282 = _T_1270 != 9'h0; // @[NV_NVDLA_CDMA_dc.scala 1058:82:@5219.4]
  assign io_dc_dat2mcif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 584:30:@4559.4]
  assign io_dc_dat2mcif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 584:30:@4558.4]
  assign io_mcif2dc_dat_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 593:47:@4570.4]
  assign io_dc_dat2cvif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 586:38:@4562.4]
  assign io_dc_dat2cvif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 586:38:@4561.4]
  assign io_cvif2dc_dat_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 595:55:@4573.4]
  assign io_dc2cvt_dat_wr_sel = _T_1157; // @[NV_NVDLA_CDMA_dc.scala 987:34:@5049.4]
  assign io_dc2cvt_dat_wr_addr_valid = _T_1165; // @[NV_NVDLA_CDMA_dc.scala 989:33:@5062.4]
  assign io_dc2cvt_dat_wr_addr_bits = _T_1172; // @[NV_NVDLA_CDMA_dc.scala 990:32:@5075.4]
  assign io_dc2cvt_dat_wr_data = _T_1179; // @[NV_NVDLA_CDMA_dc.scala 992:31:@5088.4]
  assign io_dc2cvt_dat_wr_info_pd = _T_1186; // @[NV_NVDLA_CDMA_dc.scala 994:30:@5101.4]
  assign io_dp2reg_dc_rd_stall = NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1037:27:@5188.4]
  assign io_dp2reg_dc_rd_latency = NV_COUNTER_STAGE_histogram_2_io_cnt_cur; // @[NV_NVDLA_CDMA_dc.scala 1067:29:@5229.4]
  assign io_dc2status_state = _T_148; // @[NV_NVDLA_CDMA_dc.scala 145:24:@3965.4]
  assign io_dc2status_dat_updt_valid = _T_1222; // @[NV_NVDLA_CDMA_dc.scala 1017:33:@5142.4]
  assign io_dc2status_dat_updt_bits_entries = _T_1229; // @[NV_NVDLA_CDMA_dc.scala 1018:40:@5155.4]
  assign io_dc2status_dat_updt_bits_slices = _T_1236; // @[NV_NVDLA_CDMA_dc.scala 1019:39:@5168.4]
  assign io_dc2sbuf_p0_wr_addr_valid = _T_842 & _T_746; // @[NV_NVDLA_CDMA_dc.scala 700:33:@4712.4]
  assign io_dc2sbuf_p0_wr_addr_bits = _T_864 | _T_870; // @[NV_NVDLA_CDMA_dc.scala 701:32:@4713.4]
  assign io_dc2sbuf_p0_wr_data = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits[255:0]; // @[NV_NVDLA_CDMA_dc.scala 702:27:@4715.4]
  assign io_dc2sbuf_p0_rd_addr_valid = _T_1041; // @[NV_NVDLA_CDMA_dc.scala 909:33:@4937.4]
  assign io_dc2sbuf_p0_rd_addr_bits = _T_1044; // @[NV_NVDLA_CDMA_dc.scala 910:32:@4942.4]
  assign NV_NVDLA_DMAIF_rdreq_reset = reset; // @[:@4552.4]
  assign NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 577:47:@4553.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid = _T_671 & _T_642; // @[NV_NVDLA_CDMA_dc.scala 580:54:@4555.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits = {_T_731,_T_742}; // @[NV_NVDLA_CDMA_dc.scala 582:53:@4557.4]
  assign NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready = io_dc_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 584:30:@4560.4]
  assign NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready = io_dc_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dc.scala 586:38:@4563.4]
  assign NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type = io_reg2dp_datain_ram_type; // @[NV_NVDLA_CDMA_dc.scala 578:52:@4554.4]
  assign NV_NVDLA_DMAIF_rdrsp_reset = reset; // @[:@4566.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 591:47:@4567.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid = io_mcif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 593:47:@4569.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits = io_mcif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 593:47:@4568.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid = io_cvif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dc.scala 595:55:@4572.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits = io_cvif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dc.scala 595:55:@4571.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready = ~ _T_738; // @[NV_NVDLA_CDMA_dc.scala 600:54:@4574.4]
  assign NV_NVDLA_fifo_clock = io_nvdla_core_clk; // @[:@4591.4]
  assign NV_NVDLA_fifo_reset = reset; // @[:@4592.4]
  assign NV_NVDLA_fifo_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 618:19:@4593.4]
  assign NV_NVDLA_fifo_io_wr_pvld = _T_642 & _T_673; // @[NV_NVDLA_CDMA_dc.scala 620:23:@4595.4]
  assign NV_NVDLA_fifo_io_wr_pd = {_T_657,_T_651}; // @[NV_NVDLA_CDMA_dc.scala 622:21:@4597.4]
  assign NV_NVDLA_fifo_io_rd_prdy = _T_768 & _T_764; // @[NV_NVDLA_CDMA_dc.scala 624:23:@4598.4]
  assign NV_COUNTER_STAGE_histogram_reset = reset; // @[:@5182.4]
  assign NV_COUNTER_STAGE_histogram_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 1032:16:@5183.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_inc = _T_1242; // @[NV_NVDLA_CDMA_dc.scala 1033:25:@5184.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_clr = _T_1246; // @[NV_NVDLA_CDMA_dc.scala 1035:25:@5186.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_cen = _T_1250; // @[NV_NVDLA_CDMA_dc.scala 1036:25:@5187.4]
  assign NV_COUNTER_STAGE_histogram_1_reset = reset; // @[:@5209.4]
  assign NV_COUNTER_STAGE_histogram_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 1050:18:@5210.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc = _T_1272 & _T_1257; // @[NV_NVDLA_CDMA_dc.scala 1051:27:@5211.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec = _T_1272 & _T_1261; // @[NV_NVDLA_CDMA_dc.scala 1052:27:@5212.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr = _T_1264; // @[NV_NVDLA_CDMA_dc.scala 1053:27:@5213.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen = _T_1268; // @[NV_NVDLA_CDMA_dc.scala 1054:27:@5214.4]
  assign NV_COUNTER_STAGE_histogram_2_reset = reset; // @[:@5223.4]
  assign NV_COUNTER_STAGE_histogram_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dc.scala 1062:18:@5224.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc = _T_1280 & _T_1282; // @[NV_NVDLA_CDMA_dc.scala 1063:27:@5225.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr = _T_1264; // @[NV_NVDLA_CDMA_dc.scala 1065:27:@5227.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen = _T_1268; // @[NV_NVDLA_CDMA_dc.scala 1066:27:@5228.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_85 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_91 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_116 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_119 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_154 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_151 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_893 = _RAND_6[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_201 = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_108 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_148 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_195 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_198 = _RAND_11[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_204 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_207 = _RAND_13[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_210 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_213 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_216 = _RAND_16[38:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_219 = _RAND_17[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_254 = _RAND_18[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_257 = _RAND_19[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_260 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_263 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_298 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_350 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_320 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_323 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_286 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_289 = _RAND_27[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_292 = _RAND_28[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_295 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_314 = _RAND_30[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_317 = _RAND_31[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_326 = _RAND_32[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_329 = _RAND_33[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_332 = _RAND_34[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_335 = _RAND_35[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_338 = _RAND_36[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_341 = _RAND_37[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_344 = _RAND_38[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_374 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_423 = _RAND_40[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_464 = _RAND_41[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_461 = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_458 = _RAND_43[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_455 = _RAND_44[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_420 = _RAND_45[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_411 = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_452 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  _T_611 = _RAND_48[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_648 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_642 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  _T_602 = _RAND_51[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {2{`RANDOM}};
  _T_605 = _RAND_52[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  _T_608 = _RAND_53[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {2{`RANDOM}};
  _T_645 = _RAND_54[58:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_651 = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_654 = _RAND_56[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_657 = _RAND_57[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_738 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_753 = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_775 = _RAND_60[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_778 = _RAND_61[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_781 = _RAND_62[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_784 = _RAND_63[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_879 = _RAND_64[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1017 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_896 = _RAND_66[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_973 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_956 = _RAND_68[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_927 = _RAND_69[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_930 = _RAND_70[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_916 = _RAND_71[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1014 = _RAND_72[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1041 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1044 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1047 = _RAND_75[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1050 = _RAND_76[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1053 = _RAND_77[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1095 = _RAND_78[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1098 = _RAND_79[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1101 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1132 = _RAND_81[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1135 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1153 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1155 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1157 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1161 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1163 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1165 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1168 = _RAND_89[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1170 = _RAND_90[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1172 = _RAND_91[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {8{`RANDOM}};
  _T_1175 = _RAND_92[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {8{`RANDOM}};
  _T_1177 = _RAND_93[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {8{`RANDOM}};
  _T_1179 = _RAND_94[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1182 = _RAND_95[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1184 = _RAND_96[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1186 = _RAND_97[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1189 = _RAND_98[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1218 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1220 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1222 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1225 = _RAND_102[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1227 = _RAND_103[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1229 = _RAND_104[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1232 = _RAND_105[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1234 = _RAND_106[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1236 = _RAND_107[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1242 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1246 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1250 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1257 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1261 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1264 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1268 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_85 <= 1'h0;
    end else begin
      if (_T_157) begin
        _T_85 <= _T_158;
      end
    end
    if (reset) begin
      _T_116 <= 5'h1f;
    end else begin
      if (_T_157) begin
        _T_116 <= io_reg2dp_data_bank;
      end
    end
    if (reset) begin
      _T_119 <= 1'h0;
    end else begin
      if (_T_157) begin
        _T_119 <= _T_130;
      end
    end
    if (reset) begin
      _T_154 <= 1'h0;
    end else begin
      if (_T_157) begin
        _T_154 <= _T_151;
      end
    end
    if (reset) begin
      _T_151 <= 1'h0;
    end else begin
      if (_T_157) begin
        _T_151 <= io_sc2cdma_dat_pending_req;
      end
    end
  end
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_91 <= 2'h0;
    end else begin
      if (_T_94) begin
        if (_T_95) begin
          _T_91 <= 2'h1;
        end else begin
          if (_T_98) begin
            _T_91 <= 2'h3;
          end else begin
            if (_T_130) begin
              _T_91 <= 2'h2;
            end else begin
              _T_91 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_99) begin
          if (_T_156) begin
            _T_91 <= 2'h2;
          end else begin
            _T_91 <= 2'h0;
          end
        end else begin
          if (_T_100) begin
            if (_T_122) begin
              _T_91 <= 2'h3;
            end else begin
              _T_91 <= 2'h0;
            end
          end else begin
            _T_91 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_893 <= 14'h0;
    end else begin
      if (_T_138) begin
        _T_893 <= 14'h0;
      end else begin
        if (_T_1004) begin
          _T_893 <= _T_900;
        end
      end
    end
    if (reset) begin
      _T_201 <= 14'h0;
    end else begin
      if (_T_138) begin
        _T_201 <= _T_231;
      end
    end
    if (reset) begin
      _T_108 <= 5'h0;
    end else begin
      if (_T_131) begin
        _T_108 <= 5'h0;
      end else begin
        if (_T_911) begin
          _T_108 <= _T_135;
        end
      end
    end
    if (reset) begin
      _T_148 <= 2'h0;
    end else begin
      if (_T_94) begin
        if (_T_95) begin
          _T_148 <= 2'h1;
        end else begin
          if (_T_98) begin
            _T_148 <= 2'h3;
          end else begin
            if (_T_130) begin
              _T_148 <= 2'h2;
            end else begin
              _T_148 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_99) begin
          if (_T_156) begin
            _T_148 <= 2'h2;
          end else begin
            _T_148 <= 2'h0;
          end
        end else begin
          if (_T_100) begin
            if (_T_122) begin
              _T_148 <= 2'h3;
            end else begin
              _T_148 <= 2'h0;
            end
          end else begin
            _T_148 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_195 <= 16'h0;
    end else begin
      if (_T_138) begin
        _T_195 <= {{2'd0}, _GEN_23};
      end
    end
    if (reset) begin
      _T_198 <= 15'h0;
    end else begin
      if (_T_138) begin
        _T_198 <= {{2'd0}, _T_244};
      end
    end
    if (reset) begin
      _T_204 <= 6'h0;
    end else begin
      if (_T_138) begin
        _T_204 <= _T_246;
      end
    end
    if (reset) begin
      _T_207 <= 18'h0;
    end else begin
      if (_T_138) begin
        _T_207 <= {{1'd0}, _T_249};
      end
    end
    if (reset) begin
      _T_210 <= 13'h0;
    end else begin
      if (_T_138) begin
        _T_210 <= {{1'd0}, _T_239};
      end
    end
    if (reset) begin
      _T_213 <= 11'h0;
    end else begin
      if (_T_138) begin
        _T_213 <= {{2'd0}, _T_233};
      end
    end
    if (reset) begin
      _T_216 <= 39'h0;
    end else begin
      if (_T_138) begin
        _T_216 <= _T_240;
      end
    end
    if (reset) begin
      _T_219 <= 6'h0;
    end else begin
      if (_T_138) begin
        _T_219 <= _T_251;
      end
    end
    if (reset) begin
      _T_254 <= 14'h0;
    end else begin
      if (_T_138) begin
        _T_254 <= 14'h0;
      end else begin
        if (_T_270) begin
          _T_254 <= _T_278;
        end
      end
    end
    if (reset) begin
      _T_257 <= 14'h0;
    end else begin
      if (_T_270) begin
        if (_T_274) begin
          _T_257 <= _T_273;
        end else begin
          _T_257 <= {{1'd0}, _T_210};
        end
      end
    end
    if (reset) begin
      _T_260 <= 1'h0;
    end else begin
      if (_T_270) begin
        _T_260 <= _T_274;
      end
    end
    if (reset) begin
      _T_263 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_263 <= 1'h0;
      end else begin
        if (_T_268) begin
          _T_263 <= 1'h1;
        end else begin
          if (_T_306) begin
            _T_263 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_298 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_298 <= 1'h0;
      end else begin
        if (_T_263) begin
          _T_298 <= 1'h1;
        end else begin
          if (_T_365) begin
            _T_298 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_350 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_350 <= 1'h0;
      end else begin
        if (_T_366) begin
          _T_350 <= _T_401;
        end
      end
    end
    if (reset) begin
      _T_320 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_320 <= 1'h0;
      end else begin
        if (_T_356) begin
          _T_320 <= 1'h1;
        end else begin
          if (_T_381) begin
            _T_320 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_323 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_323 <= 1'h0;
      end else begin
        if (_T_359) begin
          _T_323 <= 1'h1;
        end else begin
          if (_T_389) begin
            _T_323 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_286 <= 1'h0;
    end else begin
      _T_286 <= _GEN_40[0];
    end
    if (reset) begin
      _T_289 <= 18'h0;
    end else begin
      if (_T_307) begin
        _T_289 <= _T_304;
      end
    end
    if (reset) begin
      _T_292 <= 14'h0;
    end else begin
      if (!(_T_371)) begin
        if (_T_307) begin
          _T_292 <= _T_257;
        end
      end
    end
    if (reset) begin
      _T_295 <= 1'h0;
    end else begin
      if (_T_307) begin
        _T_295 <= _T_260;
      end
    end
    if (reset) begin
      _T_314 <= 14'h0;
    end else begin
      if (_T_356) begin
        _T_314 <= {{13'd0}, _T_286};
      end
    end
    if (reset) begin
      _T_317 <= 14'h0;
    end else begin
      if (_T_359) begin
        _T_317 <= {{13'd0}, _T_286};
      end
    end
    if (reset) begin
      _T_326 <= 18'h0;
    end else begin
      if (_T_356) begin
        _T_326 <= _T_352;
      end
    end
    if (reset) begin
      _T_329 <= 18'h0;
    end else begin
      if (_T_359) begin
        _T_329 <= _T_352;
      end
    end
    if (reset) begin
      _T_332 <= 18'h0;
    end else begin
      if (_T_369) begin
        _T_332 <= _T_352;
      end
    end
    if (reset) begin
      _T_335 <= 18'h0;
    end else begin
      if (_T_371) begin
        _T_335 <= _T_352;
      end
    end
    if (reset) begin
      _T_338 <= 18'h0;
    end else begin
      if (_T_369) begin
        _T_338 <= _T_289;
      end
    end
    if (reset) begin
      _T_341 <= 18'h0;
    end else begin
      if (_T_371) begin
        _T_341 <= _T_289;
      end
    end
    if (reset) begin
      _T_344 <= 14'h0;
    end else begin
      if (_T_369) begin
        _T_344 <= _T_292;
      end
    end
    if (reset) begin
      _T_374 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_374 <= 1'h0;
      end else begin
        if (_T_725) begin
          _T_374 <= _T_404;
        end
      end
    end
    if (reset) begin
      _T_423 <= 3'h0;
    end else begin
      if (_T_447) begin
        if (_T_448) begin
          _T_423 <= 3'h1;
        end else begin
          _T_423 <= _T_449;
        end
      end
    end
    if (reset) begin
      _T_464 <= 14'h0;
    end else begin
      if (_T_599) begin
        if (_T_570) begin
          _T_464 <= 14'h0;
        end else begin
          _T_464 <= _T_532;
        end
      end
    end
    if (reset) begin
      _T_461 <= 14'h0;
    end else begin
      if (_T_598) begin
        if (_T_570) begin
          _T_461 <= 14'h0;
        end else begin
          _T_461 <= _T_532;
        end
      end
    end
    if (reset) begin
      _T_458 <= 14'h0;
    end else begin
      if (_T_597) begin
        if (_T_570) begin
          _T_458 <= 14'h0;
        end else begin
          _T_458 <= _T_532;
        end
      end
    end
    if (reset) begin
      _T_455 <= 14'h0;
    end else begin
      if (_T_596) begin
        if (_T_570) begin
          _T_455 <= 14'h0;
        end else begin
          _T_455 <= _T_532;
        end
      end
    end
    if (reset) begin
      _T_420 <= 11'h0;
    end else begin
      if (_T_138) begin
        _T_420 <= 11'h0;
      end else begin
        if (_T_723) begin
          if (_T_446) begin
            _T_420 <= 11'h0;
          end else begin
            _T_420 <= _T_442;
          end
        end
      end
    end
    if (reset) begin
      _T_411 <= 5'h0;
    end else begin
      if (_T_138) begin
        _T_411 <= 5'h0;
      end else begin
        if (_T_724) begin
          if (_T_417) begin
            _T_411 <= 5'h0;
          end else begin
            _T_411 <= _T_416;
          end
        end
      end
    end
    if (reset) begin
      _T_452 <= 2'h0;
    end else begin
      if (_T_131) begin
        _T_452 <= 2'h0;
      end else begin
        if (_T_683) begin
          if (_T_591) begin
            _T_452 <= 2'h0;
          end else begin
            _T_452 <= _T_595;
          end
        end
      end
    end
    if (reset) begin
      _T_611 <= 59'h0;
    end else begin
      if (_T_639) begin
        if (_T_145) begin
          _T_611 <= _T_612;
        end else begin
          if (_T_630) begin
            _T_611 <= _T_614;
          end else begin
            if (_T_629) begin
              _T_611 <= _T_616;
            end else begin
              if (_T_517) begin
                _T_611 <= _T_619;
              end else begin
                if (_T_588) begin
                  _T_611 <= _T_608;
                end else begin
                  _T_611 <= _T_621;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_648 <= 1'h0;
    end else begin
      if (_T_1212) begin
        _T_648 <= 1'h0;
      end else begin
        _T_648 <= _T_1207;
      end
    end
    if (reset) begin
      _T_642 <= 1'h0;
    end else begin
      if (_T_131) begin
        _T_642 <= 1'h0;
      end else begin
        if (_T_665) begin
          _T_642 <= 1'h1;
        end else begin
          if (_T_674) begin
            _T_642 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_602 <= 59'h0;
    end else begin
      if (_T_639) begin
        if (_T_145) begin
          _T_602 <= _T_612;
        end else begin
          _T_602 <= _T_614;
        end
      end
    end
    if (reset) begin
      _T_605 <= 59'h0;
    end else begin
      if (_T_639) begin
        if (_T_145) begin
          _T_605 <= _T_612;
        end else begin
          if (_T_417) begin
            _T_605 <= _T_614;
          end else begin
            _T_605 <= _T_616;
          end
        end
      end
    end
    if (reset) begin
      _T_608 <= 59'h0;
    end else begin
      if (_T_639) begin
        if (_T_145) begin
          _T_608 <= _T_612;
        end else begin
          if (_T_625) begin
            _T_608 <= _T_614;
          end else begin
            if (_T_446) begin
              _T_608 <= _T_616;
            end else begin
              _T_608 <= _T_619;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_645 <= 59'h0;
    end else begin
      if (_T_680) begin
        _T_645 <= _T_638;
      end
    end
    if (reset) begin
      _T_651 <= 4'h0;
    end else begin
      if (_T_680) begin
        if (_T_562) begin
          _T_651 <= _T_563;
        end else begin
          if (_T_554) begin
            _T_651 <= _T_559;
          end else begin
            _T_651 <= 4'h8;
          end
        end
      end
    end
    if (reset) begin
      _T_654 <= 3'h0;
    end else begin
      _T_654 <= _GEN_85[2:0];
    end
    if (reset) begin
      _T_657 <= 2'h0;
    end else begin
      if (_T_680) begin
        _T_657 <= _T_452;
      end
    end
    if (reset) begin
      _T_738 <= 1'h0;
    end else begin
      if (_T_1034) begin
        _T_738 <= 1'h0;
      end else begin
        _T_738 <= _T_1038;
      end
    end
    if (reset) begin
      _T_753 <= 4'h0;
    end else begin
      if (_T_768) begin
        if (_T_764) begin
          _T_753 <= 4'h0;
        end else begin
          _T_753 <= _T_763;
        end
      end
    end
    if (reset) begin
      _T_775 <= 6'h0;
    end else begin
      if (_T_138) begin
        _T_775 <= 6'h0;
      end else begin
        if (_T_800) begin
          _T_775 <= _T_815;
        end
      end
    end
    if (reset) begin
      _T_778 <= 6'h0;
    end else begin
      if (!(_T_138)) begin
        if (_T_804) begin
          _T_778 <= _T_817;
        end
      end
    end
    if (reset) begin
      _T_781 <= 6'h0;
    end else begin
      if (!(_T_138)) begin
        if (_T_808) begin
          _T_781 <= _T_819;
        end
      end
    end
    if (reset) begin
      _T_784 <= 6'h0;
    end else begin
      if (!(_T_138)) begin
        if (_T_812) begin
          _T_784 <= _T_821;
        end
      end
    end
    if (reset) begin
      _T_879 <= 5'h0;
    end else begin
      if (_T_138) begin
        _T_879 <= 5'h0;
      end else begin
        if (_T_885) begin
          _T_879 <= _T_890;
        end
      end
    end
    if (reset) begin
      _T_1017 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_GEN_115) begin
          if (_T_1023) begin
            _T_1017 <= 1'h0;
          end else begin
            _T_1017 <= _T_1018;
          end
        end else begin
          _T_1017 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_896 <= 13'h0;
    end else begin
      if (!(_T_138)) begin
        if (_T_913) begin
          if (_T_905) begin
            _T_896 <= {{1'd0}, _T_239};
          end else begin
            _T_896 <= _T_906;
          end
        end
      end
    end
    if (reset) begin
      _T_973 <= 16'h0;
    end else begin
      if (_T_138) begin
        _T_973 <= 16'h0;
      end else begin
        if (_GEN_115) begin
          if (_T_988) begin
            _T_973 <= 16'h0;
          end else begin
            _T_973 <= _T_984;
          end
        end
      end
    end
    if (reset) begin
      _T_956 <= 12'h0;
    end else begin
      if (_T_138) begin
        _T_956 <= 12'h0;
      end else begin
        if (_T_1001) begin
          if (_T_970) begin
            _T_956 <= 12'h0;
          end else begin
            _T_956 <= _T_965;
          end
        end
      end
    end
    if (reset) begin
      _T_927 <= 11'h0;
    end else begin
      if (_T_138) begin
        _T_927 <= 11'h0;
      end else begin
        if (_T_1002) begin
          if (_T_948) begin
            _T_927 <= 11'h0;
          end else begin
            _T_927 <= _T_936;
          end
        end
      end
    end
    if (reset) begin
      _T_930 <= 3'h0;
    end else begin
      if (_T_953) begin
        if (_T_942) begin
          _T_930 <= 3'h1;
        end else begin
          _T_930 <= _T_943;
        end
      end
    end
    if (reset) begin
      _T_916 <= 5'h0;
    end else begin
      if (_T_138) begin
        _T_916 <= 5'h0;
      end else begin
        if (_T_1003) begin
          if (_T_917) begin
            _T_916 <= 5'h0;
          end else begin
            _T_916 <= _T_924;
          end
        end
      end
    end
    if (reset) begin
      _T_1014 <= 6'h0;
    end else begin
      if (_T_138) begin
        _T_1014 <= 6'h0;
      end else begin
        if (_T_1019) begin
          _T_1014 <= _T_1027;
        end
      end
    end
    if (reset) begin
      _T_1041 <= 1'h0;
    end else begin
      if (_T_1008) begin
        _T_1041 <= _T_1006;
      end else begin
        _T_1041 <= 1'h0;
      end
    end
    if (reset) begin
      _T_1044 <= 8'h0;
    end else begin
      if (_GEN_115) begin
        _T_1044 <= _T_1032;
      end
    end
    if (reset) begin
      _T_1047 <= 18'h0;
    end else begin
      if (_T_1127) begin
        if (_T_138) begin
          _T_1047 <= 18'h0;
        end else begin
          if (_T_948) begin
            if (_T_1080) begin
              _T_1047 <= 18'h0;
            end else begin
              _T_1047 <= _T_1083;
            end
          end else begin
            if (_T_1077) begin
              _T_1047 <= _T_1072;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1050 <= 18'h0;
    end else begin
      if (_T_1127) begin
        if (_T_1080) begin
          _T_1050 <= 18'h0;
        end else begin
          _T_1050 <= _T_1083;
        end
      end
    end
    if (reset) begin
      _T_1053 <= 18'h0;
    end else begin
      if (_T_1127) begin
        if (_T_138) begin
          _T_1053 <= 18'h0;
        end else begin
          if (_T_970) begin
            if (_T_138) begin
              _T_1053 <= 18'h0;
            end else begin
              if (_T_948) begin
                if (_T_1080) begin
                  _T_1053 <= 18'h0;
                end else begin
                  _T_1053 <= _T_1083;
                end
              end else begin
                if (_T_1077) begin
                  _T_1053 <= _T_1072;
                end else begin
                  _T_1053 <= _T_1047;
                end
              end
            end
          end else begin
            if (_T_908) begin
              _T_1053 <= _T_1087;
            end else begin
              _T_1053 <= _T_1089;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1095 <= 15'h0;
    end else begin
      if (_T_145) begin
        _T_1095 <= io_status2dma_wr_idx;
      end
    end
    if (reset) begin
      _T_1098 <= 18'h0;
    end else begin
      if (_T_1004) begin
        _T_1098 <= _T_1129;
      end else begin
        if (_T_145) begin
          _T_1098 <= 18'h0;
        end
      end
    end
    if (reset) begin
      _T_1101 <= 1'h0;
    end else begin
      if (_T_1008) begin
        _T_1101 <= _T_1006;
      end else begin
        _T_1101 <= 1'h0;
      end
    end
    if (reset) begin
      _T_1132 <= 17'h0;
    end else begin
      _T_1132 <= _GEN_130[16:0];
    end
    if (reset) begin
      _T_1135 <= 1'h0;
    end else begin
      if (_GEN_115) begin
        _T_1135 <= _T_1068;
      end
    end
    if (reset) begin
      _T_1153 <= 1'h0;
    end else begin
      if (_T_1101) begin
        _T_1153 <= _T_1135;
      end
    end
    if (reset) begin
      _T_1155 <= 1'h0;
    end else begin
      if (_T_1101) begin
        _T_1155 <= _T_1153;
      end
    end
    if (reset) begin
      _T_1157 <= 1'h0;
    end else begin
      if (_T_1101) begin
        _T_1157 <= _T_1155;
      end
    end
    if (reset) begin
      _T_1161 <= 1'h0;
    end else begin
      _T_1161 <= _T_1101;
    end
    if (reset) begin
      _T_1163 <= 1'h0;
    end else begin
      _T_1163 <= _T_1161;
    end
    if (reset) begin
      _T_1165 <= 1'h0;
    end else begin
      _T_1165 <= _T_1163;
    end
    if (reset) begin
      _T_1168 <= 17'h0;
    end else begin
      if (_T_1101) begin
        _T_1168 <= _T_1132;
      end
    end
    if (reset) begin
      _T_1170 <= 17'h0;
    end else begin
      if (_T_1101) begin
        _T_1170 <= _T_1168;
      end
    end
    if (reset) begin
      _T_1172 <= 17'h0;
    end else begin
      if (_T_1101) begin
        _T_1172 <= _T_1170;
      end
    end
    if (reset) begin
      _T_1175 <= 256'h0;
    end else begin
      if (_T_1101) begin
        _T_1175 <= io_dc2sbuf_p0_rd_data;
      end
    end
    if (reset) begin
      _T_1177 <= 256'h0;
    end else begin
      if (_T_1101) begin
        _T_1177 <= _T_1175;
      end
    end
    if (reset) begin
      _T_1179 <= 256'h0;
    end else begin
      if (_T_1101) begin
        _T_1179 <= _T_1177;
      end
    end
    if (reset) begin
      _T_1182 <= 12'h0;
    end else begin
      if (_T_1101) begin
        _T_1182 <= _T_1150;
      end
    end
    if (reset) begin
      _T_1184 <= 12'h0;
    end else begin
      if (_T_1101) begin
        _T_1184 <= _T_1182;
      end
    end
    if (reset) begin
      _T_1186 <= 12'h0;
    end else begin
      if (_T_1101) begin
        _T_1186 <= _T_1184;
      end
    end
    if (reset) begin
      _T_1189 <= 15'h0;
    end else begin
      if (_T_1200) begin
        _T_1189 <= _T_1205;
      end
    end
    if (reset) begin
      _T_1218 <= 1'h0;
    end else begin
      _T_1218 <= _T_1004;
    end
    if (reset) begin
      _T_1220 <= 1'h0;
    end else begin
      _T_1220 <= _T_1218;
    end
    if (reset) begin
      _T_1222 <= 1'h0;
    end else begin
      _T_1222 <= _T_1220;
    end
    if (reset) begin
      _T_1225 <= 15'h0;
    end else begin
      _T_1225 <= _GEN_151[14:0];
    end
    if (reset) begin
      _T_1227 <= 15'h0;
    end else begin
      if (_T_1004) begin
        _T_1227 <= _T_1225;
      end
    end
    if (reset) begin
      _T_1229 <= 15'h0;
    end else begin
      if (_T_1004) begin
        _T_1229 <= _T_1227;
      end
    end
    if (reset) begin
      _T_1232 <= 14'h0;
    end else begin
      if (_T_1004) begin
        if (_T_908) begin
          _T_1232 <= 14'h0;
        end else begin
          _T_1232 <= _T_344;
        end
      end
    end
    if (reset) begin
      _T_1234 <= 14'h0;
    end else begin
      if (_T_1004) begin
        _T_1234 <= _T_1232;
      end
    end
    if (reset) begin
      _T_1236 <= 14'h0;
    end else begin
      if (_T_1004) begin
        _T_1236 <= _T_1234;
      end
    end
    if (reset) begin
      _T_1242 <= 1'h0;
    end else begin
      _T_1242 <= _T_1239;
    end
    if (reset) begin
      _T_1246 <= 1'h0;
    end else begin
      _T_1246 <= _T_1243;
    end
    if (reset) begin
      _T_1250 <= 1'h0;
    end else begin
      _T_1250 <= _T_1247;
    end
    if (reset) begin
      _T_1257 <= 1'h0;
    end else begin
      _T_1257 <= _T_1239;
    end
    if (reset) begin
      _T_1261 <= 1'h0;
    end else begin
      _T_1261 <= _T_1258;
    end
    if (reset) begin
      _T_1264 <= 1'h0;
    end else begin
      _T_1264 <= io_status2dma_fsm_switch;
    end
    if (reset) begin
      _T_1268 <= 1'h0;
    end else begin
      _T_1268 <= _T_1247;
    end
  end
endmodule
module NV_NVDLA_slcg_1( // @[:@5231.2]
  input   io_nvdla_clock_nvdla_core_clk, // @[:@5234.4]
  output  io_nvdla_core_gated_clk // @[:@5234.4]
);
  assign io_nvdla_core_gated_clk = io_nvdla_clock_nvdla_core_clk; // @[slcg.scala 23:31:@5236.4]
endmodule
module NV_NVDLA_CDMA_IMG_ctrl( // @[:@5238.2]
  input         reset, // @[:@5240.4]
  input         io_nvdla_core_clk, // @[:@5241.4]
  input         io_nvdla_core_ng_clk, // @[:@5241.4]
  input         io_pack_is_done, // @[:@5241.4]
  input         io_sc2cdma_dat_pending_req, // @[:@5241.4]
  input         io_sg_is_done, // @[:@5241.4]
  output [1:0]  io_img2status_state, // @[:@5241.4]
  output        io_is_running, // @[:@5241.4]
  output        io_layer_st, // @[:@5241.4]
  output [5:0]  io_pixel_bank, // @[:@5241.4]
  output        io_pixel_early_end, // @[:@5241.4]
  output [10:0] io_pixel_order, // @[:@5241.4]
  output        io_pixel_packed_10b, // @[:@5241.4]
  output        io_pixel_planar, // @[:@5241.4]
  output [1:0]  io_pixel_precision, // @[:@5241.4]
  output        io_pixel_uint, // @[:@5241.4]
  output [3:0]  io_pixel_planar0_bundle_limit, // @[:@5241.4]
  output [3:0]  io_pixel_planar0_bundle_limit_1st, // @[:@5241.4]
  output [4:0]  io_pixel_planar0_byte_sft, // @[:@5241.4]
  output [3:0]  io_pixel_planar0_lp_burst, // @[:@5241.4]
  output        io_pixel_planar0_lp_vld, // @[:@5241.4]
  output [3:0]  io_pixel_planar0_rp_burst, // @[:@5241.4]
  output        io_pixel_planar0_rp_vld, // @[:@5241.4]
  output [2:0]  io_pixel_planar0_sft, // @[:@5241.4]
  output [13:0] io_pixel_planar0_width_burst, // @[:@5241.4]
  output [4:0]  io_pixel_planar1_bundle_limit, // @[:@5241.4]
  output [4:0]  io_pixel_planar1_bundle_limit_1st, // @[:@5241.4]
  output [4:0]  io_pixel_planar1_byte_sft, // @[:@5241.4]
  output [2:0]  io_pixel_planar1_lp_burst, // @[:@5241.4]
  output        io_pixel_planar1_lp_vld, // @[:@5241.4]
  output [2:0]  io_pixel_planar1_rp_burst, // @[:@5241.4]
  output        io_pixel_planar1_rp_vld, // @[:@5241.4]
  output [2:0]  io_pixel_planar1_sft, // @[:@5241.4]
  output [13:0] io_pixel_planar1_width_burst, // @[:@5241.4]
  input         io_reg2dp_op_en, // @[:@5241.4]
  input         io_reg2dp_conv_mode, // @[:@5241.4]
  input         io_reg2dp_datain_format, // @[:@5241.4]
  input  [5:0]  io_reg2dp_pixel_format, // @[:@5241.4]
  input         io_reg2dp_pixel_sign_override, // @[:@5241.4]
  input  [12:0] io_reg2dp_datain_width, // @[:@5241.4]
  input         io_reg2dp_data_reuse, // @[:@5241.4]
  input         io_reg2dp_skip_data_rls, // @[:@5241.4]
  input  [4:0]  io_reg2dp_data_bank, // @[:@5241.4]
  input  [4:0]  io_reg2dp_pixel_x_offset, // @[:@5241.4]
  input  [4:0]  io_reg2dp_pad_left, // @[:@5241.4]
  input  [5:0]  io_reg2dp_pad_right // @[:@5241.4]
);
  reg  _T_117; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 103:69:@5245.4]
  reg [31:0] _RAND_0;
  reg [1:0] _T_129; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 109:28:@5249.4]
  reg [31:0] _RAND_1;
  wire  _T_132; // @[Conditional.scala 37:30:@5252.4]
  wire  _T_215; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 185:38:@5359.4]
  wire  _T_218; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 187:31:@5361.4]
  wire  _T_219; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 187:39:@5362.4]
  reg [4:0] _T_163; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 148:65:@5308.4]
  reg [31:0] _RAND_2;
  wire  _T_212; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 183:37:@5355.4]
  wire  _T_133; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 114:22:@5254.6]
  wire  _T_134; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:27:@5259.8]
  wire  _T_135; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:50:@5260.8]
  reg  _T_156; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 147:59:@5306.4]
  reg [31:0] _RAND_3;
  wire  _T_213; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 184:26:@5357.4]
  wire  _T_136; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:71:@5261.8]
  wire [1:0] _GEN_0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 116:28:@5266.10]
  wire [1:0] _GEN_1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:85:@5262.8]
  wire [1:0] _GEN_2; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 114:38:@5255.6]
  wire  _T_137; // @[Conditional.scala 37:30:@5271.6]
  reg  _T_169; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 150:65:@5310.4]
  reg [31:0] _RAND_4;
  reg  _T_166; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 149:62:@5309.4]
  reg [31:0] _RAND_5;
  wire  _T_170; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 151:41:@5311.4]
  wire  _T_171; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 151:39:@5312.4]
  wire [1:0] _GEN_3; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 119:32:@5273.8]
  wire  _T_138; // @[Conditional.scala 37:30:@5278.8]
  reg  _T_142; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 132:32:@5292.4]
  reg [31:0] _RAND_6;
  wire  _T_149; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 140:44:@5300.4]
  wire  _T_150; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 140:42:@5301.4]
  wire  _T_198; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:35:@5343.4]
  wire  _T_199; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:33:@5344.4]
  wire  _T_200; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:53:@5345.4]
  wire  _T_201; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:69:@5346.4]
  reg [4:0] _T_197; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 176:28:@5342.4]
  reg [31:0] _RAND_7;
  wire  _T_203; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 180:38:@5347.4]
  wire  _T_204; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 180:25:@5348.4]
  wire [1:0] _GEN_4; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 122:25:@5280.10]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@5279.8]
  wire [1:0] _GEN_8; // @[Conditional.scala 39:67:@5272.6]
  wire [1:0] _GEN_9; // @[Conditional.scala 40:58:@5253.4]
  wire  _T_143; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 134:30:@5293.4]
  wire  _T_146; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 137:30:@5297.4]
  reg [1:0] _T_153; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 143:35:@5303.4]
  reg [31:0] _RAND_8;
  wire  _T_172; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:26:@5314.4]
  wire  _T_173; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 156:38:@5318.6]
  wire  _GEN_10; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  wire [4:0] _GEN_11; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  wire  _GEN_12; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  wire  _T_205; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 181:27:@5350.4]
  wire [5:0] _T_208; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:45:@5351.4]
  wire [4:0] _T_209; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:45:@5352.4]
  wire [4:0] _T_210; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:26:@5353.4]
  wire [5:0] _T_211; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 181:26:@5354.4]
  wire  _T_220; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 189:18:@5364.4]
  wire [5:0] _GEN_15; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 189:28:@5365.4]
  wire  _T_246; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:33:@5384.4]
  wire  _T_250; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:38:@5390.6]
  wire  _T_253; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:38:@5395.8]
  wire  _T_256; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:38:@5400.10]
  wire  _T_259; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:38:@5405.12]
  wire  _T_262; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:38:@5410.14]
  wire  _T_265; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:38:@5415.16]
  wire  _T_268; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:38:@5420.18]
  wire  _T_271; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:38:@5425.20]
  wire  _T_274; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:38:@5430.22]
  wire  _T_277; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:38:@5435.24]
  wire  _T_280; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:38:@5440.26]
  wire [2:0] _GEN_17; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  wire [4:0] _GEN_19; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  wire [4:0] _GEN_20; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  wire  _GEN_21; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [10:0] _GEN_22; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [2:0] _GEN_23; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [2:0] _GEN_24; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [4:0] _GEN_26; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  wire [10:0] _GEN_27; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire  _GEN_28; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire [2:0] _GEN_29; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire [2:0] _GEN_30; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire [4:0] _GEN_31; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire [4:0] _GEN_32; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  wire [10:0] _GEN_33; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire  _GEN_34; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire [2:0] _GEN_35; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire [2:0] _GEN_36; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire [4:0] _GEN_37; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire [4:0] _GEN_38; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  wire [10:0] _GEN_39; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire  _GEN_40; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire [2:0] _GEN_41; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire [2:0] _GEN_42; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire [4:0] _GEN_43; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire [4:0] _GEN_44; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  wire [10:0] _GEN_45; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire  _GEN_46; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire [2:0] _GEN_47; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire [2:0] _GEN_48; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire [4:0] _GEN_49; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire [4:0] _GEN_50; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  wire [10:0] _GEN_51; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire  _GEN_52; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire [2:0] _GEN_53; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire [2:0] _GEN_54; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire [4:0] _GEN_55; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire [4:0] _GEN_56; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  wire [10:0] _GEN_57; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire  _GEN_58; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire [2:0] _GEN_59; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire [2:0] _GEN_60; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire [4:0] _GEN_61; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire [4:0] _GEN_62; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  wire [10:0] _GEN_63; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire  _GEN_64; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire [2:0] _GEN_65; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire [2:0] _GEN_66; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire [4:0] _GEN_67; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire [4:0] _GEN_68; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  wire [10:0] _GEN_69; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire  _GEN_70; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire [2:0] _GEN_71; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire [2:0] _GEN_72; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire [4:0] _GEN_73; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire [4:0] _GEN_74; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  wire [10:0] _GEN_75; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire  _GEN_76; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire [2:0] _GEN_77; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire [2:0] _GEN_78; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire [4:0] _GEN_79; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire [4:0] _GEN_80; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  wire [10:0] _GEN_81; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire  _GEN_82; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire [2:0] _GEN_83; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire [2:0] _GEN_84; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire [4:0] _GEN_85; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire [4:0] _GEN_86; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  wire [2:0] _GEN_87; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire [4:0] _GEN_88; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire [10:0] _GEN_89; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire  _GEN_90; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire [2:0] _GEN_91; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire [4:0] _GEN_92; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  wire  _T_299; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 283:57:@5458.4]
  wire [4:0] _T_300; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 284:60:@5459.4]
  wire [4:0] _T_301; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 285:54:@5460.4]
  wire [4:0] _T_302; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 286:54:@5461.4]
  wire  _T_303; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 287:65:@5462.4]
  wire [4:0] _T_304; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:24:@5463.4]
  wire [3:0] _T_306; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:93:@5464.4]
  wire [4:0] _T_307; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:69:@5465.4]
  wire [4:0] _T_308; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 287:39:@5466.4]
  wire [3:0] _T_309; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:99:@5467.4]
  wire  _T_310; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 289:65:@5468.4]
  wire [4:0] _T_311; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:24:@5469.4]
  wire [3:0] _T_313; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:93:@5470.4]
  wire [4:0] _T_314; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:69:@5471.4]
  wire [4:0] _T_315; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 289:39:@5472.4]
  wire [2:0] _T_316; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:99:@5473.4]
  wire [12:0] _GEN_120; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 291:60:@5474.4]
  wire [13:0] _T_317; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 291:60:@5474.4]
  wire [12:0] _GEN_121; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 292:60:@5475.4]
  wire [13:0] _T_318; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 292:60:@5475.4]
  wire [13:0] _T_319; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 293:66:@5476.4]
  wire [14:0] _T_321; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 293:92:@5477.4]
  wire [13:0] _T_322; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 294:66:@5478.4]
  wire [14:0] _T_324; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 294:92:@5479.4]
  wire [12:0] _GEN_122; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:48:@5480.4]
  wire [13:0] _T_325; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:48:@5480.4]
  wire [13:0] _GEN_123; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:74:@5481.4]
  wire [14:0] _T_326; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:74:@5481.4]
  wire [14:0] _T_327; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 296:57:@5482.4]
  wire [15:0] _T_329; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 296:83:@5483.4]
  wire [15:0] _GEN_124; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5486.4]
  wire [16:0] _T_333; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5486.4]
  wire [16:0] _T_334; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5487.4]
  wire [16:0] _GEN_125; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5488.4]
  wire [17:0] _T_335; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5488.4]
  wire [17:0] _T_336; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5489.4]
  wire [3:0] _T_337; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:123:@5490.4]
  wire [2:0] _T_342; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 299:123:@5495.4]
  wire [4:0] _T_349; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:52:@5499.4]
  wire [5:0] _T_350; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:27:@5500.4]
  wire [6:0] _T_351; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:82:@5501.4]
  wire [7:0] _T_353; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:105:@5502.4]
  wire [4:0] _T_354; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:112:@5503.4]
  wire [7:0] _T_355; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:36:@5504.4]
  wire [8:0] _T_361; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:53:@5506.4]
  wire [2:0] _T_362; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:93:@5507.4]
  wire  _T_364; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 313:34:@5508.4]
  wire  _T_366; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 314:33:@5509.4]
  wire  _T_367; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 313:42:@5510.4]
  wire  _T_369; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 315:34:@5511.4]
  wire [5:0] _T_371; // @[Cat.scala 30:58:@5512.4]
  wire  _T_373; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 316:43:@5513.4]
  wire  _T_374; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 315:42:@5514.4]
  wire  _T_375; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 314:41:@5515.4]
  wire  _T_376; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 312:46:@5516.4]
  wire [5:0] _T_378; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:57:@5518.4]
  wire [5:0] _T_379; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:57:@5519.4]
  wire [4:0] _T_380; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:97:@5520.4]
  wire [9:0] _T_386; // @[Cat.scala 30:58:@5522.4]
  wire [9:0] _T_387; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 321:90:@5523.4]
  wire [4:0] _T_388; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 321:115:@5524.4]
  wire [9:0] _T_395; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 322:90:@5527.4]
  wire [4:0] _T_396; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 322:115:@5528.4]
  wire  _T_403; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 330:59:@5530.4]
  wire  _T_405; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 331:59:@5531.4]
  wire  _T_407; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 332:59:@5532.4]
  wire  _T_409; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 333:59:@5533.4]
  reg  _T_412; // @[Reg.scala 19:20:@5534.4]
  reg [31:0] _RAND_9;
  wire  _GEN_93; // @[Reg.scala 20:19:@5535.4]
  reg [1:0] _T_415; // @[Reg.scala 19:20:@5539.4]
  reg [31:0] _RAND_10;
  wire [1:0] _GEN_94; // @[Reg.scala 20:19:@5540.4]
  reg [10:0] _T_418; // @[Reg.scala 19:20:@5544.4]
  reg [31:0] _RAND_11;
  wire [10:0] _GEN_95; // @[Reg.scala 20:19:@5545.4]
  reg  _T_421; // @[Reg.scala 19:20:@5549.4]
  reg [31:0] _RAND_12;
  wire  _GEN_96; // @[Reg.scala 20:19:@5550.4]
  reg  _T_430; // @[Reg.scala 19:20:@5564.4]
  reg [31:0] _RAND_13;
  wire  _GEN_99; // @[Reg.scala 20:19:@5565.4]
  reg [2:0] _T_433; // @[Reg.scala 19:20:@5569.4]
  reg [31:0] _RAND_14;
  wire [2:0] _GEN_100; // @[Reg.scala 20:19:@5570.4]
  wire  _T_435; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 343:92:@5574.4]
  reg [2:0] _T_437; // @[Reg.scala 19:20:@5575.4]
  reg [31:0] _RAND_15;
  wire [2:0] _GEN_101; // @[Reg.scala 20:19:@5576.4]
  reg [3:0] _T_440; // @[Reg.scala 19:20:@5580.4]
  reg [31:0] _RAND_16;
  wire [3:0] _GEN_102; // @[Reg.scala 20:19:@5581.4]
  reg [2:0] _T_444; // @[Reg.scala 19:20:@5586.4]
  reg [31:0] _RAND_17;
  wire [2:0] _GEN_103; // @[Reg.scala 20:19:@5587.4]
  reg  _T_447; // @[Reg.scala 19:20:@5591.4]
  reg [31:0] _RAND_18;
  wire  _GEN_104; // @[Reg.scala 20:19:@5592.4]
  reg  _T_451; // @[Reg.scala 19:20:@5597.4]
  reg [31:0] _RAND_19;
  wire  _GEN_105; // @[Reg.scala 20:19:@5598.4]
  reg [13:0] _T_454; // @[Reg.scala 19:20:@5602.4]
  reg [31:0] _RAND_20;
  wire [14:0] _GEN_106; // @[Reg.scala 20:19:@5603.4]
  reg [13:0] _T_458; // @[Reg.scala 19:20:@5608.4]
  reg [31:0] _RAND_21;
  wire [14:0] _GEN_107; // @[Reg.scala 20:19:@5609.4]
  reg [3:0] _T_461; // @[Reg.scala 19:20:@5613.4]
  reg [31:0] _RAND_22;
  wire [3:0] _GEN_108; // @[Reg.scala 20:19:@5614.4]
  reg [2:0] _T_465; // @[Reg.scala 19:20:@5619.4]
  reg [31:0] _RAND_23;
  wire [2:0] _GEN_109; // @[Reg.scala 20:19:@5620.4]
  reg  _T_468; // @[Reg.scala 19:20:@5624.4]
  reg [31:0] _RAND_24;
  wire  _GEN_110; // @[Reg.scala 20:19:@5625.4]
  reg  _T_472; // @[Reg.scala 19:20:@5630.4]
  reg [31:0] _RAND_25;
  wire  _GEN_111; // @[Reg.scala 20:19:@5631.4]
  reg  _T_476; // @[Reg.scala 19:20:@5636.4]
  reg [31:0] _RAND_26;
  wire  _GEN_112; // @[Reg.scala 20:19:@5637.4]
  reg [4:0] _T_479; // @[Reg.scala 19:20:@5641.4]
  reg [31:0] _RAND_27;
  wire [4:0] _GEN_113; // @[Reg.scala 20:19:@5642.4]
  reg [4:0] _T_483; // @[Reg.scala 19:20:@5647.4]
  reg [31:0] _RAND_28;
  wire [4:0] _GEN_114; // @[Reg.scala 20:19:@5648.4]
  wire [5:0] _T_485; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 357:52:@5652.4]
  reg [5:0] _T_488; // @[Reg.scala 19:20:@5653.4]
  reg [31:0] _RAND_29;
  wire [5:0] _GEN_115; // @[Reg.scala 20:19:@5654.4]
  reg [3:0] _T_491; // @[Reg.scala 19:20:@5658.4]
  reg [31:0] _RAND_30;
  wire [3:0] _GEN_116; // @[Reg.scala 20:19:@5659.4]
  reg [4:0] _T_495; // @[Reg.scala 19:20:@5664.4]
  reg [31:0] _RAND_31;
  wire [4:0] _GEN_117; // @[Reg.scala 20:19:@5665.4]
  reg [3:0] _T_498; // @[Reg.scala 19:20:@5669.4]
  reg [31:0] _RAND_32;
  wire [3:0] _GEN_118; // @[Reg.scala 20:19:@5670.4]
  reg [4:0] _T_502; // @[Reg.scala 19:20:@5675.4]
  reg [31:0] _RAND_33;
  wire [4:0] _GEN_119; // @[Reg.scala 20:19:@5676.4]
  assign _T_132 = 2'h0 == _T_129; // @[Conditional.scala 37:30:@5252.4]
  assign _T_215 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 185:38:@5359.4]
  assign _T_218 = io_reg2dp_op_en & _T_215; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 187:31:@5361.4]
  assign _T_219 = _T_218 & io_reg2dp_datain_format; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 187:39:@5362.4]
  assign _T_212 = _T_163 != io_reg2dp_data_bank; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 183:37:@5355.4]
  assign _T_133 = _T_219 & _T_212; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 114:22:@5254.6]
  assign _T_134 = _T_219 & io_reg2dp_data_reuse; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:27:@5259.8]
  assign _T_135 = _T_134 & _T_117; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:50:@5260.8]
  assign _T_213 = _T_219 & _T_156; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 184:26:@5357.4]
  assign _T_136 = _T_135 & _T_213; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:71:@5261.8]
  assign _GEN_0 = _T_219 ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 116:28:@5266.10]
  assign _GEN_1 = _T_136 ? 2'h3 : _GEN_0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 115:85:@5262.8]
  assign _GEN_2 = _T_133 ? 2'h1 : _GEN_1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 114:38:@5255.6]
  assign _T_137 = 2'h1 == _T_129; // @[Conditional.scala 37:30:@5271.6]
  assign _T_170 = ~ _T_166; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 151:41:@5311.4]
  assign _T_171 = _T_169 & _T_170; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 151:39:@5312.4]
  assign _GEN_3 = _T_171 ? 2'h2 : 2'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 119:32:@5273.8]
  assign _T_138 = 2'h2 == _T_129; // @[Conditional.scala 37:30:@5278.8]
  assign _T_149 = _T_142 == 1'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 140:44:@5300.4]
  assign _T_150 = io_is_running & _T_149; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 140:42:@5301.4]
  assign _T_198 = ~ _T_150; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:35:@5343.4]
  assign _T_199 = io_is_running & _T_198; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:33:@5344.4]
  assign _T_200 = _T_199 & io_sg_is_done; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:53:@5345.4]
  assign _T_201 = _T_200 & io_pack_is_done; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 178:69:@5346.4]
  assign _T_203 = _T_197 == 5'h9; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 180:38:@5347.4]
  assign _T_204 = _T_201 & _T_203; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 180:25:@5348.4]
  assign _GEN_4 = _T_204 ? 2'h3 : 2'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 122:25:@5280.10]
  assign _GEN_7 = _T_138 ? _GEN_4 : 2'h0; // @[Conditional.scala 39:67:@5279.8]
  assign _GEN_8 = _T_137 ? _GEN_3 : _GEN_7; // @[Conditional.scala 39:67:@5272.6]
  assign _GEN_9 = _T_132 ? _GEN_2 : _GEN_8; // @[Conditional.scala 40:58:@5253.4]
  assign _T_143 = _T_129 == 2'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 134:30:@5293.4]
  assign _T_146 = _T_129 == 2'h3; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 137:30:@5297.4]
  assign _T_172 = io_reg2dp_op_en & _T_143; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:26:@5314.4]
  assign _T_173 = _T_219 & io_reg2dp_skip_data_rls; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 156:38:@5318.6]
  assign _GEN_10 = _T_172 ? _T_219 : _T_156; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  assign _GEN_11 = _T_172 ? io_reg2dp_data_bank : _T_163; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  assign _GEN_12 = _T_172 ? _T_173 : _T_117; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 153:36:@5315.4]
  assign _T_205 = ~ io_is_running; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 181:27:@5350.4]
  assign _T_208 = _T_197 + 5'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:45:@5351.4]
  assign _T_209 = _T_197 + 5'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:45:@5352.4]
  assign _T_210 = _T_201 ? _T_209 : _T_197; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 182:26:@5353.4]
  assign _T_211 = _T_205 ? 6'h0 : {{1'd0}, _T_210}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 181:26:@5354.4]
  assign _T_220 = _T_201 | _T_146; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 189:18:@5364.4]
  assign _GEN_15 = _T_220 ? _T_211 : {{1'd0}, _T_197}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 189:28:@5365.4]
  assign _T_246 = io_reg2dp_pixel_format == 6'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:33:@5384.4]
  assign _T_250 = io_reg2dp_pixel_format == 6'hc; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:38:@5390.6]
  assign _T_253 = io_reg2dp_pixel_format == 6'hd; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:38:@5395.8]
  assign _T_256 = io_reg2dp_pixel_format == 6'he; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:38:@5400.10]
  assign _T_259 = io_reg2dp_pixel_format == 6'hf; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:38:@5405.12]
  assign _T_262 = io_reg2dp_pixel_format == 6'h10; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:38:@5410.14]
  assign _T_265 = io_reg2dp_pixel_format == 6'h11; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:38:@5415.16]
  assign _T_268 = io_reg2dp_pixel_format == 6'h12; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:38:@5420.18]
  assign _T_271 = io_reg2dp_pixel_format == 6'h13; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:38:@5425.20]
  assign _T_274 = io_reg2dp_pixel_format == 6'h1a; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:38:@5430.22]
  assign _T_277 = io_reg2dp_pixel_format == 6'h1b; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:38:@5435.24]
  assign _T_280 = io_reg2dp_pixel_format == 6'h1c; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:38:@5440.26]
  assign _GEN_17 = _T_280 ? 3'h5 : 3'h3; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  assign _GEN_18 = _T_280 ? 3'h4 : 3'h3; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  assign _GEN_19 = _T_280 ? 5'h1f : 5'h7; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  assign _GEN_20 = _T_280 ? 5'hf : 5'h7; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 270:60:@5451.28]
  assign _GEN_21 = _T_280 ? 1'h1 : _T_280; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_22 = _T_280 ? 11'h200 : 11'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_23 = _T_280 ? 3'h5 : _GEN_17; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_24 = _T_280 ? 3'h4 : _GEN_18; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_25 = _T_280 ? 5'h1f : _GEN_19; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_26 = _T_280 ? 5'hf : _GEN_20; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 261:60:@5441.26]
  assign _GEN_27 = _T_277 ? 11'h8 : _GEN_22; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_28 = _T_277 ? 1'h0 : _GEN_21; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_29 = _T_277 ? 3'h3 : _GEN_23; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_30 = _T_277 ? 3'h3 : _GEN_24; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_31 = _T_277 ? 5'h7 : _GEN_25; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_32 = _T_277 ? 5'h7 : _GEN_26; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 257:60:@5436.24]
  assign _GEN_33 = _T_274 ? 11'h2 : _GEN_27; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_34 = _T_274 ? 1'h0 : _GEN_28; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_35 = _T_274 ? 3'h3 : _GEN_29; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_36 = _T_274 ? 3'h3 : _GEN_30; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_37 = _T_274 ? 5'h7 : _GEN_31; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_38 = _T_274 ? 5'h7 : _GEN_32; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 253:60:@5431.22]
  assign _GEN_39 = _T_271 ? 11'h20 : _GEN_33; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_40 = _T_271 ? 1'h0 : _GEN_34; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_41 = _T_271 ? 3'h3 : _GEN_35; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_42 = _T_271 ? 3'h3 : _GEN_36; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_43 = _T_271 ? 5'h7 : _GEN_37; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_44 = _T_271 ? 5'h7 : _GEN_38; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 249:60:@5426.20]
  assign _GEN_45 = _T_268 ? 11'h8 : _GEN_39; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_46 = _T_268 ? 1'h0 : _GEN_40; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_47 = _T_268 ? 3'h3 : _GEN_41; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_48 = _T_268 ? 3'h3 : _GEN_42; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_49 = _T_268 ? 5'h7 : _GEN_43; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_50 = _T_268 ? 5'h7 : _GEN_44; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 245:60:@5421.18]
  assign _GEN_51 = _T_265 ? 11'h2 : _GEN_45; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_52 = _T_265 ? 1'h0 : _GEN_46; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_53 = _T_265 ? 3'h3 : _GEN_47; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_54 = _T_265 ? 3'h3 : _GEN_48; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_55 = _T_265 ? 5'h7 : _GEN_49; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_56 = _T_265 ? 5'h7 : _GEN_50; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 241:60:@5416.16]
  assign _GEN_57 = _T_262 ? 11'h1 : _GEN_51; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_58 = _T_262 ? 1'h0 : _GEN_52; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_59 = _T_262 ? 3'h3 : _GEN_53; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_60 = _T_262 ? 3'h3 : _GEN_54; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_61 = _T_262 ? 5'h7 : _GEN_55; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_62 = _T_262 ? 5'h7 : _GEN_56; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 237:60:@5411.14]
  assign _GEN_63 = _T_259 ? 11'h20 : _GEN_57; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_64 = _T_259 ? 1'h0 : _GEN_58; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_65 = _T_259 ? 3'h3 : _GEN_59; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_66 = _T_259 ? 3'h3 : _GEN_60; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_67 = _T_259 ? 5'h7 : _GEN_61; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_68 = _T_259 ? 5'h7 : _GEN_62; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 233:59:@5406.12]
  assign _GEN_69 = _T_256 ? 11'h8 : _GEN_63; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_70 = _T_256 ? 1'h0 : _GEN_64; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_71 = _T_256 ? 3'h3 : _GEN_65; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_72 = _T_256 ? 3'h3 : _GEN_66; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_73 = _T_256 ? 5'h7 : _GEN_67; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_74 = _T_256 ? 5'h7 : _GEN_68; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 229:59:@5401.10]
  assign _GEN_75 = _T_253 ? 11'h2 : _GEN_69; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_76 = _T_253 ? 1'h0 : _GEN_70; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_77 = _T_253 ? 3'h3 : _GEN_71; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_78 = _T_253 ? 3'h3 : _GEN_72; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_79 = _T_253 ? 5'h7 : _GEN_73; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_80 = _T_253 ? 5'h7 : _GEN_74; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 225:59:@5396.8]
  assign _GEN_81 = _T_250 ? 11'h1 : _GEN_75; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_82 = _T_250 ? 1'h0 : _GEN_76; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_83 = _T_250 ? 3'h3 : _GEN_77; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_84 = _T_250 ? 3'h3 : _GEN_78; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_85 = _T_250 ? 5'h7 : _GEN_79; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_86 = _T_250 ? 5'h7 : _GEN_80; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 221:59:@5391.6]
  assign _GEN_87 = _T_246 ? 3'h5 : _GEN_83; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _GEN_88 = _T_246 ? 5'h1f : _GEN_85; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _GEN_89 = _T_246 ? 11'h1 : _GEN_81; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _GEN_90 = _T_246 ? 1'h0 : _GEN_82; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _GEN_91 = _T_246 ? 3'h3 : _GEN_84; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _GEN_92 = _T_246 ? 5'h7 : _GEN_86; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 216:54:@5385.4]
  assign _T_299 = io_reg2dp_pixel_sign_override == 1'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 283:57:@5458.4]
  assign _T_300 = io_reg2dp_pixel_x_offset & _GEN_92; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 284:60:@5459.4]
  assign _T_301 = io_reg2dp_pad_left & _GEN_88; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 285:54:@5460.4]
  assign _T_302 = io_reg2dp_pad_left & _GEN_92; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 286:54:@5461.4]
  assign _T_303 = io_reg2dp_pixel_x_offset >= _T_301; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 287:65:@5462.4]
  assign _T_304 = io_reg2dp_pad_left >> _GEN_87; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:24:@5463.4]
  assign _T_306 = _GEN_87 + 3'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:93:@5464.4]
  assign _T_307 = io_reg2dp_pad_left >> _T_306; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:69:@5465.4]
  assign _T_308 = _T_303 ? _T_304 : _T_307; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 287:39:@5466.4]
  assign _T_309 = _T_308[3:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 288:99:@5467.4]
  assign _T_310 = io_reg2dp_pixel_x_offset >= _T_302; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 289:65:@5468.4]
  assign _T_311 = io_reg2dp_pad_left >> _GEN_91; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:24:@5469.4]
  assign _T_313 = _GEN_91 + 3'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:93:@5470.4]
  assign _T_314 = io_reg2dp_pad_left >> _T_313; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:69:@5471.4]
  assign _T_315 = _T_310 ? _T_311 : _T_314; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 289:39:@5472.4]
  assign _T_316 = _T_315[2:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 290:99:@5473.4]
  assign _GEN_120 = {{8'd0}, io_reg2dp_pixel_x_offset}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 291:60:@5474.4]
  assign _T_317 = io_reg2dp_datain_width + _GEN_120; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 291:60:@5474.4]
  assign _GEN_121 = {{8'd0}, _T_300}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 292:60:@5475.4]
  assign _T_318 = io_reg2dp_datain_width + _GEN_121; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 292:60:@5475.4]
  assign _T_319 = _T_317 >> _GEN_87; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 293:66:@5476.4]
  assign _T_321 = _T_319 + 14'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 293:92:@5477.4]
  assign _T_322 = _T_318 >> _GEN_91; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 294:66:@5478.4]
  assign _T_324 = _T_322 + 14'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 294:92:@5479.4]
  assign _GEN_122 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:48:@5480.4]
  assign _T_325 = _GEN_122 + io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:48:@5480.4]
  assign _GEN_123 = {{8'd0}, io_reg2dp_pad_right}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:74:@5481.4]
  assign _T_326 = _T_325 + _GEN_123; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 295:74:@5481.4]
  assign _T_327 = _T_326 >> _GEN_87; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 296:57:@5482.4]
  assign _T_329 = _T_327 + 15'h2; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 296:83:@5483.4]
  assign _GEN_124 = {{12'd0}, _T_309}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5486.4]
  assign _T_333 = _T_329 - _GEN_124; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5486.4]
  assign _T_334 = $unsigned(_T_333); // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:64:@5487.4]
  assign _GEN_125 = {{2'd0}, _T_321}; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5488.4]
  assign _T_335 = _T_334 - _GEN_125; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5488.4]
  assign _T_336 = $unsigned(_T_335); // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:92:@5489.4]
  assign _T_337 = _T_336[3:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 298:123:@5490.4]
  assign _T_342 = _T_336[2:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 299:123:@5495.4]
  assign _T_349 = io_reg2dp_datain_width[4:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:52:@5499.4]
  assign _T_350 = io_reg2dp_pad_left + _T_349; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:27:@5500.4]
  assign _T_351 = _T_350 + io_reg2dp_pad_right; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:82:@5501.4]
  assign _T_353 = _T_351 + 7'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:105:@5502.4]
  assign _T_354 = _T_353[4:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 306:112:@5503.4]
  assign _T_355 = _T_354 * 5'h3; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:36:@5504.4]
  assign _T_361 = _T_355 + 8'h1f; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:53:@5506.4]
  assign _T_362 = _T_361[7:5]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 309:93:@5507.4]
  assign _T_364 = _T_362 == 3'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 313:34:@5508.4]
  assign _T_366 = _T_362 == 3'h4; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 314:33:@5509.4]
  assign _T_367 = _T_364 | _T_366; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 313:42:@5510.4]
  assign _T_369 = _T_362 == 3'h2; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 315:34:@5511.4]
  assign _T_371 = {_T_354,1'h0}; // @[Cat.scala 30:58:@5512.4]
  assign _T_373 = _T_371 > 6'h20; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 316:43:@5513.4]
  assign _T_374 = _T_369 & _T_373; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 315:42:@5514.4]
  assign _T_375 = _T_367 | _T_374; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 314:41:@5515.4]
  assign _T_376 = _GEN_90 & _T_375; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 312:46:@5516.4]
  assign _T_378 = io_reg2dp_pixel_x_offset - io_reg2dp_pad_left; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:57:@5518.4]
  assign _T_379 = $unsigned(_T_378); // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:57:@5519.4]
  assign _T_380 = _T_379[4:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 320:97:@5520.4]
  assign _T_386 = {_T_380,5'h0}; // @[Cat.scala 30:58:@5522.4]
  assign _T_387 = _T_386 >> _GEN_87; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 321:90:@5523.4]
  assign _T_388 = _T_387[4:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 321:115:@5524.4]
  assign _T_395 = _T_386 >> _GEN_91; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 322:90:@5527.4]
  assign _T_396 = _T_395[4:0]; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 322:115:@5528.4]
  assign _T_403 = _T_309 != 4'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 330:59:@5530.4]
  assign _T_405 = _T_316 != 3'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 331:59:@5531.4]
  assign _T_407 = _T_337 != 4'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 332:59:@5532.4]
  assign _T_409 = _T_342 != 3'h0; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 333:59:@5533.4]
  assign _GEN_93 = io_layer_st ? _GEN_90 : _T_412; // @[Reg.scala 20:19:@5535.4]
  assign _GEN_94 = io_layer_st ? 2'h0 : _T_415; // @[Reg.scala 20:19:@5540.4]
  assign _GEN_95 = io_layer_st ? _GEN_89 : _T_418; // @[Reg.scala 20:19:@5545.4]
  assign _GEN_96 = io_layer_st ? 1'h0 : _T_421; // @[Reg.scala 20:19:@5550.4]
  assign _GEN_99 = io_layer_st ? _T_299 : _T_430; // @[Reg.scala 20:19:@5565.4]
  assign _GEN_100 = io_layer_st ? _GEN_87 : _T_433; // @[Reg.scala 20:19:@5570.4]
  assign _T_435 = io_layer_st & _GEN_90; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 343:92:@5574.4]
  assign _GEN_101 = _T_435 ? _GEN_91 : _T_437; // @[Reg.scala 20:19:@5576.4]
  assign _GEN_102 = io_layer_st ? _T_309 : _T_440; // @[Reg.scala 20:19:@5581.4]
  assign _GEN_103 = _T_435 ? _T_316 : _T_444; // @[Reg.scala 20:19:@5587.4]
  assign _GEN_104 = io_layer_st ? _T_403 : _T_447; // @[Reg.scala 20:19:@5592.4]
  assign _GEN_105 = _T_435 ? _T_405 : _T_451; // @[Reg.scala 20:19:@5598.4]
  assign _GEN_106 = io_layer_st ? _T_321 : {{1'd0}, _T_454}; // @[Reg.scala 20:19:@5603.4]
  assign _GEN_107 = _T_435 ? _T_324 : {{1'd0}, _T_458}; // @[Reg.scala 20:19:@5609.4]
  assign _GEN_108 = io_layer_st ? _T_337 : _T_461; // @[Reg.scala 20:19:@5614.4]
  assign _GEN_109 = _T_435 ? _T_342 : _T_465; // @[Reg.scala 20:19:@5620.4]
  assign _GEN_110 = io_layer_st ? _T_407 : _T_468; // @[Reg.scala 20:19:@5625.4]
  assign _GEN_111 = _T_435 ? _T_409 : _T_472; // @[Reg.scala 20:19:@5631.4]
  assign _GEN_112 = _T_435 ? _T_376 : _T_476; // @[Reg.scala 20:19:@5637.4]
  assign _GEN_113 = io_layer_st ? _T_388 : _T_479; // @[Reg.scala 20:19:@5642.4]
  assign _GEN_114 = _T_435 ? _T_396 : _T_483; // @[Reg.scala 20:19:@5648.4]
  assign _T_485 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 357:52:@5652.4]
  assign _GEN_115 = io_layer_st ? _T_485 : _T_488; // @[Reg.scala 20:19:@5654.4]
  assign _GEN_116 = io_layer_st ? 4'h8 : _T_491; // @[Reg.scala 20:19:@5659.4]
  assign _GEN_117 = _T_435 ? 5'h10 : _T_495; // @[Reg.scala 20:19:@5665.4]
  assign _GEN_118 = io_layer_st ? 4'h9 : _T_498; // @[Reg.scala 20:19:@5670.4]
  assign _GEN_119 = _T_435 ? 5'h11 : _T_502; // @[Reg.scala 20:19:@5676.4]
  assign io_img2status_state = _T_153; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 143:25:@5305.4]
  assign io_is_running = _T_129 == 2'h2; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 136:19:@5296.4]
  assign io_layer_st = _T_219 & _T_143; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 139:17:@5299.4]
  assign io_pixel_bank = _T_488; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 357:19:@5657.4]
  assign io_pixel_early_end = _T_476; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 354:24:@5640.4]
  assign io_pixel_order = _T_418; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 337:20:@5548.4]
  assign io_pixel_packed_10b = _T_421; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 338:25:@5553.4]
  assign io_pixel_planar = _T_412; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 335:21:@5538.4]
  assign io_pixel_precision = _T_415; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 336:24:@5543.4]
  assign io_pixel_uint = _T_430; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 341:19:@5568.4]
  assign io_pixel_planar0_bundle_limit = _T_491; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 358:35:@5662.4]
  assign io_pixel_planar0_bundle_limit_1st = _T_498; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 360:39:@5673.4]
  assign io_pixel_planar0_byte_sft = _T_479; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 355:31:@5645.4]
  assign io_pixel_planar0_lp_burst = _T_440; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 344:31:@5584.4]
  assign io_pixel_planar0_lp_vld = _T_447; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 346:29:@5595.4]
  assign io_pixel_planar0_rp_burst = _T_461; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 350:31:@5617.4]
  assign io_pixel_planar0_rp_vld = _T_468; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 352:29:@5628.4]
  assign io_pixel_planar0_sft = _T_433; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 342:26:@5573.4]
  assign io_pixel_planar0_width_burst = _T_454; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 348:34:@5606.4]
  assign io_pixel_planar1_bundle_limit = _T_495; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 359:35:@5668.4]
  assign io_pixel_planar1_bundle_limit_1st = _T_502; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 361:39:@5679.4]
  assign io_pixel_planar1_byte_sft = _T_483; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 356:31:@5651.4]
  assign io_pixel_planar1_lp_burst = _T_444; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 345:31:@5590.4]
  assign io_pixel_planar1_lp_vld = _T_451; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 347:29:@5601.4]
  assign io_pixel_planar1_rp_burst = _T_465; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 351:31:@5623.4]
  assign io_pixel_planar1_rp_vld = _T_472; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 353:29:@5634.4]
  assign io_pixel_planar1_sft = _T_437; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 343:26:@5579.4]
  assign io_pixel_planar1_width_burst = _T_458; // @[NV_NVDLA_CDMA_IMG_ctrl.scala 349:34:@5612.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_117 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_163 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_156 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_169 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_166 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_142 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_197 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_153 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_412 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_415 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_418 = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_421 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_430 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_433 = _RAND_14[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_437 = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_440 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_444 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_447 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_451 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_454 = _RAND_20[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_458 = _RAND_21[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_461 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_465 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_468 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_472 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_476 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_479 = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_483 = _RAND_28[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_488 = _RAND_29[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_491 = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_495 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_498 = _RAND_32[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_502 = _RAND_33[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_117 <= 1'h0;
    end else begin
      if (_T_172) begin
        _T_117 <= _T_173;
      end
    end
    if (reset) begin
      _T_163 <= 5'h1f;
    end else begin
      if (_T_172) begin
        _T_163 <= io_reg2dp_data_bank;
      end
    end
    if (reset) begin
      _T_156 <= 1'h0;
    end else begin
      if (_T_172) begin
        _T_156 <= _T_219;
      end
    end
    if (reset) begin
      _T_169 <= 1'h0;
    end else begin
      _T_169 <= _T_166;
    end
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= io_sc2cdma_dat_pending_req;
    end
  end
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_129 <= 2'h0;
    end else begin
      if (_T_132) begin
        if (_T_133) begin
          _T_129 <= 2'h1;
        end else begin
          if (_T_136) begin
            _T_129 <= 2'h3;
          end else begin
            if (_T_219) begin
              _T_129 <= 2'h2;
            end else begin
              _T_129 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_137) begin
          if (_T_171) begin
            _T_129 <= 2'h2;
          end else begin
            _T_129 <= 2'h0;
          end
        end else begin
          if (_T_138) begin
            if (_T_204) begin
              _T_129 <= 2'h3;
            end else begin
              _T_129 <= 2'h0;
            end
          end else begin
            _T_129 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      _T_142 <= io_is_running;
    end
    if (reset) begin
      _T_197 <= 5'h0;
    end else begin
      _T_197 <= _GEN_15[4:0];
    end
    if (reset) begin
      _T_153 <= 2'h0;
    end else begin
      if (_T_132) begin
        if (_T_133) begin
          _T_153 <= 2'h1;
        end else begin
          if (_T_136) begin
            _T_153 <= 2'h3;
          end else begin
            if (_T_219) begin
              _T_153 <= 2'h2;
            end else begin
              _T_153 <= 2'h0;
            end
          end
        end
      end else begin
        if (_T_137) begin
          if (_T_171) begin
            _T_153 <= 2'h2;
          end else begin
            _T_153 <= 2'h0;
          end
        end else begin
          if (_T_138) begin
            if (_T_204) begin
              _T_153 <= 2'h3;
            end else begin
              _T_153 <= 2'h0;
            end
          end else begin
            _T_153 <= 2'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_412 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        if (_T_246) begin
          _T_412 <= 1'h0;
        end else begin
          if (_T_250) begin
            _T_412 <= 1'h0;
          end else begin
            if (_T_253) begin
              _T_412 <= 1'h0;
            end else begin
              if (_T_256) begin
                _T_412 <= 1'h0;
              end else begin
                if (_T_259) begin
                  _T_412 <= 1'h0;
                end else begin
                  if (_T_262) begin
                    _T_412 <= 1'h0;
                  end else begin
                    if (_T_265) begin
                      _T_412 <= 1'h0;
                    end else begin
                      if (_T_268) begin
                        _T_412 <= 1'h0;
                      end else begin
                        if (_T_271) begin
                          _T_412 <= 1'h0;
                        end else begin
                          if (_T_274) begin
                            _T_412 <= 1'h0;
                          end else begin
                            if (_T_277) begin
                              _T_412 <= 1'h0;
                            end else begin
                              if (_T_280) begin
                                _T_412 <= 1'h1;
                              end else begin
                                _T_412 <= _T_280;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_415 <= 2'h0;
    end else begin
      if (io_layer_st) begin
        _T_415 <= 2'h0;
      end
    end
    if (reset) begin
      _T_418 <= 11'h0;
    end else begin
      if (io_layer_st) begin
        if (_T_246) begin
          _T_418 <= 11'h1;
        end else begin
          if (_T_250) begin
            _T_418 <= 11'h1;
          end else begin
            if (_T_253) begin
              _T_418 <= 11'h2;
            end else begin
              if (_T_256) begin
                _T_418 <= 11'h8;
              end else begin
                if (_T_259) begin
                  _T_418 <= 11'h20;
                end else begin
                  if (_T_262) begin
                    _T_418 <= 11'h1;
                  end else begin
                    if (_T_265) begin
                      _T_418 <= 11'h2;
                    end else begin
                      if (_T_268) begin
                        _T_418 <= 11'h8;
                      end else begin
                        if (_T_271) begin
                          _T_418 <= 11'h20;
                        end else begin
                          if (_T_274) begin
                            _T_418 <= 11'h2;
                          end else begin
                            if (_T_277) begin
                              _T_418 <= 11'h8;
                            end else begin
                              if (_T_280) begin
                                _T_418 <= 11'h200;
                              end else begin
                                _T_418 <= 11'h1;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_421 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        _T_421 <= 1'h0;
      end
    end
    if (reset) begin
      _T_430 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        _T_430 <= _T_299;
      end
    end
    if (reset) begin
      _T_433 <= 3'h0;
    end else begin
      if (io_layer_st) begin
        if (_T_246) begin
          _T_433 <= 3'h5;
        end else begin
          if (_T_250) begin
            _T_433 <= 3'h3;
          end else begin
            if (_T_253) begin
              _T_433 <= 3'h3;
            end else begin
              if (_T_256) begin
                _T_433 <= 3'h3;
              end else begin
                if (_T_259) begin
                  _T_433 <= 3'h3;
                end else begin
                  if (_T_262) begin
                    _T_433 <= 3'h3;
                  end else begin
                    if (_T_265) begin
                      _T_433 <= 3'h3;
                    end else begin
                      if (_T_268) begin
                        _T_433 <= 3'h3;
                      end else begin
                        if (_T_271) begin
                          _T_433 <= 3'h3;
                        end else begin
                          if (_T_274) begin
                            _T_433 <= 3'h3;
                          end else begin
                            if (_T_277) begin
                              _T_433 <= 3'h3;
                            end else begin
                              if (_T_280) begin
                                _T_433 <= 3'h5;
                              end else begin
                                if (_T_280) begin
                                  _T_433 <= 3'h5;
                                end else begin
                                  _T_433 <= 3'h3;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_437 <= 3'h0;
    end else begin
      if (_T_435) begin
        if (_T_246) begin
          _T_437 <= 3'h3;
        end else begin
          if (_T_250) begin
            _T_437 <= 3'h3;
          end else begin
            if (_T_253) begin
              _T_437 <= 3'h3;
            end else begin
              if (_T_256) begin
                _T_437 <= 3'h3;
              end else begin
                if (_T_259) begin
                  _T_437 <= 3'h3;
                end else begin
                  if (_T_262) begin
                    _T_437 <= 3'h3;
                  end else begin
                    if (_T_265) begin
                      _T_437 <= 3'h3;
                    end else begin
                      if (_T_268) begin
                        _T_437 <= 3'h3;
                      end else begin
                        if (_T_271) begin
                          _T_437 <= 3'h3;
                        end else begin
                          if (_T_274) begin
                            _T_437 <= 3'h3;
                          end else begin
                            if (_T_277) begin
                              _T_437 <= 3'h3;
                            end else begin
                              if (_T_280) begin
                                _T_437 <= 3'h4;
                              end else begin
                                if (_T_280) begin
                                  _T_437 <= 3'h4;
                                end else begin
                                  _T_437 <= 3'h3;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_440 <= 4'h0;
    end else begin
      if (io_layer_st) begin
        _T_440 <= _T_309;
      end
    end
    if (reset) begin
      _T_444 <= 3'h0;
    end else begin
      if (_T_435) begin
        _T_444 <= _T_316;
      end
    end
    if (reset) begin
      _T_447 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        _T_447 <= _T_403;
      end
    end
    if (reset) begin
      _T_451 <= 1'h0;
    end else begin
      if (_T_435) begin
        _T_451 <= _T_405;
      end
    end
    if (reset) begin
      _T_454 <= 14'h0;
    end else begin
      _T_454 <= _GEN_106[13:0];
    end
    if (reset) begin
      _T_458 <= 14'h0;
    end else begin
      _T_458 <= _GEN_107[13:0];
    end
    if (reset) begin
      _T_461 <= 4'h0;
    end else begin
      if (io_layer_st) begin
        _T_461 <= _T_337;
      end
    end
    if (reset) begin
      _T_465 <= 3'h0;
    end else begin
      if (_T_435) begin
        _T_465 <= _T_342;
      end
    end
    if (reset) begin
      _T_468 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        _T_468 <= _T_407;
      end
    end
    if (reset) begin
      _T_472 <= 1'h0;
    end else begin
      if (_T_435) begin
        _T_472 <= _T_409;
      end
    end
    if (reset) begin
      _T_476 <= 1'h0;
    end else begin
      if (_T_435) begin
        _T_476 <= _T_376;
      end
    end
    if (reset) begin
      _T_479 <= 5'h0;
    end else begin
      if (io_layer_st) begin
        _T_479 <= _T_388;
      end
    end
    if (reset) begin
      _T_483 <= 5'h0;
    end else begin
      if (_T_435) begin
        _T_483 <= _T_396;
      end
    end
    if (reset) begin
      _T_488 <= 6'h0;
    end else begin
      if (io_layer_st) begin
        _T_488 <= _T_485;
      end
    end
    if (reset) begin
      _T_491 <= 4'h0;
    end else begin
      if (io_layer_st) begin
        _T_491 <= 4'h8;
      end
    end
    if (reset) begin
      _T_495 <= 5'h0;
    end else begin
      if (_T_435) begin
        _T_495 <= 5'h10;
      end
    end
    if (reset) begin
      _T_498 <= 4'h0;
    end else begin
      if (io_layer_st) begin
        _T_498 <= 4'h9;
      end
    end
    if (reset) begin
      _T_502 <= 5'h0;
    end else begin
      if (_T_435) begin
        _T_502 <= 5'h11;
      end
    end
  end
endmodule
module nv_ram_rwsp_3( // @[:@6026.2]
  input         io_clk, // @[:@6029.4]
  input         io_re, // @[:@6029.4]
  input         io_we, // @[:@6029.4]
  input         io_ore, // @[:@6029.4]
  input  [6:0]  io_ra, // @[:@6029.4]
  input  [6:0]  io_wa, // @[:@6029.4]
  input  [10:0] io_di, // @[:@6029.4]
  output [10:0] io_dout // @[:@6029.4]
);
  reg [10:0] _T_26_0; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_0;
  reg [10:0] _T_26_1; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_1;
  reg [10:0] _T_26_2; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_2;
  reg [10:0] _T_26_3; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_3;
  reg [10:0] _T_26_4; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_4;
  reg [10:0] _T_26_5; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_5;
  reg [10:0] _T_26_6; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_6;
  reg [10:0] _T_26_7; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_7;
  reg [10:0] _T_26_8; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_8;
  reg [10:0] _T_26_9; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_9;
  reg [10:0] _T_26_10; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_10;
  reg [10:0] _T_26_11; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_11;
  reg [10:0] _T_26_12; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_12;
  reg [10:0] _T_26_13; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_13;
  reg [10:0] _T_26_14; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_14;
  reg [10:0] _T_26_15; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_15;
  reg [10:0] _T_26_16; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_16;
  reg [10:0] _T_26_17; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_17;
  reg [10:0] _T_26_18; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_18;
  reg [10:0] _T_26_19; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_19;
  reg [10:0] _T_26_20; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_20;
  reg [10:0] _T_26_21; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_21;
  reg [10:0] _T_26_22; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_22;
  reg [10:0] _T_26_23; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_23;
  reg [10:0] _T_26_24; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_24;
  reg [10:0] _T_26_25; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_25;
  reg [10:0] _T_26_26; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_26;
  reg [10:0] _T_26_27; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_27;
  reg [10:0] _T_26_28; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_28;
  reg [10:0] _T_26_29; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_29;
  reg [10:0] _T_26_30; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_30;
  reg [10:0] _T_26_31; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_31;
  reg [10:0] _T_26_32; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_32;
  reg [10:0] _T_26_33; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_33;
  reg [10:0] _T_26_34; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_34;
  reg [10:0] _T_26_35; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_35;
  reg [10:0] _T_26_36; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_36;
  reg [10:0] _T_26_37; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_37;
  reg [10:0] _T_26_38; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_38;
  reg [10:0] _T_26_39; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_39;
  reg [10:0] _T_26_40; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_40;
  reg [10:0] _T_26_41; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_41;
  reg [10:0] _T_26_42; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_42;
  reg [10:0] _T_26_43; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_43;
  reg [10:0] _T_26_44; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_44;
  reg [10:0] _T_26_45; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_45;
  reg [10:0] _T_26_46; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_46;
  reg [10:0] _T_26_47; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_47;
  reg [10:0] _T_26_48; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_48;
  reg [10:0] _T_26_49; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_49;
  reg [10:0] _T_26_50; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_50;
  reg [10:0] _T_26_51; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_51;
  reg [10:0] _T_26_52; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_52;
  reg [10:0] _T_26_53; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_53;
  reg [10:0] _T_26_54; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_54;
  reg [10:0] _T_26_55; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_55;
  reg [10:0] _T_26_56; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_56;
  reg [10:0] _T_26_57; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_57;
  reg [10:0] _T_26_58; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_58;
  reg [10:0] _T_26_59; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_59;
  reg [10:0] _T_26_60; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_60;
  reg [10:0] _T_26_61; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_61;
  reg [10:0] _T_26_62; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_62;
  reg [10:0] _T_26_63; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_63;
  reg [10:0] _T_26_64; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_64;
  reg [10:0] _T_26_65; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_65;
  reg [10:0] _T_26_66; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_66;
  reg [10:0] _T_26_67; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_67;
  reg [10:0] _T_26_68; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_68;
  reg [10:0] _T_26_69; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_69;
  reg [10:0] _T_26_70; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_70;
  reg [10:0] _T_26_71; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_71;
  reg [10:0] _T_26_72; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_72;
  reg [10:0] _T_26_73; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_73;
  reg [10:0] _T_26_74; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_74;
  reg [10:0] _T_26_75; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_75;
  reg [10:0] _T_26_76; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_76;
  reg [10:0] _T_26_77; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_77;
  reg [10:0] _T_26_78; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_78;
  reg [10:0] _T_26_79; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_79;
  reg [10:0] _T_26_80; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_80;
  reg [10:0] _T_26_81; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_81;
  reg [10:0] _T_26_82; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_82;
  reg [10:0] _T_26_83; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_83;
  reg [10:0] _T_26_84; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_84;
  reg [10:0] _T_26_85; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_85;
  reg [10:0] _T_26_86; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_86;
  reg [10:0] _T_26_87; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_87;
  reg [10:0] _T_26_88; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_88;
  reg [10:0] _T_26_89; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_89;
  reg [10:0] _T_26_90; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_90;
  reg [10:0] _T_26_91; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_91;
  reg [10:0] _T_26_92; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_92;
  reg [10:0] _T_26_93; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_93;
  reg [10:0] _T_26_94; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_94;
  reg [10:0] _T_26_95; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_95;
  reg [10:0] _T_26_96; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_96;
  reg [10:0] _T_26_97; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_97;
  reg [10:0] _T_26_98; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_98;
  reg [10:0] _T_26_99; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_99;
  reg [10:0] _T_26_100; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_100;
  reg [10:0] _T_26_101; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_101;
  reg [10:0] _T_26_102; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_102;
  reg [10:0] _T_26_103; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_103;
  reg [10:0] _T_26_104; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_104;
  reg [10:0] _T_26_105; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_105;
  reg [10:0] _T_26_106; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_106;
  reg [10:0] _T_26_107; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_107;
  reg [10:0] _T_26_108; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_108;
  reg [10:0] _T_26_109; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_109;
  reg [10:0] _T_26_110; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_110;
  reg [10:0] _T_26_111; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_111;
  reg [10:0] _T_26_112; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_112;
  reg [10:0] _T_26_113; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_113;
  reg [10:0] _T_26_114; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_114;
  reg [10:0] _T_26_115; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_115;
  reg [10:0] _T_26_116; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_116;
  reg [10:0] _T_26_117; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_117;
  reg [10:0] _T_26_118; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_118;
  reg [10:0] _T_26_119; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_119;
  reg [10:0] _T_26_120; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_120;
  reg [10:0] _T_26_121; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_121;
  reg [10:0] _T_26_122; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_122;
  reg [10:0] _T_26_123; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_123;
  reg [10:0] _T_26_124; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_124;
  reg [10:0] _T_26_125; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_125;
  reg [10:0] _T_26_126; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_126;
  reg [10:0] _T_26_127; // @[nv_ram_rwsp.scala 31:18:@6031.4]
  reg [31:0] _RAND_127;
  reg [6:0] _T_158; // @[nv_ram_rwsp.scala 32:19:@6032.4]
  reg [31:0] _RAND_128;
  reg [10:0] _T_160; // @[nv_ram_rwsp.scala 33:21:@6033.4]
  reg [31:0] _RAND_129;
  wire [10:0] _GEN_0; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_1; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_2; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_3; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_4; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_5; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_6; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_7; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_8; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_9; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_10; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_11; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_12; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_13; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_14; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_15; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_16; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_17; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_18; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_19; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_20; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_21; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_22; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_23; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_24; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_25; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_26; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_27; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_28; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_29; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_30; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_31; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_32; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_33; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_34; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_35; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_36; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_37; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_38; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_39; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_40; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_41; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_42; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_43; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_44; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_45; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_46; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_47; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_48; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_49; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_50; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_51; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_52; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_53; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_54; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_55; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_56; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_57; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_58; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_59; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_60; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_61; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_62; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_63; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_64; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_65; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_66; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_67; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_68; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_69; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_70; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_71; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_72; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_73; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_74; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_75; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_76; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_77; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_78; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_79; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_80; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_81; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_82; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_83; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_84; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_85; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_86; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_87; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_88; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_89; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_90; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_91; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_92; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_93; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_94; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_95; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_96; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_97; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_98; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_99; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_100; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_101; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_102; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_103; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_104; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_105; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_106; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_107; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_108; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_109; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_110; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_111; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_112; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_113; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_114; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_115; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_116; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_117; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_118; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_119; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_120; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_121; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_122; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_123; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_124; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_125; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_126; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_127; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  wire [10:0] _GEN_258; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_259; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_260; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_261; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_262; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_263; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_264; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_265; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_266; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_267; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_268; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_269; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_270; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_271; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_272; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_273; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_274; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_275; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_276; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_277; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_278; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_279; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_280; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_281; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_282; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_283; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_284; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_285; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_286; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_287; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_288; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_289; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_290; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_291; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_292; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_293; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_294; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_295; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_296; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_297; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_298; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_299; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_300; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_301; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_302; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_303; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_304; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_305; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_306; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_307; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_308; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_309; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_310; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_311; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_312; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_313; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_314; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_315; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_316; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_317; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_318; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_319; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_320; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_321; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_322; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_323; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_324; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_325; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_326; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_327; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_328; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_329; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_330; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_331; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_332; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_333; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_334; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_335; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_336; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_337; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_338; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_339; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_340; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_341; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_342; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_343; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_344; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_345; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_346; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_347; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_348; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_349; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_350; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_351; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_352; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_353; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_354; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_355; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_356; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_357; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_358; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_359; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_360; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_361; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_362; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_363; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_364; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_365; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_366; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_367; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_368; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_369; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_370; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_371; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_372; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_373; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_374; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_375; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_376; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_377; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_378; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_379; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_380; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_381; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_382; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_383; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  wire [10:0] _GEN_384; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_0 = 7'h0 == io_wa ? io_di : _T_26_0; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_1 = 7'h1 == io_wa ? io_di : _T_26_1; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_2 = 7'h2 == io_wa ? io_di : _T_26_2; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_3 = 7'h3 == io_wa ? io_di : _T_26_3; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_4 = 7'h4 == io_wa ? io_di : _T_26_4; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_5 = 7'h5 == io_wa ? io_di : _T_26_5; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_6 = 7'h6 == io_wa ? io_di : _T_26_6; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_7 = 7'h7 == io_wa ? io_di : _T_26_7; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_8 = 7'h8 == io_wa ? io_di : _T_26_8; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_9 = 7'h9 == io_wa ? io_di : _T_26_9; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_10 = 7'ha == io_wa ? io_di : _T_26_10; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_11 = 7'hb == io_wa ? io_di : _T_26_11; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_12 = 7'hc == io_wa ? io_di : _T_26_12; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_13 = 7'hd == io_wa ? io_di : _T_26_13; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_14 = 7'he == io_wa ? io_di : _T_26_14; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_15 = 7'hf == io_wa ? io_di : _T_26_15; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_16 = 7'h10 == io_wa ? io_di : _T_26_16; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_17 = 7'h11 == io_wa ? io_di : _T_26_17; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_18 = 7'h12 == io_wa ? io_di : _T_26_18; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_19 = 7'h13 == io_wa ? io_di : _T_26_19; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_20 = 7'h14 == io_wa ? io_di : _T_26_20; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_21 = 7'h15 == io_wa ? io_di : _T_26_21; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_22 = 7'h16 == io_wa ? io_di : _T_26_22; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_23 = 7'h17 == io_wa ? io_di : _T_26_23; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_24 = 7'h18 == io_wa ? io_di : _T_26_24; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_25 = 7'h19 == io_wa ? io_di : _T_26_25; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_26 = 7'h1a == io_wa ? io_di : _T_26_26; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_27 = 7'h1b == io_wa ? io_di : _T_26_27; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_28 = 7'h1c == io_wa ? io_di : _T_26_28; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_29 = 7'h1d == io_wa ? io_di : _T_26_29; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_30 = 7'h1e == io_wa ? io_di : _T_26_30; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_31 = 7'h1f == io_wa ? io_di : _T_26_31; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_32 = 7'h20 == io_wa ? io_di : _T_26_32; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_33 = 7'h21 == io_wa ? io_di : _T_26_33; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_34 = 7'h22 == io_wa ? io_di : _T_26_34; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_35 = 7'h23 == io_wa ? io_di : _T_26_35; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_36 = 7'h24 == io_wa ? io_di : _T_26_36; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_37 = 7'h25 == io_wa ? io_di : _T_26_37; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_38 = 7'h26 == io_wa ? io_di : _T_26_38; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_39 = 7'h27 == io_wa ? io_di : _T_26_39; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_40 = 7'h28 == io_wa ? io_di : _T_26_40; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_41 = 7'h29 == io_wa ? io_di : _T_26_41; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_42 = 7'h2a == io_wa ? io_di : _T_26_42; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_43 = 7'h2b == io_wa ? io_di : _T_26_43; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_44 = 7'h2c == io_wa ? io_di : _T_26_44; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_45 = 7'h2d == io_wa ? io_di : _T_26_45; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_46 = 7'h2e == io_wa ? io_di : _T_26_46; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_47 = 7'h2f == io_wa ? io_di : _T_26_47; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_48 = 7'h30 == io_wa ? io_di : _T_26_48; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_49 = 7'h31 == io_wa ? io_di : _T_26_49; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_50 = 7'h32 == io_wa ? io_di : _T_26_50; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_51 = 7'h33 == io_wa ? io_di : _T_26_51; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_52 = 7'h34 == io_wa ? io_di : _T_26_52; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_53 = 7'h35 == io_wa ? io_di : _T_26_53; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_54 = 7'h36 == io_wa ? io_di : _T_26_54; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_55 = 7'h37 == io_wa ? io_di : _T_26_55; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_56 = 7'h38 == io_wa ? io_di : _T_26_56; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_57 = 7'h39 == io_wa ? io_di : _T_26_57; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_58 = 7'h3a == io_wa ? io_di : _T_26_58; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_59 = 7'h3b == io_wa ? io_di : _T_26_59; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_60 = 7'h3c == io_wa ? io_di : _T_26_60; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_61 = 7'h3d == io_wa ? io_di : _T_26_61; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_62 = 7'h3e == io_wa ? io_di : _T_26_62; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_63 = 7'h3f == io_wa ? io_di : _T_26_63; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_64 = 7'h40 == io_wa ? io_di : _T_26_64; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_65 = 7'h41 == io_wa ? io_di : _T_26_65; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_66 = 7'h42 == io_wa ? io_di : _T_26_66; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_67 = 7'h43 == io_wa ? io_di : _T_26_67; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_68 = 7'h44 == io_wa ? io_di : _T_26_68; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_69 = 7'h45 == io_wa ? io_di : _T_26_69; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_70 = 7'h46 == io_wa ? io_di : _T_26_70; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_71 = 7'h47 == io_wa ? io_di : _T_26_71; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_72 = 7'h48 == io_wa ? io_di : _T_26_72; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_73 = 7'h49 == io_wa ? io_di : _T_26_73; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_74 = 7'h4a == io_wa ? io_di : _T_26_74; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_75 = 7'h4b == io_wa ? io_di : _T_26_75; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_76 = 7'h4c == io_wa ? io_di : _T_26_76; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_77 = 7'h4d == io_wa ? io_di : _T_26_77; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_78 = 7'h4e == io_wa ? io_di : _T_26_78; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_79 = 7'h4f == io_wa ? io_di : _T_26_79; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_80 = 7'h50 == io_wa ? io_di : _T_26_80; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_81 = 7'h51 == io_wa ? io_di : _T_26_81; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_82 = 7'h52 == io_wa ? io_di : _T_26_82; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_83 = 7'h53 == io_wa ? io_di : _T_26_83; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_84 = 7'h54 == io_wa ? io_di : _T_26_84; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_85 = 7'h55 == io_wa ? io_di : _T_26_85; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_86 = 7'h56 == io_wa ? io_di : _T_26_86; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_87 = 7'h57 == io_wa ? io_di : _T_26_87; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_88 = 7'h58 == io_wa ? io_di : _T_26_88; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_89 = 7'h59 == io_wa ? io_di : _T_26_89; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_90 = 7'h5a == io_wa ? io_di : _T_26_90; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_91 = 7'h5b == io_wa ? io_di : _T_26_91; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_92 = 7'h5c == io_wa ? io_di : _T_26_92; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_93 = 7'h5d == io_wa ? io_di : _T_26_93; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_94 = 7'h5e == io_wa ? io_di : _T_26_94; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_95 = 7'h5f == io_wa ? io_di : _T_26_95; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_96 = 7'h60 == io_wa ? io_di : _T_26_96; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_97 = 7'h61 == io_wa ? io_di : _T_26_97; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_98 = 7'h62 == io_wa ? io_di : _T_26_98; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_99 = 7'h63 == io_wa ? io_di : _T_26_99; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_100 = 7'h64 == io_wa ? io_di : _T_26_100; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_101 = 7'h65 == io_wa ? io_di : _T_26_101; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_102 = 7'h66 == io_wa ? io_di : _T_26_102; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_103 = 7'h67 == io_wa ? io_di : _T_26_103; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_104 = 7'h68 == io_wa ? io_di : _T_26_104; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_105 = 7'h69 == io_wa ? io_di : _T_26_105; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_106 = 7'h6a == io_wa ? io_di : _T_26_106; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_107 = 7'h6b == io_wa ? io_di : _T_26_107; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_108 = 7'h6c == io_wa ? io_di : _T_26_108; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_109 = 7'h6d == io_wa ? io_di : _T_26_109; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_110 = 7'h6e == io_wa ? io_di : _T_26_110; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_111 = 7'h6f == io_wa ? io_di : _T_26_111; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_112 = 7'h70 == io_wa ? io_di : _T_26_112; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_113 = 7'h71 == io_wa ? io_di : _T_26_113; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_114 = 7'h72 == io_wa ? io_di : _T_26_114; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_115 = 7'h73 == io_wa ? io_di : _T_26_115; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_116 = 7'h74 == io_wa ? io_di : _T_26_116; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_117 = 7'h75 == io_wa ? io_di : _T_26_117; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_118 = 7'h76 == io_wa ? io_di : _T_26_118; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_119 = 7'h77 == io_wa ? io_di : _T_26_119; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_120 = 7'h78 == io_wa ? io_di : _T_26_120; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_121 = 7'h79 == io_wa ? io_di : _T_26_121; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_122 = 7'h7a == io_wa ? io_di : _T_26_122; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_123 = 7'h7b == io_wa ? io_di : _T_26_123; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_124 = 7'h7c == io_wa ? io_di : _T_26_124; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_125 = 7'h7d == io_wa ? io_di : _T_26_125; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_126 = 7'h7e == io_wa ? io_di : _T_26_126; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_127 = 7'h7f == io_wa ? io_di : _T_26_127; // @[nv_ram_rwsp.scala 36:20:@6035.6]
  assign _GEN_258 = 7'h1 == _T_158 ? _T_26_1 : _T_26_0; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_259 = 7'h2 == _T_158 ? _T_26_2 : _GEN_258; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_260 = 7'h3 == _T_158 ? _T_26_3 : _GEN_259; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_261 = 7'h4 == _T_158 ? _T_26_4 : _GEN_260; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_262 = 7'h5 == _T_158 ? _T_26_5 : _GEN_261; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_263 = 7'h6 == _T_158 ? _T_26_6 : _GEN_262; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_264 = 7'h7 == _T_158 ? _T_26_7 : _GEN_263; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_265 = 7'h8 == _T_158 ? _T_26_8 : _GEN_264; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_266 = 7'h9 == _T_158 ? _T_26_9 : _GEN_265; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_267 = 7'ha == _T_158 ? _T_26_10 : _GEN_266; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_268 = 7'hb == _T_158 ? _T_26_11 : _GEN_267; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_269 = 7'hc == _T_158 ? _T_26_12 : _GEN_268; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_270 = 7'hd == _T_158 ? _T_26_13 : _GEN_269; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_271 = 7'he == _T_158 ? _T_26_14 : _GEN_270; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_272 = 7'hf == _T_158 ? _T_26_15 : _GEN_271; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_273 = 7'h10 == _T_158 ? _T_26_16 : _GEN_272; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_274 = 7'h11 == _T_158 ? _T_26_17 : _GEN_273; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_275 = 7'h12 == _T_158 ? _T_26_18 : _GEN_274; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_276 = 7'h13 == _T_158 ? _T_26_19 : _GEN_275; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_277 = 7'h14 == _T_158 ? _T_26_20 : _GEN_276; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_278 = 7'h15 == _T_158 ? _T_26_21 : _GEN_277; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_279 = 7'h16 == _T_158 ? _T_26_22 : _GEN_278; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_280 = 7'h17 == _T_158 ? _T_26_23 : _GEN_279; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_281 = 7'h18 == _T_158 ? _T_26_24 : _GEN_280; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_282 = 7'h19 == _T_158 ? _T_26_25 : _GEN_281; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_283 = 7'h1a == _T_158 ? _T_26_26 : _GEN_282; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_284 = 7'h1b == _T_158 ? _T_26_27 : _GEN_283; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_285 = 7'h1c == _T_158 ? _T_26_28 : _GEN_284; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_286 = 7'h1d == _T_158 ? _T_26_29 : _GEN_285; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_287 = 7'h1e == _T_158 ? _T_26_30 : _GEN_286; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_288 = 7'h1f == _T_158 ? _T_26_31 : _GEN_287; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_289 = 7'h20 == _T_158 ? _T_26_32 : _GEN_288; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_290 = 7'h21 == _T_158 ? _T_26_33 : _GEN_289; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_291 = 7'h22 == _T_158 ? _T_26_34 : _GEN_290; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_292 = 7'h23 == _T_158 ? _T_26_35 : _GEN_291; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_293 = 7'h24 == _T_158 ? _T_26_36 : _GEN_292; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_294 = 7'h25 == _T_158 ? _T_26_37 : _GEN_293; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_295 = 7'h26 == _T_158 ? _T_26_38 : _GEN_294; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_296 = 7'h27 == _T_158 ? _T_26_39 : _GEN_295; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_297 = 7'h28 == _T_158 ? _T_26_40 : _GEN_296; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_298 = 7'h29 == _T_158 ? _T_26_41 : _GEN_297; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_299 = 7'h2a == _T_158 ? _T_26_42 : _GEN_298; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_300 = 7'h2b == _T_158 ? _T_26_43 : _GEN_299; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_301 = 7'h2c == _T_158 ? _T_26_44 : _GEN_300; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_302 = 7'h2d == _T_158 ? _T_26_45 : _GEN_301; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_303 = 7'h2e == _T_158 ? _T_26_46 : _GEN_302; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_304 = 7'h2f == _T_158 ? _T_26_47 : _GEN_303; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_305 = 7'h30 == _T_158 ? _T_26_48 : _GEN_304; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_306 = 7'h31 == _T_158 ? _T_26_49 : _GEN_305; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_307 = 7'h32 == _T_158 ? _T_26_50 : _GEN_306; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_308 = 7'h33 == _T_158 ? _T_26_51 : _GEN_307; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_309 = 7'h34 == _T_158 ? _T_26_52 : _GEN_308; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_310 = 7'h35 == _T_158 ? _T_26_53 : _GEN_309; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_311 = 7'h36 == _T_158 ? _T_26_54 : _GEN_310; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_312 = 7'h37 == _T_158 ? _T_26_55 : _GEN_311; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_313 = 7'h38 == _T_158 ? _T_26_56 : _GEN_312; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_314 = 7'h39 == _T_158 ? _T_26_57 : _GEN_313; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_315 = 7'h3a == _T_158 ? _T_26_58 : _GEN_314; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_316 = 7'h3b == _T_158 ? _T_26_59 : _GEN_315; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_317 = 7'h3c == _T_158 ? _T_26_60 : _GEN_316; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_318 = 7'h3d == _T_158 ? _T_26_61 : _GEN_317; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_319 = 7'h3e == _T_158 ? _T_26_62 : _GEN_318; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_320 = 7'h3f == _T_158 ? _T_26_63 : _GEN_319; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_321 = 7'h40 == _T_158 ? _T_26_64 : _GEN_320; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_322 = 7'h41 == _T_158 ? _T_26_65 : _GEN_321; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_323 = 7'h42 == _T_158 ? _T_26_66 : _GEN_322; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_324 = 7'h43 == _T_158 ? _T_26_67 : _GEN_323; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_325 = 7'h44 == _T_158 ? _T_26_68 : _GEN_324; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_326 = 7'h45 == _T_158 ? _T_26_69 : _GEN_325; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_327 = 7'h46 == _T_158 ? _T_26_70 : _GEN_326; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_328 = 7'h47 == _T_158 ? _T_26_71 : _GEN_327; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_329 = 7'h48 == _T_158 ? _T_26_72 : _GEN_328; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_330 = 7'h49 == _T_158 ? _T_26_73 : _GEN_329; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_331 = 7'h4a == _T_158 ? _T_26_74 : _GEN_330; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_332 = 7'h4b == _T_158 ? _T_26_75 : _GEN_331; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_333 = 7'h4c == _T_158 ? _T_26_76 : _GEN_332; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_334 = 7'h4d == _T_158 ? _T_26_77 : _GEN_333; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_335 = 7'h4e == _T_158 ? _T_26_78 : _GEN_334; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_336 = 7'h4f == _T_158 ? _T_26_79 : _GEN_335; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_337 = 7'h50 == _T_158 ? _T_26_80 : _GEN_336; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_338 = 7'h51 == _T_158 ? _T_26_81 : _GEN_337; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_339 = 7'h52 == _T_158 ? _T_26_82 : _GEN_338; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_340 = 7'h53 == _T_158 ? _T_26_83 : _GEN_339; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_341 = 7'h54 == _T_158 ? _T_26_84 : _GEN_340; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_342 = 7'h55 == _T_158 ? _T_26_85 : _GEN_341; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_343 = 7'h56 == _T_158 ? _T_26_86 : _GEN_342; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_344 = 7'h57 == _T_158 ? _T_26_87 : _GEN_343; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_345 = 7'h58 == _T_158 ? _T_26_88 : _GEN_344; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_346 = 7'h59 == _T_158 ? _T_26_89 : _GEN_345; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_347 = 7'h5a == _T_158 ? _T_26_90 : _GEN_346; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_348 = 7'h5b == _T_158 ? _T_26_91 : _GEN_347; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_349 = 7'h5c == _T_158 ? _T_26_92 : _GEN_348; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_350 = 7'h5d == _T_158 ? _T_26_93 : _GEN_349; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_351 = 7'h5e == _T_158 ? _T_26_94 : _GEN_350; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_352 = 7'h5f == _T_158 ? _T_26_95 : _GEN_351; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_353 = 7'h60 == _T_158 ? _T_26_96 : _GEN_352; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_354 = 7'h61 == _T_158 ? _T_26_97 : _GEN_353; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_355 = 7'h62 == _T_158 ? _T_26_98 : _GEN_354; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_356 = 7'h63 == _T_158 ? _T_26_99 : _GEN_355; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_357 = 7'h64 == _T_158 ? _T_26_100 : _GEN_356; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_358 = 7'h65 == _T_158 ? _T_26_101 : _GEN_357; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_359 = 7'h66 == _T_158 ? _T_26_102 : _GEN_358; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_360 = 7'h67 == _T_158 ? _T_26_103 : _GEN_359; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_361 = 7'h68 == _T_158 ? _T_26_104 : _GEN_360; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_362 = 7'h69 == _T_158 ? _T_26_105 : _GEN_361; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_363 = 7'h6a == _T_158 ? _T_26_106 : _GEN_362; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_364 = 7'h6b == _T_158 ? _T_26_107 : _GEN_363; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_365 = 7'h6c == _T_158 ? _T_26_108 : _GEN_364; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_366 = 7'h6d == _T_158 ? _T_26_109 : _GEN_365; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_367 = 7'h6e == _T_158 ? _T_26_110 : _GEN_366; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_368 = 7'h6f == _T_158 ? _T_26_111 : _GEN_367; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_369 = 7'h70 == _T_158 ? _T_26_112 : _GEN_368; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_370 = 7'h71 == _T_158 ? _T_26_113 : _GEN_369; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_371 = 7'h72 == _T_158 ? _T_26_114 : _GEN_370; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_372 = 7'h73 == _T_158 ? _T_26_115 : _GEN_371; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_373 = 7'h74 == _T_158 ? _T_26_116 : _GEN_372; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_374 = 7'h75 == _T_158 ? _T_26_117 : _GEN_373; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_375 = 7'h76 == _T_158 ? _T_26_118 : _GEN_374; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_376 = 7'h77 == _T_158 ? _T_26_119 : _GEN_375; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_377 = 7'h78 == _T_158 ? _T_26_120 : _GEN_376; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_378 = 7'h79 == _T_158 ? _T_26_121 : _GEN_377; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_379 = 7'h7a == _T_158 ? _T_26_122 : _GEN_378; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_380 = 7'h7b == _T_158 ? _T_26_123 : _GEN_379; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_381 = 7'h7c == _T_158 ? _T_26_124 : _GEN_380; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_382 = 7'h7d == _T_158 ? _T_26_125 : _GEN_381; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_383 = 7'h7e == _T_158 ? _T_26_126 : _GEN_382; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign _GEN_384 = 7'h7f == _T_158 ? _T_26_127 : _GEN_383; // @[nv_ram_rwsp.scala 43:16:@6041.6]
  assign io_dout = _T_160; // @[nv_ram_rwsp.scala 45:13:@6043.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26_0 = _RAND_0[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26_1 = _RAND_1[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_26_2 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_26_3 = _RAND_3[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_26_4 = _RAND_4[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_26_5 = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_26_6 = _RAND_6[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_26_7 = _RAND_7[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_26_8 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_26_9 = _RAND_9[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_26_10 = _RAND_10[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_26_11 = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_26_12 = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_26_13 = _RAND_13[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_26_14 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_26_15 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_26_16 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_26_17 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_26_18 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_26_19 = _RAND_19[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_26_20 = _RAND_20[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_26_21 = _RAND_21[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_26_22 = _RAND_22[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_26_23 = _RAND_23[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_26_24 = _RAND_24[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_26_25 = _RAND_25[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26_26 = _RAND_26[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_26_27 = _RAND_27[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_26_28 = _RAND_28[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_26_29 = _RAND_29[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_26_30 = _RAND_30[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_26_31 = _RAND_31[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_26_32 = _RAND_32[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_26_33 = _RAND_33[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_26_34 = _RAND_34[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_26_35 = _RAND_35[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_26_36 = _RAND_36[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_26_37 = _RAND_37[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_26_38 = _RAND_38[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_26_39 = _RAND_39[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_26_40 = _RAND_40[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_26_41 = _RAND_41[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_26_42 = _RAND_42[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_26_43 = _RAND_43[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_26_44 = _RAND_44[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_26_45 = _RAND_45[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_26_46 = _RAND_46[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_26_47 = _RAND_47[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_26_48 = _RAND_48[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_26_49 = _RAND_49[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_26_50 = _RAND_50[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_26_51 = _RAND_51[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_26_52 = _RAND_52[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_26_53 = _RAND_53[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_26_54 = _RAND_54[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_26_55 = _RAND_55[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_26_56 = _RAND_56[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_26_57 = _RAND_57[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_26_58 = _RAND_58[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_26_59 = _RAND_59[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_26_60 = _RAND_60[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_26_61 = _RAND_61[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_26_62 = _RAND_62[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_26_63 = _RAND_63[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_26_64 = _RAND_64[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_26_65 = _RAND_65[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_26_66 = _RAND_66[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_26_67 = _RAND_67[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_26_68 = _RAND_68[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_26_69 = _RAND_69[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_26_70 = _RAND_70[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_26_71 = _RAND_71[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_26_72 = _RAND_72[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_26_73 = _RAND_73[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_26_74 = _RAND_74[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_26_75 = _RAND_75[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_26_76 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_26_77 = _RAND_77[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_26_78 = _RAND_78[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_26_79 = _RAND_79[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_26_80 = _RAND_80[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_26_81 = _RAND_81[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_26_82 = _RAND_82[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_26_83 = _RAND_83[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_26_84 = _RAND_84[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_26_85 = _RAND_85[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_26_86 = _RAND_86[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_26_87 = _RAND_87[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_26_88 = _RAND_88[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_26_89 = _RAND_89[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_26_90 = _RAND_90[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_26_91 = _RAND_91[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_26_92 = _RAND_92[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_26_93 = _RAND_93[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_26_94 = _RAND_94[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_26_95 = _RAND_95[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_26_96 = _RAND_96[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_26_97 = _RAND_97[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_26_98 = _RAND_98[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_26_99 = _RAND_99[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_26_100 = _RAND_100[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_26_101 = _RAND_101[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_26_102 = _RAND_102[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_26_103 = _RAND_103[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_26_104 = _RAND_104[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_26_105 = _RAND_105[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_26_106 = _RAND_106[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_26_107 = _RAND_107[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_26_108 = _RAND_108[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_26_109 = _RAND_109[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_26_110 = _RAND_110[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_26_111 = _RAND_111[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_26_112 = _RAND_112[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_26_113 = _RAND_113[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_26_114 = _RAND_114[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_26_115 = _RAND_115[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_26_116 = _RAND_116[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_26_117 = _RAND_117[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_26_118 = _RAND_118[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_26_119 = _RAND_119[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_26_120 = _RAND_120[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_26_121 = _RAND_121[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_26_122 = _RAND_122[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_26_123 = _RAND_123[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_26_124 = _RAND_124[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_26_125 = _RAND_125[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_26_126 = _RAND_126[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_26_127 = _RAND_127[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_158 = _RAND_128[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_160 = _RAND_129[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (7'h0 == io_wa) begin
        _T_26_0 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1 == io_wa) begin
        _T_26_1 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2 == io_wa) begin
        _T_26_2 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3 == io_wa) begin
        _T_26_3 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4 == io_wa) begin
        _T_26_4 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5 == io_wa) begin
        _T_26_5 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6 == io_wa) begin
        _T_26_6 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7 == io_wa) begin
        _T_26_7 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h8 == io_wa) begin
        _T_26_8 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h9 == io_wa) begin
        _T_26_9 <= io_di;
      end
    end
    if (io_we) begin
      if (7'ha == io_wa) begin
        _T_26_10 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hb == io_wa) begin
        _T_26_11 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hc == io_wa) begin
        _T_26_12 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hd == io_wa) begin
        _T_26_13 <= io_di;
      end
    end
    if (io_we) begin
      if (7'he == io_wa) begin
        _T_26_14 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hf == io_wa) begin
        _T_26_15 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h10 == io_wa) begin
        _T_26_16 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h11 == io_wa) begin
        _T_26_17 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h12 == io_wa) begin
        _T_26_18 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h13 == io_wa) begin
        _T_26_19 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h14 == io_wa) begin
        _T_26_20 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h15 == io_wa) begin
        _T_26_21 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h16 == io_wa) begin
        _T_26_22 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h17 == io_wa) begin
        _T_26_23 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h18 == io_wa) begin
        _T_26_24 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h19 == io_wa) begin
        _T_26_25 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1a == io_wa) begin
        _T_26_26 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1b == io_wa) begin
        _T_26_27 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1c == io_wa) begin
        _T_26_28 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1d == io_wa) begin
        _T_26_29 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1e == io_wa) begin
        _T_26_30 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1f == io_wa) begin
        _T_26_31 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h20 == io_wa) begin
        _T_26_32 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h21 == io_wa) begin
        _T_26_33 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h22 == io_wa) begin
        _T_26_34 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h23 == io_wa) begin
        _T_26_35 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h24 == io_wa) begin
        _T_26_36 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h25 == io_wa) begin
        _T_26_37 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h26 == io_wa) begin
        _T_26_38 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h27 == io_wa) begin
        _T_26_39 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h28 == io_wa) begin
        _T_26_40 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h29 == io_wa) begin
        _T_26_41 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2a == io_wa) begin
        _T_26_42 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2b == io_wa) begin
        _T_26_43 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2c == io_wa) begin
        _T_26_44 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2d == io_wa) begin
        _T_26_45 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2e == io_wa) begin
        _T_26_46 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2f == io_wa) begin
        _T_26_47 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h30 == io_wa) begin
        _T_26_48 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h31 == io_wa) begin
        _T_26_49 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h32 == io_wa) begin
        _T_26_50 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h33 == io_wa) begin
        _T_26_51 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h34 == io_wa) begin
        _T_26_52 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h35 == io_wa) begin
        _T_26_53 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h36 == io_wa) begin
        _T_26_54 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h37 == io_wa) begin
        _T_26_55 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h38 == io_wa) begin
        _T_26_56 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h39 == io_wa) begin
        _T_26_57 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3a == io_wa) begin
        _T_26_58 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3b == io_wa) begin
        _T_26_59 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3c == io_wa) begin
        _T_26_60 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3d == io_wa) begin
        _T_26_61 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3e == io_wa) begin
        _T_26_62 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3f == io_wa) begin
        _T_26_63 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h40 == io_wa) begin
        _T_26_64 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h41 == io_wa) begin
        _T_26_65 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h42 == io_wa) begin
        _T_26_66 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h43 == io_wa) begin
        _T_26_67 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h44 == io_wa) begin
        _T_26_68 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h45 == io_wa) begin
        _T_26_69 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h46 == io_wa) begin
        _T_26_70 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h47 == io_wa) begin
        _T_26_71 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h48 == io_wa) begin
        _T_26_72 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h49 == io_wa) begin
        _T_26_73 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4a == io_wa) begin
        _T_26_74 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4b == io_wa) begin
        _T_26_75 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4c == io_wa) begin
        _T_26_76 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4d == io_wa) begin
        _T_26_77 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4e == io_wa) begin
        _T_26_78 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4f == io_wa) begin
        _T_26_79 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h50 == io_wa) begin
        _T_26_80 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h51 == io_wa) begin
        _T_26_81 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h52 == io_wa) begin
        _T_26_82 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h53 == io_wa) begin
        _T_26_83 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h54 == io_wa) begin
        _T_26_84 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h55 == io_wa) begin
        _T_26_85 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h56 == io_wa) begin
        _T_26_86 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h57 == io_wa) begin
        _T_26_87 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h58 == io_wa) begin
        _T_26_88 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h59 == io_wa) begin
        _T_26_89 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5a == io_wa) begin
        _T_26_90 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5b == io_wa) begin
        _T_26_91 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5c == io_wa) begin
        _T_26_92 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5d == io_wa) begin
        _T_26_93 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5e == io_wa) begin
        _T_26_94 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5f == io_wa) begin
        _T_26_95 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h60 == io_wa) begin
        _T_26_96 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h61 == io_wa) begin
        _T_26_97 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h62 == io_wa) begin
        _T_26_98 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h63 == io_wa) begin
        _T_26_99 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h64 == io_wa) begin
        _T_26_100 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h65 == io_wa) begin
        _T_26_101 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h66 == io_wa) begin
        _T_26_102 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h67 == io_wa) begin
        _T_26_103 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h68 == io_wa) begin
        _T_26_104 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h69 == io_wa) begin
        _T_26_105 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6a == io_wa) begin
        _T_26_106 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6b == io_wa) begin
        _T_26_107 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6c == io_wa) begin
        _T_26_108 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6d == io_wa) begin
        _T_26_109 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6e == io_wa) begin
        _T_26_110 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6f == io_wa) begin
        _T_26_111 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h70 == io_wa) begin
        _T_26_112 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h71 == io_wa) begin
        _T_26_113 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h72 == io_wa) begin
        _T_26_114 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h73 == io_wa) begin
        _T_26_115 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h74 == io_wa) begin
        _T_26_116 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h75 == io_wa) begin
        _T_26_117 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h76 == io_wa) begin
        _T_26_118 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h77 == io_wa) begin
        _T_26_119 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h78 == io_wa) begin
        _T_26_120 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h79 == io_wa) begin
        _T_26_121 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7a == io_wa) begin
        _T_26_122 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7b == io_wa) begin
        _T_26_123 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7c == io_wa) begin
        _T_26_124 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7d == io_wa) begin
        _T_26_125 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7e == io_wa) begin
        _T_26_126 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7f == io_wa) begin
        _T_26_127 <= io_di;
      end
    end
    if (io_re) begin
      _T_158 <= io_ra;
    end
    if (io_ore) begin
      if (7'h7f == _T_158) begin
        _T_160 <= _T_26_127;
      end else begin
        if (7'h7e == _T_158) begin
          _T_160 <= _T_26_126;
        end else begin
          if (7'h7d == _T_158) begin
            _T_160 <= _T_26_125;
          end else begin
            if (7'h7c == _T_158) begin
              _T_160 <= _T_26_124;
            end else begin
              if (7'h7b == _T_158) begin
                _T_160 <= _T_26_123;
              end else begin
                if (7'h7a == _T_158) begin
                  _T_160 <= _T_26_122;
                end else begin
                  if (7'h79 == _T_158) begin
                    _T_160 <= _T_26_121;
                  end else begin
                    if (7'h78 == _T_158) begin
                      _T_160 <= _T_26_120;
                    end else begin
                      if (7'h77 == _T_158) begin
                        _T_160 <= _T_26_119;
                      end else begin
                        if (7'h76 == _T_158) begin
                          _T_160 <= _T_26_118;
                        end else begin
                          if (7'h75 == _T_158) begin
                            _T_160 <= _T_26_117;
                          end else begin
                            if (7'h74 == _T_158) begin
                              _T_160 <= _T_26_116;
                            end else begin
                              if (7'h73 == _T_158) begin
                                _T_160 <= _T_26_115;
                              end else begin
                                if (7'h72 == _T_158) begin
                                  _T_160 <= _T_26_114;
                                end else begin
                                  if (7'h71 == _T_158) begin
                                    _T_160 <= _T_26_113;
                                  end else begin
                                    if (7'h70 == _T_158) begin
                                      _T_160 <= _T_26_112;
                                    end else begin
                                      if (7'h6f == _T_158) begin
                                        _T_160 <= _T_26_111;
                                      end else begin
                                        if (7'h6e == _T_158) begin
                                          _T_160 <= _T_26_110;
                                        end else begin
                                          if (7'h6d == _T_158) begin
                                            _T_160 <= _T_26_109;
                                          end else begin
                                            if (7'h6c == _T_158) begin
                                              _T_160 <= _T_26_108;
                                            end else begin
                                              if (7'h6b == _T_158) begin
                                                _T_160 <= _T_26_107;
                                              end else begin
                                                if (7'h6a == _T_158) begin
                                                  _T_160 <= _T_26_106;
                                                end else begin
                                                  if (7'h69 == _T_158) begin
                                                    _T_160 <= _T_26_105;
                                                  end else begin
                                                    if (7'h68 == _T_158) begin
                                                      _T_160 <= _T_26_104;
                                                    end else begin
                                                      if (7'h67 == _T_158) begin
                                                        _T_160 <= _T_26_103;
                                                      end else begin
                                                        if (7'h66 == _T_158) begin
                                                          _T_160 <= _T_26_102;
                                                        end else begin
                                                          if (7'h65 == _T_158) begin
                                                            _T_160 <= _T_26_101;
                                                          end else begin
                                                            if (7'h64 == _T_158) begin
                                                              _T_160 <= _T_26_100;
                                                            end else begin
                                                              if (7'h63 == _T_158) begin
                                                                _T_160 <= _T_26_99;
                                                              end else begin
                                                                if (7'h62 == _T_158) begin
                                                                  _T_160 <= _T_26_98;
                                                                end else begin
                                                                  if (7'h61 == _T_158) begin
                                                                    _T_160 <= _T_26_97;
                                                                  end else begin
                                                                    if (7'h60 == _T_158) begin
                                                                      _T_160 <= _T_26_96;
                                                                    end else begin
                                                                      if (7'h5f == _T_158) begin
                                                                        _T_160 <= _T_26_95;
                                                                      end else begin
                                                                        if (7'h5e == _T_158) begin
                                                                          _T_160 <= _T_26_94;
                                                                        end else begin
                                                                          if (7'h5d == _T_158) begin
                                                                            _T_160 <= _T_26_93;
                                                                          end else begin
                                                                            if (7'h5c == _T_158) begin
                                                                              _T_160 <= _T_26_92;
                                                                            end else begin
                                                                              if (7'h5b == _T_158) begin
                                                                                _T_160 <= _T_26_91;
                                                                              end else begin
                                                                                if (7'h5a == _T_158) begin
                                                                                  _T_160 <= _T_26_90;
                                                                                end else begin
                                                                                  if (7'h59 == _T_158) begin
                                                                                    _T_160 <= _T_26_89;
                                                                                  end else begin
                                                                                    if (7'h58 == _T_158) begin
                                                                                      _T_160 <= _T_26_88;
                                                                                    end else begin
                                                                                      if (7'h57 == _T_158) begin
                                                                                        _T_160 <= _T_26_87;
                                                                                      end else begin
                                                                                        if (7'h56 == _T_158) begin
                                                                                          _T_160 <= _T_26_86;
                                                                                        end else begin
                                                                                          if (7'h55 == _T_158) begin
                                                                                            _T_160 <= _T_26_85;
                                                                                          end else begin
                                                                                            if (7'h54 == _T_158) begin
                                                                                              _T_160 <= _T_26_84;
                                                                                            end else begin
                                                                                              if (7'h53 == _T_158) begin
                                                                                                _T_160 <= _T_26_83;
                                                                                              end else begin
                                                                                                if (7'h52 == _T_158) begin
                                                                                                  _T_160 <= _T_26_82;
                                                                                                end else begin
                                                                                                  if (7'h51 == _T_158) begin
                                                                                                    _T_160 <= _T_26_81;
                                                                                                  end else begin
                                                                                                    if (7'h50 == _T_158) begin
                                                                                                      _T_160 <= _T_26_80;
                                                                                                    end else begin
                                                                                                      if (7'h4f == _T_158) begin
                                                                                                        _T_160 <= _T_26_79;
                                                                                                      end else begin
                                                                                                        if (7'h4e == _T_158) begin
                                                                                                          _T_160 <= _T_26_78;
                                                                                                        end else begin
                                                                                                          if (7'h4d == _T_158) begin
                                                                                                            _T_160 <= _T_26_77;
                                                                                                          end else begin
                                                                                                            if (7'h4c == _T_158) begin
                                                                                                              _T_160 <= _T_26_76;
                                                                                                            end else begin
                                                                                                              if (7'h4b == _T_158) begin
                                                                                                                _T_160 <= _T_26_75;
                                                                                                              end else begin
                                                                                                                if (7'h4a == _T_158) begin
                                                                                                                  _T_160 <= _T_26_74;
                                                                                                                end else begin
                                                                                                                  if (7'h49 == _T_158) begin
                                                                                                                    _T_160 <= _T_26_73;
                                                                                                                  end else begin
                                                                                                                    if (7'h48 == _T_158) begin
                                                                                                                      _T_160 <= _T_26_72;
                                                                                                                    end else begin
                                                                                                                      if (7'h47 == _T_158) begin
                                                                                                                        _T_160 <= _T_26_71;
                                                                                                                      end else begin
                                                                                                                        if (7'h46 == _T_158) begin
                                                                                                                          _T_160 <= _T_26_70;
                                                                                                                        end else begin
                                                                                                                          if (7'h45 == _T_158) begin
                                                                                                                            _T_160 <= _T_26_69;
                                                                                                                          end else begin
                                                                                                                            if (7'h44 == _T_158) begin
                                                                                                                              _T_160 <= _T_26_68;
                                                                                                                            end else begin
                                                                                                                              if (7'h43 == _T_158) begin
                                                                                                                                _T_160 <= _T_26_67;
                                                                                                                              end else begin
                                                                                                                                if (7'h42 == _T_158) begin
                                                                                                                                  _T_160 <= _T_26_66;
                                                                                                                                end else begin
                                                                                                                                  if (7'h41 == _T_158) begin
                                                                                                                                    _T_160 <= _T_26_65;
                                                                                                                                  end else begin
                                                                                                                                    if (7'h40 == _T_158) begin
                                                                                                                                      _T_160 <= _T_26_64;
                                                                                                                                    end else begin
                                                                                                                                      if (7'h3f == _T_158) begin
                                                                                                                                        _T_160 <= _T_26_63;
                                                                                                                                      end else begin
                                                                                                                                        if (7'h3e == _T_158) begin
                                                                                                                                          _T_160 <= _T_26_62;
                                                                                                                                        end else begin
                                                                                                                                          if (7'h3d == _T_158) begin
                                                                                                                                            _T_160 <= _T_26_61;
                                                                                                                                          end else begin
                                                                                                                                            if (7'h3c == _T_158) begin
                                                                                                                                              _T_160 <= _T_26_60;
                                                                                                                                            end else begin
                                                                                                                                              if (7'h3b == _T_158) begin
                                                                                                                                                _T_160 <= _T_26_59;
                                                                                                                                              end else begin
                                                                                                                                                if (7'h3a == _T_158) begin
                                                                                                                                                  _T_160 <= _T_26_58;
                                                                                                                                                end else begin
                                                                                                                                                  if (7'h39 == _T_158) begin
                                                                                                                                                    _T_160 <= _T_26_57;
                                                                                                                                                  end else begin
                                                                                                                                                    if (7'h38 == _T_158) begin
                                                                                                                                                      _T_160 <= _T_26_56;
                                                                                                                                                    end else begin
                                                                                                                                                      if (7'h37 == _T_158) begin
                                                                                                                                                        _T_160 <= _T_26_55;
                                                                                                                                                      end else begin
                                                                                                                                                        if (7'h36 == _T_158) begin
                                                                                                                                                          _T_160 <= _T_26_54;
                                                                                                                                                        end else begin
                                                                                                                                                          if (7'h35 == _T_158) begin
                                                                                                                                                            _T_160 <= _T_26_53;
                                                                                                                                                          end else begin
                                                                                                                                                            if (7'h34 == _T_158) begin
                                                                                                                                                              _T_160 <= _T_26_52;
                                                                                                                                                            end else begin
                                                                                                                                                              if (7'h33 == _T_158) begin
                                                                                                                                                                _T_160 <= _T_26_51;
                                                                                                                                                              end else begin
                                                                                                                                                                if (7'h32 == _T_158) begin
                                                                                                                                                                  _T_160 <= _T_26_50;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (7'h31 == _T_158) begin
                                                                                                                                                                    _T_160 <= _T_26_49;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (7'h30 == _T_158) begin
                                                                                                                                                                      _T_160 <= _T_26_48;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (7'h2f == _T_158) begin
                                                                                                                                                                        _T_160 <= _T_26_47;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (7'h2e == _T_158) begin
                                                                                                                                                                          _T_160 <= _T_26_46;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (7'h2d == _T_158) begin
                                                                                                                                                                            _T_160 <= _T_26_45;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (7'h2c == _T_158) begin
                                                                                                                                                                              _T_160 <= _T_26_44;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (7'h2b == _T_158) begin
                                                                                                                                                                                _T_160 <= _T_26_43;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (7'h2a == _T_158) begin
                                                                                                                                                                                  _T_160 <= _T_26_42;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (7'h29 == _T_158) begin
                                                                                                                                                                                    _T_160 <= _T_26_41;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (7'h28 == _T_158) begin
                                                                                                                                                                                      _T_160 <= _T_26_40;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (7'h27 == _T_158) begin
                                                                                                                                                                                        _T_160 <= _T_26_39;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (7'h26 == _T_158) begin
                                                                                                                                                                                          _T_160 <= _T_26_38;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (7'h25 == _T_158) begin
                                                                                                                                                                                            _T_160 <= _T_26_37;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (7'h24 == _T_158) begin
                                                                                                                                                                                              _T_160 <= _T_26_36;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (7'h23 == _T_158) begin
                                                                                                                                                                                                _T_160 <= _T_26_35;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (7'h22 == _T_158) begin
                                                                                                                                                                                                  _T_160 <= _T_26_34;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (7'h21 == _T_158) begin
                                                                                                                                                                                                    _T_160 <= _T_26_33;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (7'h20 == _T_158) begin
                                                                                                                                                                                                      _T_160 <= _T_26_32;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (7'h1f == _T_158) begin
                                                                                                                                                                                                        _T_160 <= _T_26_31;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (7'h1e == _T_158) begin
                                                                                                                                                                                                          _T_160 <= _T_26_30;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (7'h1d == _T_158) begin
                                                                                                                                                                                                            _T_160 <= _T_26_29;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (7'h1c == _T_158) begin
                                                                                                                                                                                                              _T_160 <= _T_26_28;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (7'h1b == _T_158) begin
                                                                                                                                                                                                                _T_160 <= _T_26_27;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (7'h1a == _T_158) begin
                                                                                                                                                                                                                  _T_160 <= _T_26_26;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (7'h19 == _T_158) begin
                                                                                                                                                                                                                    _T_160 <= _T_26_25;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (7'h18 == _T_158) begin
                                                                                                                                                                                                                      _T_160 <= _T_26_24;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (7'h17 == _T_158) begin
                                                                                                                                                                                                                        _T_160 <= _T_26_23;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (7'h16 == _T_158) begin
                                                                                                                                                                                                                          _T_160 <= _T_26_22;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (7'h15 == _T_158) begin
                                                                                                                                                                                                                            _T_160 <= _T_26_21;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (7'h14 == _T_158) begin
                                                                                                                                                                                                                              _T_160 <= _T_26_20;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (7'h13 == _T_158) begin
                                                                                                                                                                                                                                _T_160 <= _T_26_19;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (7'h12 == _T_158) begin
                                                                                                                                                                                                                                  _T_160 <= _T_26_18;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (7'h11 == _T_158) begin
                                                                                                                                                                                                                                    _T_160 <= _T_26_17;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (7'h10 == _T_158) begin
                                                                                                                                                                                                                                      _T_160 <= _T_26_16;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (7'hf == _T_158) begin
                                                                                                                                                                                                                                        _T_160 <= _T_26_15;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (7'he == _T_158) begin
                                                                                                                                                                                                                                          _T_160 <= _T_26_14;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (7'hd == _T_158) begin
                                                                                                                                                                                                                                            _T_160 <= _T_26_13;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (7'hc == _T_158) begin
                                                                                                                                                                                                                                              _T_160 <= _T_26_12;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (7'hb == _T_158) begin
                                                                                                                                                                                                                                                _T_160 <= _T_26_11;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (7'ha == _T_158) begin
                                                                                                                                                                                                                                                  _T_160 <= _T_26_10;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (7'h9 == _T_158) begin
                                                                                                                                                                                                                                                    _T_160 <= _T_26_9;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (7'h8 == _T_158) begin
                                                                                                                                                                                                                                                      _T_160 <= _T_26_8;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (7'h7 == _T_158) begin
                                                                                                                                                                                                                                                        _T_160 <= _T_26_7;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (7'h6 == _T_158) begin
                                                                                                                                                                                                                                                          _T_160 <= _T_26_6;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (7'h5 == _T_158) begin
                                                                                                                                                                                                                                                            _T_160 <= _T_26_5;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (7'h4 == _T_158) begin
                                                                                                                                                                                                                                                              _T_160 <= _T_26_4;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (7'h3 == _T_158) begin
                                                                                                                                                                                                                                                                _T_160 <= _T_26_3;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (7'h2 == _T_158) begin
                                                                                                                                                                                                                                                                  _T_160 <= _T_26_2;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  if (7'h1 == _T_158) begin
                                                                                                                                                                                                                                                                    _T_160 <= _T_26_1;
                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                    _T_160 <= _T_26_0;
                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_fifo_3( // @[:@6045.2]
  input         clock, // @[:@6046.4]
  input         reset, // @[:@6047.4]
  input         io_clk, // @[:@6048.4]
  input         io_wr_pvld, // @[:@6048.4]
  output        io_wr_prdy, // @[:@6048.4]
  input  [10:0] io_wr_pd, // @[:@6048.4]
  output        io_rd_pvld, // @[:@6048.4]
  input         io_rd_prdy, // @[:@6048.4]
  output [10:0] io_rd_pd // @[:@6048.4]
);
  wire  nv_ram_rwsp_io_clk; // @[FIFO.scala 270:29:@6122.4]
  wire  nv_ram_rwsp_io_re; // @[FIFO.scala 270:29:@6122.4]
  wire  nv_ram_rwsp_io_we; // @[FIFO.scala 270:29:@6122.4]
  wire  nv_ram_rwsp_io_ore; // @[FIFO.scala 270:29:@6122.4]
  wire [6:0] nv_ram_rwsp_io_ra; // @[FIFO.scala 270:29:@6122.4]
  wire [6:0] nv_ram_rwsp_io_wa; // @[FIFO.scala 270:29:@6122.4]
  wire [10:0] nv_ram_rwsp_io_di; // @[FIFO.scala 270:29:@6122.4]
  wire [10:0] nv_ram_rwsp_io_dout; // @[FIFO.scala 270:29:@6122.4]
  reg  _T_26; // @[FIFO.scala 156:56:@6057.4]
  reg [31:0] _RAND_0;
  reg  _T_29; // @[FIFO.scala 158:52:@6058.4]
  reg [31:0] _RAND_1;
  reg [10:0] _T_31; // @[FIFO.scala 159:64:@6059.4]
  reg [31:0] _RAND_2;
  reg  _T_34; // @[FIFO.scala 160:52:@6060.4]
  reg [31:0] _RAND_3;
  wire  _T_125; // @[FIFO.scala 331:38:@6153.4]
  wire  _T_54; // @[FIFO.scala 183:39:@6081.4]
  wire  _T_55; // @[FIFO.scala 183:36:@6082.4]
  reg [7:0] _T_60; // @[FIFO.scala 186:53:@6085.4]
  reg [31:0] _RAND_4;
  wire [8:0] _T_67; // @[FIFO.scala 191:69:@6090.4]
  wire [7:0] _T_68; // @[FIFO.scala 191:69:@6091.4]
  wire [7:0] _T_69; // @[FIFO.scala 191:46:@6092.4]
  wire  _T_72; // @[FIFO.scala 194:80:@6094.4]
  wire  _T_74; // @[FIFO.scala 195:40:@6095.4]
  wire [8:0] _T_62; // @[FIFO.scala 190:76:@6086.4]
  wire [8:0] _T_63; // @[FIFO.scala 190:76:@6087.4]
  wire [7:0] _T_64; // @[FIFO.scala 190:76:@6088.4]
  wire [7:0] _T_65; // @[FIFO.scala 190:43:@6089.4]
  wire [7:0] _T_70; // @[FIFO.scala 192:32:@6093.4]
  wire  _T_37; // @[FIFO.scala 166:60:@6062.4]
  wire  _T_39; // @[FIFO.scala 166:80:@6063.4]
  wire  _T_40; // @[FIFO.scala 166:77:@6064.4]
  wire  _T_41; // @[FIFO.scala 167:38:@6065.4]
  wire  _T_42; // @[FIFO.scala 168:45:@6066.4]
  wire  _T_44; // @[FIFO.scala 171:18:@6068.4]
  wire  _T_46; // @[FIFO.scala 172:45:@6070.6]
  wire  _T_47; // @[FIFO.scala 172:42:@6071.6]
  wire  _GEN_0; // @[FIFO.scala 171:34:@6069.4]
  wire  _T_50; // @[FIFO.scala 176:34:@6075.4]
  wire  _T_82; // @[FIFO.scala 202:27:@6103.4]
  wire [7:0] _GEN_2; // @[FIFO.scala 202:40:@6104.4]
  reg [6:0] _T_85; // @[FIFO.scala 215:68:@6107.4]
  reg [31:0] _RAND_5;
  wire [7:0] _T_87; // @[FIFO.scala 217:42:@6108.4]
  wire [6:0] _T_88; // @[FIFO.scala 217:42:@6109.4]
  wire [6:0] _GEN_3; // @[FIFO.scala 218:29:@6110.4]
  reg [6:0] _T_93; // @[FIFO.scala 224:63:@6114.4]
  reg [31:0] _RAND_6;
  wire [7:0] _T_95; // @[FIFO.scala 225:42:@6115.4]
  wire [6:0] _T_96; // @[FIFO.scala 225:42:@6116.4]
  wire [6:0] _GEN_4; // @[FIFO.scala 227:29:@6117.4]
  reg  _T_104; // @[FIFO.scala 289:73:@6136.4]
  reg [31:0] _RAND_7;
  reg  _T_107; // @[FIFO.scala 295:72:@6138.4]
  reg [31:0] _RAND_8;
  reg  _T_110; // @[FIFO.scala 297:97:@6139.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_113; // @[FIFO.scala 299:53:@6140.4]
  reg [31:0] _RAND_10;
  wire [8:0] _T_115; // @[FIFO.scala 300:74:@6141.4]
  wire [8:0] _T_116; // @[FIFO.scala 300:74:@6142.4]
  wire [7:0] _T_117; // @[FIFO.scala 300:74:@6143.4]
  wire [7:0] _T_118; // @[FIFO.scala 300:43:@6144.4]
  wire [8:0] _T_120; // @[FIFO.scala 301:68:@6145.4]
  wire [7:0] _T_121; // @[FIFO.scala 301:68:@6146.4]
  wire [7:0] _T_122; // @[FIFO.scala 301:46:@6147.4]
  wire [7:0] _T_123; // @[FIFO.scala 302:32:@6148.4]
  wire  _T_124; // @[FIFO.scala 303:25:@6149.4]
  wire [7:0] _GEN_5; // @[FIFO.scala 303:39:@6150.4]
  wire  _T_127; // @[FIFO.scala 333:77:@6155.4]
  wire  _T_129; // @[FIFO.scala 334:83:@6156.4]
  wire  _T_130; // @[FIFO.scala 335:44:@6157.4]
  wire  _T_131; // @[FIFO.scala 336:60:@6158.4]
  wire  _T_133; // @[FIFO.scala 336:81:@6160.4]
  wire  _GEN_6; // @[FIFO.scala 338:43:@6164.4]
  wire  _T_137; // @[FIFO.scala 341:66:@6167.4]
  wire  _T_138; // @[FIFO.scala 341:63:@6168.4]
  wire  _T_139; // @[FIFO.scala 341:43:@6169.4]
  nv_ram_rwsp_3 nv_ram_rwsp ( // @[FIFO.scala 270:29:@6122.4]
    .io_clk(nv_ram_rwsp_io_clk),
    .io_re(nv_ram_rwsp_io_re),
    .io_we(nv_ram_rwsp_io_we),
    .io_ore(nv_ram_rwsp_io_ore),
    .io_ra(nv_ram_rwsp_io_ra),
    .io_wa(nv_ram_rwsp_io_wa),
    .io_di(nv_ram_rwsp_io_di),
    .io_dout(nv_ram_rwsp_io_dout)
  );
  assign _T_125 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 331:38:@6153.4]
  assign _T_54 = _T_26 == 1'h0; // @[FIFO.scala 183:39:@6081.4]
  assign _T_55 = _T_29 & _T_54; // @[FIFO.scala 183:36:@6082.4]
  assign _T_67 = _T_60 + 8'h1; // @[FIFO.scala 191:69:@6090.4]
  assign _T_68 = _T_60 + 8'h1; // @[FIFO.scala 191:69:@6091.4]
  assign _T_69 = _T_55 ? _T_68 : _T_60; // @[FIFO.scala 191:46:@6092.4]
  assign _T_72 = _T_69 == 8'h80; // @[FIFO.scala 194:80:@6094.4]
  assign _T_74 = _T_125 ? 1'h0 : _T_72; // @[FIFO.scala 195:40:@6095.4]
  assign _T_62 = _T_60 - 8'h1; // @[FIFO.scala 190:76:@6086.4]
  assign _T_63 = $unsigned(_T_62); // @[FIFO.scala 190:76:@6087.4]
  assign _T_64 = _T_63[7:0]; // @[FIFO.scala 190:76:@6088.4]
  assign _T_65 = _T_55 ? _T_60 : _T_64; // @[FIFO.scala 190:43:@6089.4]
  assign _T_70 = _T_125 ? _T_65 : _T_69; // @[FIFO.scala 192:32:@6093.4]
  assign _T_37 = _T_29 & _T_74; // @[FIFO.scala 166:60:@6062.4]
  assign _T_39 = _T_55 == 1'h0; // @[FIFO.scala 166:80:@6063.4]
  assign _T_40 = _T_37 & _T_39; // @[FIFO.scala 166:77:@6064.4]
  assign _T_41 = io_wr_pvld ? _T_74 : _T_40; // @[FIFO.scala 167:38:@6065.4]
  assign _T_42 = _T_29 & _T_26; // @[FIFO.scala 168:45:@6066.4]
  assign _T_44 = _T_42 == 1'h0; // @[FIFO.scala 171:18:@6068.4]
  assign _T_46 = _T_34 == 1'h0; // @[FIFO.scala 172:45:@6070.6]
  assign _T_47 = io_wr_pvld & _T_46; // @[FIFO.scala 172:42:@6071.6]
  assign _GEN_0 = _T_44 ? _T_47 : _T_29; // @[FIFO.scala 171:34:@6069.4]
  assign _T_50 = _T_46 & io_wr_pvld; // @[FIFO.scala 176:34:@6075.4]
  assign _T_82 = _T_55 ^ _T_125; // @[FIFO.scala 202:27:@6103.4]
  assign _GEN_2 = _T_82 ? _T_70 : _T_60; // @[FIFO.scala 202:40:@6104.4]
  assign _T_87 = _T_85 + 7'h1; // @[FIFO.scala 217:42:@6108.4]
  assign _T_88 = _T_85 + 7'h1; // @[FIFO.scala 217:42:@6109.4]
  assign _GEN_3 = _T_55 ? _T_88 : _T_85; // @[FIFO.scala 218:29:@6110.4]
  assign _T_95 = _T_93 + 7'h1; // @[FIFO.scala 225:42:@6115.4]
  assign _T_96 = _T_93 + 7'h1; // @[FIFO.scala 225:42:@6116.4]
  assign _GEN_4 = _T_125 ? _T_96 : _T_93; // @[FIFO.scala 227:29:@6117.4]
  assign _T_115 = _T_113 - 8'h1; // @[FIFO.scala 300:74:@6141.4]
  assign _T_116 = $unsigned(_T_115); // @[FIFO.scala 300:74:@6142.4]
  assign _T_117 = _T_116[7:0]; // @[FIFO.scala 300:74:@6143.4]
  assign _T_118 = _T_104 ? _T_113 : _T_117; // @[FIFO.scala 300:43:@6144.4]
  assign _T_120 = _T_113 + 8'h1; // @[FIFO.scala 301:68:@6145.4]
  assign _T_121 = _T_113 + 8'h1; // @[FIFO.scala 301:68:@6146.4]
  assign _T_122 = _T_104 ? _T_121 : _T_113; // @[FIFO.scala 301:46:@6147.4]
  assign _T_123 = _T_125 ? _T_118 : _T_122; // @[FIFO.scala 302:32:@6148.4]
  assign _T_124 = _T_104 | _T_125; // @[FIFO.scala 303:25:@6149.4]
  assign _GEN_5 = _T_124 ? _T_123 : _T_113; // @[FIFO.scala 303:39:@6150.4]
  assign _T_127 = _T_118 != 8'h0; // @[FIFO.scala 333:77:@6155.4]
  assign _T_129 = _T_122 != 8'h0; // @[FIFO.scala 334:83:@6156.4]
  assign _T_130 = _T_125 ? _T_127 : _T_129; // @[FIFO.scala 335:44:@6157.4]
  assign _T_131 = ~ _T_107; // @[FIFO.scala 336:60:@6158.4]
  assign _T_133 = _T_131 | _T_125; // @[FIFO.scala 336:81:@6160.4]
  assign _GEN_6 = _T_124 ? _T_130 : _T_107; // @[FIFO.scala 338:43:@6164.4]
  assign _T_137 = io_rd_prdy == 1'h0; // @[FIFO.scala 341:66:@6167.4]
  assign _T_138 = _T_110 & _T_137; // @[FIFO.scala 341:63:@6168.4]
  assign _T_139 = _T_107 | _T_138; // @[FIFO.scala 341:43:@6169.4]
  assign io_wr_prdy = _T_34 == 1'h0; // @[FIFO.scala 182:20:@6080.4]
  assign io_rd_pvld = _T_110; // @[FIFO.scala 344:24:@6171.4]
  assign io_rd_pd = nv_ram_rwsp_io_dout; // @[FIFO.scala 345:22:@6172.4]
  assign nv_ram_rwsp_io_clk = io_clk; // @[FIFO.scala 271:24:@6125.4]
  assign nv_ram_rwsp_io_re = _T_130 & _T_133; // @[FIFO.scala 279:23:@6132.4]
  assign nv_ram_rwsp_io_we = _T_29 & _T_54; // @[FIFO.scala 276:23:@6128.4]
  assign nv_ram_rwsp_io_ore = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 280:24:@6133.4]
  assign nv_ram_rwsp_io_ra = _T_125 ? _T_96 : _T_93; // @[FIFO.scala 278:23:@6131.4]
  assign nv_ram_rwsp_io_wa = _T_85; // @[FIFO.scala 274:27:@6127.4]
  assign nv_ram_rwsp_io_di = _T_31; // @[FIFO.scala 277:23:@6129.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_26 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_31 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_34 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_60 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_85 = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_93 = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_104 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_107 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_110 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_113 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_125) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_72;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_29 <= _T_47;
      end
    end
    if (_T_50) begin
      _T_31 <= io_wr_pd;
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (io_wr_pvld) begin
        if (_T_125) begin
          _T_34 <= 1'h0;
        end else begin
          _T_34 <= _T_72;
        end
      end else begin
        _T_34 <= _T_40;
      end
    end
    if (reset) begin
      _T_60 <= 8'h0;
    end else begin
      if (_T_82) begin
        if (_T_125) begin
          if (!(_T_55)) begin
            _T_60 <= _T_64;
          end
        end else begin
          if (_T_55) begin
            _T_60 <= _T_68;
          end
        end
      end
    end
    if (reset) begin
      _T_85 <= 7'h0;
    end else begin
      if (_T_55) begin
        _T_85 <= _T_88;
      end
    end
    if (reset) begin
      _T_93 <= 7'h0;
    end else begin
      if (_T_125) begin
        _T_93 <= _T_96;
      end
    end
    if (reset) begin
      _T_104 <= 1'h0;
    end else begin
      _T_104 <= _T_55;
    end
    if (reset) begin
      _T_107 <= 1'h0;
    end else begin
      if (_T_124) begin
        if (_T_125) begin
          _T_107 <= _T_127;
        end else begin
          _T_107 <= _T_129;
        end
      end
    end
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      _T_110 <= _T_139;
    end
    if (reset) begin
      _T_113 <= 8'h0;
    end else begin
      if (_T_124) begin
        if (_T_125) begin
          if (!(_T_104)) begin
            _T_113 <= _T_117;
          end
        end else begin
          if (_T_104) begin
            _T_113 <= _T_121;
          end
        end
      end
    end
  end
endmodule
module nv_flopram( // @[:@6219.2]
  input  [10:0] io_di, // @[:@6222.4]
  input  [7:0]  io_ra, // @[:@6222.4]
  output [10:0] io_dout // @[:@6222.4]
);
  wire  _T_669; // @[Mux.scala 46:19:@6874.4]
  wire [10:0] _T_670; // @[Mux.scala 46:16:@6875.4]
  wire  _T_671; // @[Mux.scala 46:19:@6876.4]
  wire [10:0] _T_672; // @[Mux.scala 46:16:@6877.4]
  wire  _T_673; // @[Mux.scala 46:19:@6878.4]
  wire [10:0] _T_674; // @[Mux.scala 46:16:@6879.4]
  wire  _T_675; // @[Mux.scala 46:19:@6880.4]
  wire [10:0] _T_676; // @[Mux.scala 46:16:@6881.4]
  wire  _T_677; // @[Mux.scala 46:19:@6882.4]
  wire [10:0] _T_678; // @[Mux.scala 46:16:@6883.4]
  wire  _T_679; // @[Mux.scala 46:19:@6884.4]
  wire [10:0] _T_680; // @[Mux.scala 46:16:@6885.4]
  wire  _T_681; // @[Mux.scala 46:19:@6886.4]
  wire [10:0] _T_682; // @[Mux.scala 46:16:@6887.4]
  wire  _T_683; // @[Mux.scala 46:19:@6888.4]
  wire [10:0] _T_684; // @[Mux.scala 46:16:@6889.4]
  wire  _T_685; // @[Mux.scala 46:19:@6890.4]
  wire [10:0] _T_686; // @[Mux.scala 46:16:@6891.4]
  wire  _T_687; // @[Mux.scala 46:19:@6892.4]
  wire [10:0] _T_688; // @[Mux.scala 46:16:@6893.4]
  wire  _T_689; // @[Mux.scala 46:19:@6894.4]
  wire [10:0] _T_690; // @[Mux.scala 46:16:@6895.4]
  wire  _T_691; // @[Mux.scala 46:19:@6896.4]
  wire [10:0] _T_692; // @[Mux.scala 46:16:@6897.4]
  wire  _T_693; // @[Mux.scala 46:19:@6898.4]
  wire [10:0] _T_694; // @[Mux.scala 46:16:@6899.4]
  wire  _T_695; // @[Mux.scala 46:19:@6900.4]
  wire [10:0] _T_696; // @[Mux.scala 46:16:@6901.4]
  wire  _T_697; // @[Mux.scala 46:19:@6902.4]
  wire [10:0] _T_698; // @[Mux.scala 46:16:@6903.4]
  wire  _T_699; // @[Mux.scala 46:19:@6904.4]
  wire [10:0] _T_700; // @[Mux.scala 46:16:@6905.4]
  wire  _T_701; // @[Mux.scala 46:19:@6906.4]
  wire [10:0] _T_702; // @[Mux.scala 46:16:@6907.4]
  wire  _T_703; // @[Mux.scala 46:19:@6908.4]
  wire [10:0] _T_704; // @[Mux.scala 46:16:@6909.4]
  wire  _T_705; // @[Mux.scala 46:19:@6910.4]
  wire [10:0] _T_706; // @[Mux.scala 46:16:@6911.4]
  wire  _T_707; // @[Mux.scala 46:19:@6912.4]
  wire [10:0] _T_708; // @[Mux.scala 46:16:@6913.4]
  wire  _T_709; // @[Mux.scala 46:19:@6914.4]
  wire [10:0] _T_710; // @[Mux.scala 46:16:@6915.4]
  wire  _T_711; // @[Mux.scala 46:19:@6916.4]
  wire [10:0] _T_712; // @[Mux.scala 46:16:@6917.4]
  wire  _T_713; // @[Mux.scala 46:19:@6918.4]
  wire [10:0] _T_714; // @[Mux.scala 46:16:@6919.4]
  wire  _T_715; // @[Mux.scala 46:19:@6920.4]
  wire [10:0] _T_716; // @[Mux.scala 46:16:@6921.4]
  wire  _T_717; // @[Mux.scala 46:19:@6922.4]
  wire [10:0] _T_718; // @[Mux.scala 46:16:@6923.4]
  wire  _T_719; // @[Mux.scala 46:19:@6924.4]
  wire [10:0] _T_720; // @[Mux.scala 46:16:@6925.4]
  wire  _T_721; // @[Mux.scala 46:19:@6926.4]
  wire [10:0] _T_722; // @[Mux.scala 46:16:@6927.4]
  wire  _T_723; // @[Mux.scala 46:19:@6928.4]
  wire [10:0] _T_724; // @[Mux.scala 46:16:@6929.4]
  wire  _T_725; // @[Mux.scala 46:19:@6930.4]
  wire [10:0] _T_726; // @[Mux.scala 46:16:@6931.4]
  wire  _T_727; // @[Mux.scala 46:19:@6932.4]
  wire [10:0] _T_728; // @[Mux.scala 46:16:@6933.4]
  wire  _T_729; // @[Mux.scala 46:19:@6934.4]
  wire [10:0] _T_730; // @[Mux.scala 46:16:@6935.4]
  wire  _T_731; // @[Mux.scala 46:19:@6936.4]
  wire [10:0] _T_732; // @[Mux.scala 46:16:@6937.4]
  wire  _T_733; // @[Mux.scala 46:19:@6938.4]
  wire [10:0] _T_734; // @[Mux.scala 46:16:@6939.4]
  wire  _T_735; // @[Mux.scala 46:19:@6940.4]
  wire [10:0] _T_736; // @[Mux.scala 46:16:@6941.4]
  wire  _T_737; // @[Mux.scala 46:19:@6942.4]
  wire [10:0] _T_738; // @[Mux.scala 46:16:@6943.4]
  wire  _T_739; // @[Mux.scala 46:19:@6944.4]
  wire [10:0] _T_740; // @[Mux.scala 46:16:@6945.4]
  wire  _T_741; // @[Mux.scala 46:19:@6946.4]
  wire [10:0] _T_742; // @[Mux.scala 46:16:@6947.4]
  wire  _T_743; // @[Mux.scala 46:19:@6948.4]
  wire [10:0] _T_744; // @[Mux.scala 46:16:@6949.4]
  wire  _T_745; // @[Mux.scala 46:19:@6950.4]
  wire [10:0] _T_746; // @[Mux.scala 46:16:@6951.4]
  wire  _T_747; // @[Mux.scala 46:19:@6952.4]
  wire [10:0] _T_748; // @[Mux.scala 46:16:@6953.4]
  wire  _T_749; // @[Mux.scala 46:19:@6954.4]
  wire [10:0] _T_750; // @[Mux.scala 46:16:@6955.4]
  wire  _T_751; // @[Mux.scala 46:19:@6956.4]
  wire [10:0] _T_752; // @[Mux.scala 46:16:@6957.4]
  wire  _T_753; // @[Mux.scala 46:19:@6958.4]
  wire [10:0] _T_754; // @[Mux.scala 46:16:@6959.4]
  wire  _T_755; // @[Mux.scala 46:19:@6960.4]
  wire [10:0] _T_756; // @[Mux.scala 46:16:@6961.4]
  wire  _T_757; // @[Mux.scala 46:19:@6962.4]
  wire [10:0] _T_758; // @[Mux.scala 46:16:@6963.4]
  wire  _T_759; // @[Mux.scala 46:19:@6964.4]
  wire [10:0] _T_760; // @[Mux.scala 46:16:@6965.4]
  wire  _T_761; // @[Mux.scala 46:19:@6966.4]
  wire [10:0] _T_762; // @[Mux.scala 46:16:@6967.4]
  wire  _T_763; // @[Mux.scala 46:19:@6968.4]
  wire [10:0] _T_764; // @[Mux.scala 46:16:@6969.4]
  wire  _T_765; // @[Mux.scala 46:19:@6970.4]
  wire [10:0] _T_766; // @[Mux.scala 46:16:@6971.4]
  wire  _T_767; // @[Mux.scala 46:19:@6972.4]
  wire [10:0] _T_768; // @[Mux.scala 46:16:@6973.4]
  wire  _T_769; // @[Mux.scala 46:19:@6974.4]
  wire [10:0] _T_770; // @[Mux.scala 46:16:@6975.4]
  wire  _T_771; // @[Mux.scala 46:19:@6976.4]
  wire [10:0] _T_772; // @[Mux.scala 46:16:@6977.4]
  wire  _T_773; // @[Mux.scala 46:19:@6978.4]
  wire [10:0] _T_774; // @[Mux.scala 46:16:@6979.4]
  wire  _T_775; // @[Mux.scala 46:19:@6980.4]
  wire [10:0] _T_776; // @[Mux.scala 46:16:@6981.4]
  wire  _T_777; // @[Mux.scala 46:19:@6982.4]
  wire [10:0] _T_778; // @[Mux.scala 46:16:@6983.4]
  wire  _T_779; // @[Mux.scala 46:19:@6984.4]
  wire [10:0] _T_780; // @[Mux.scala 46:16:@6985.4]
  wire  _T_781; // @[Mux.scala 46:19:@6986.4]
  wire [10:0] _T_782; // @[Mux.scala 46:16:@6987.4]
  wire  _T_783; // @[Mux.scala 46:19:@6988.4]
  wire [10:0] _T_784; // @[Mux.scala 46:16:@6989.4]
  wire  _T_785; // @[Mux.scala 46:19:@6990.4]
  wire [10:0] _T_786; // @[Mux.scala 46:16:@6991.4]
  wire  _T_787; // @[Mux.scala 46:19:@6992.4]
  wire [10:0] _T_788; // @[Mux.scala 46:16:@6993.4]
  wire  _T_789; // @[Mux.scala 46:19:@6994.4]
  wire [10:0] _T_790; // @[Mux.scala 46:16:@6995.4]
  wire  _T_791; // @[Mux.scala 46:19:@6996.4]
  wire [10:0] _T_792; // @[Mux.scala 46:16:@6997.4]
  wire  _T_793; // @[Mux.scala 46:19:@6998.4]
  wire [10:0] _T_794; // @[Mux.scala 46:16:@6999.4]
  wire  _T_795; // @[Mux.scala 46:19:@7000.4]
  wire [10:0] _T_796; // @[Mux.scala 46:16:@7001.4]
  wire  _T_797; // @[Mux.scala 46:19:@7002.4]
  wire [10:0] _T_798; // @[Mux.scala 46:16:@7003.4]
  wire  _T_799; // @[Mux.scala 46:19:@7004.4]
  wire [10:0] _T_800; // @[Mux.scala 46:16:@7005.4]
  wire  _T_801; // @[Mux.scala 46:19:@7006.4]
  wire [10:0] _T_802; // @[Mux.scala 46:16:@7007.4]
  wire  _T_803; // @[Mux.scala 46:19:@7008.4]
  wire [10:0] _T_804; // @[Mux.scala 46:16:@7009.4]
  wire  _T_805; // @[Mux.scala 46:19:@7010.4]
  wire [10:0] _T_806; // @[Mux.scala 46:16:@7011.4]
  wire  _T_807; // @[Mux.scala 46:19:@7012.4]
  wire [10:0] _T_808; // @[Mux.scala 46:16:@7013.4]
  wire  _T_809; // @[Mux.scala 46:19:@7014.4]
  wire [10:0] _T_810; // @[Mux.scala 46:16:@7015.4]
  wire  _T_811; // @[Mux.scala 46:19:@7016.4]
  wire [10:0] _T_812; // @[Mux.scala 46:16:@7017.4]
  wire  _T_813; // @[Mux.scala 46:19:@7018.4]
  wire [10:0] _T_814; // @[Mux.scala 46:16:@7019.4]
  wire  _T_815; // @[Mux.scala 46:19:@7020.4]
  wire [10:0] _T_816; // @[Mux.scala 46:16:@7021.4]
  wire  _T_817; // @[Mux.scala 46:19:@7022.4]
  wire [10:0] _T_818; // @[Mux.scala 46:16:@7023.4]
  wire  _T_819; // @[Mux.scala 46:19:@7024.4]
  wire [10:0] _T_820; // @[Mux.scala 46:16:@7025.4]
  wire  _T_821; // @[Mux.scala 46:19:@7026.4]
  wire [10:0] _T_822; // @[Mux.scala 46:16:@7027.4]
  wire  _T_823; // @[Mux.scala 46:19:@7028.4]
  wire [10:0] _T_824; // @[Mux.scala 46:16:@7029.4]
  wire  _T_825; // @[Mux.scala 46:19:@7030.4]
  wire [10:0] _T_826; // @[Mux.scala 46:16:@7031.4]
  wire  _T_827; // @[Mux.scala 46:19:@7032.4]
  wire [10:0] _T_828; // @[Mux.scala 46:16:@7033.4]
  wire  _T_829; // @[Mux.scala 46:19:@7034.4]
  wire [10:0] _T_830; // @[Mux.scala 46:16:@7035.4]
  wire  _T_831; // @[Mux.scala 46:19:@7036.4]
  wire [10:0] _T_832; // @[Mux.scala 46:16:@7037.4]
  wire  _T_833; // @[Mux.scala 46:19:@7038.4]
  wire [10:0] _T_834; // @[Mux.scala 46:16:@7039.4]
  wire  _T_835; // @[Mux.scala 46:19:@7040.4]
  wire [10:0] _T_836; // @[Mux.scala 46:16:@7041.4]
  wire  _T_837; // @[Mux.scala 46:19:@7042.4]
  wire [10:0] _T_838; // @[Mux.scala 46:16:@7043.4]
  wire  _T_839; // @[Mux.scala 46:19:@7044.4]
  wire [10:0] _T_840; // @[Mux.scala 46:16:@7045.4]
  wire  _T_841; // @[Mux.scala 46:19:@7046.4]
  wire [10:0] _T_842; // @[Mux.scala 46:16:@7047.4]
  wire  _T_843; // @[Mux.scala 46:19:@7048.4]
  wire [10:0] _T_844; // @[Mux.scala 46:16:@7049.4]
  wire  _T_845; // @[Mux.scala 46:19:@7050.4]
  wire [10:0] _T_846; // @[Mux.scala 46:16:@7051.4]
  wire  _T_847; // @[Mux.scala 46:19:@7052.4]
  wire [10:0] _T_848; // @[Mux.scala 46:16:@7053.4]
  wire  _T_849; // @[Mux.scala 46:19:@7054.4]
  wire [10:0] _T_850; // @[Mux.scala 46:16:@7055.4]
  wire  _T_851; // @[Mux.scala 46:19:@7056.4]
  wire [10:0] _T_852; // @[Mux.scala 46:16:@7057.4]
  wire  _T_853; // @[Mux.scala 46:19:@7058.4]
  wire [10:0] _T_854; // @[Mux.scala 46:16:@7059.4]
  wire  _T_855; // @[Mux.scala 46:19:@7060.4]
  wire [10:0] _T_856; // @[Mux.scala 46:16:@7061.4]
  wire  _T_857; // @[Mux.scala 46:19:@7062.4]
  wire [10:0] _T_858; // @[Mux.scala 46:16:@7063.4]
  wire  _T_859; // @[Mux.scala 46:19:@7064.4]
  wire [10:0] _T_860; // @[Mux.scala 46:16:@7065.4]
  wire  _T_861; // @[Mux.scala 46:19:@7066.4]
  wire [10:0] _T_862; // @[Mux.scala 46:16:@7067.4]
  wire  _T_863; // @[Mux.scala 46:19:@7068.4]
  wire [10:0] _T_864; // @[Mux.scala 46:16:@7069.4]
  wire  _T_865; // @[Mux.scala 46:19:@7070.4]
  wire [10:0] _T_866; // @[Mux.scala 46:16:@7071.4]
  wire  _T_867; // @[Mux.scala 46:19:@7072.4]
  wire [10:0] _T_868; // @[Mux.scala 46:16:@7073.4]
  wire  _T_869; // @[Mux.scala 46:19:@7074.4]
  wire [10:0] _T_870; // @[Mux.scala 46:16:@7075.4]
  wire  _T_871; // @[Mux.scala 46:19:@7076.4]
  wire [10:0] _T_872; // @[Mux.scala 46:16:@7077.4]
  wire  _T_873; // @[Mux.scala 46:19:@7078.4]
  wire [10:0] _T_874; // @[Mux.scala 46:16:@7079.4]
  wire  _T_875; // @[Mux.scala 46:19:@7080.4]
  wire [10:0] _T_876; // @[Mux.scala 46:16:@7081.4]
  wire  _T_877; // @[Mux.scala 46:19:@7082.4]
  wire [10:0] _T_878; // @[Mux.scala 46:16:@7083.4]
  wire  _T_879; // @[Mux.scala 46:19:@7084.4]
  wire [10:0] _T_880; // @[Mux.scala 46:16:@7085.4]
  wire  _T_881; // @[Mux.scala 46:19:@7086.4]
  wire [10:0] _T_882; // @[Mux.scala 46:16:@7087.4]
  wire  _T_883; // @[Mux.scala 46:19:@7088.4]
  wire [10:0] _T_884; // @[Mux.scala 46:16:@7089.4]
  wire  _T_885; // @[Mux.scala 46:19:@7090.4]
  wire [10:0] _T_886; // @[Mux.scala 46:16:@7091.4]
  wire  _T_887; // @[Mux.scala 46:19:@7092.4]
  wire [10:0] _T_888; // @[Mux.scala 46:16:@7093.4]
  wire  _T_889; // @[Mux.scala 46:19:@7094.4]
  wire [10:0] _T_890; // @[Mux.scala 46:16:@7095.4]
  wire  _T_891; // @[Mux.scala 46:19:@7096.4]
  wire [10:0] _T_892; // @[Mux.scala 46:16:@7097.4]
  wire  _T_893; // @[Mux.scala 46:19:@7098.4]
  wire [10:0] _T_894; // @[Mux.scala 46:16:@7099.4]
  wire  _T_895; // @[Mux.scala 46:19:@7100.4]
  wire [10:0] _T_896; // @[Mux.scala 46:16:@7101.4]
  wire  _T_897; // @[Mux.scala 46:19:@7102.4]
  wire [10:0] _T_898; // @[Mux.scala 46:16:@7103.4]
  wire  _T_899; // @[Mux.scala 46:19:@7104.4]
  wire [10:0] _T_900; // @[Mux.scala 46:16:@7105.4]
  wire  _T_901; // @[Mux.scala 46:19:@7106.4]
  wire [10:0] _T_902; // @[Mux.scala 46:16:@7107.4]
  wire  _T_903; // @[Mux.scala 46:19:@7108.4]
  wire [10:0] _T_904; // @[Mux.scala 46:16:@7109.4]
  wire  _T_905; // @[Mux.scala 46:19:@7110.4]
  wire [10:0] _T_906; // @[Mux.scala 46:16:@7111.4]
  wire  _T_907; // @[Mux.scala 46:19:@7112.4]
  wire [10:0] _T_908; // @[Mux.scala 46:16:@7113.4]
  wire  _T_909; // @[Mux.scala 46:19:@7114.4]
  wire [10:0] _T_910; // @[Mux.scala 46:16:@7115.4]
  wire  _T_911; // @[Mux.scala 46:19:@7116.4]
  wire [10:0] _T_912; // @[Mux.scala 46:16:@7117.4]
  wire  _T_913; // @[Mux.scala 46:19:@7118.4]
  wire [10:0] _T_914; // @[Mux.scala 46:16:@7119.4]
  wire  _T_915; // @[Mux.scala 46:19:@7120.4]
  wire [10:0] _T_916; // @[Mux.scala 46:16:@7121.4]
  wire  _T_917; // @[Mux.scala 46:19:@7122.4]
  wire [10:0] _T_918; // @[Mux.scala 46:16:@7123.4]
  wire  _T_919; // @[Mux.scala 46:19:@7124.4]
  wire [10:0] _T_920; // @[Mux.scala 46:16:@7125.4]
  wire  _T_921; // @[Mux.scala 46:19:@7126.4]
  wire [10:0] _T_922; // @[Mux.scala 46:16:@7127.4]
  wire  _T_923; // @[Mux.scala 46:19:@7128.4]
  wire [10:0] _T_924; // @[Mux.scala 46:16:@7129.4]
  wire  _T_925; // @[Mux.scala 46:19:@7130.4]
  assign _T_669 = 8'h80 == io_ra; // @[Mux.scala 46:19:@6874.4]
  assign _T_670 = _T_669 ? io_di : 11'h0; // @[Mux.scala 46:16:@6875.4]
  assign _T_671 = 8'h7f == io_ra; // @[Mux.scala 46:19:@6876.4]
  assign _T_672 = _T_671 ? 11'h0 : _T_670; // @[Mux.scala 46:16:@6877.4]
  assign _T_673 = 8'h7e == io_ra; // @[Mux.scala 46:19:@6878.4]
  assign _T_674 = _T_673 ? 11'h0 : _T_672; // @[Mux.scala 46:16:@6879.4]
  assign _T_675 = 8'h7d == io_ra; // @[Mux.scala 46:19:@6880.4]
  assign _T_676 = _T_675 ? 11'h0 : _T_674; // @[Mux.scala 46:16:@6881.4]
  assign _T_677 = 8'h7c == io_ra; // @[Mux.scala 46:19:@6882.4]
  assign _T_678 = _T_677 ? 11'h0 : _T_676; // @[Mux.scala 46:16:@6883.4]
  assign _T_679 = 8'h7b == io_ra; // @[Mux.scala 46:19:@6884.4]
  assign _T_680 = _T_679 ? 11'h0 : _T_678; // @[Mux.scala 46:16:@6885.4]
  assign _T_681 = 8'h7a == io_ra; // @[Mux.scala 46:19:@6886.4]
  assign _T_682 = _T_681 ? 11'h0 : _T_680; // @[Mux.scala 46:16:@6887.4]
  assign _T_683 = 8'h79 == io_ra; // @[Mux.scala 46:19:@6888.4]
  assign _T_684 = _T_683 ? 11'h0 : _T_682; // @[Mux.scala 46:16:@6889.4]
  assign _T_685 = 8'h78 == io_ra; // @[Mux.scala 46:19:@6890.4]
  assign _T_686 = _T_685 ? 11'h0 : _T_684; // @[Mux.scala 46:16:@6891.4]
  assign _T_687 = 8'h77 == io_ra; // @[Mux.scala 46:19:@6892.4]
  assign _T_688 = _T_687 ? 11'h0 : _T_686; // @[Mux.scala 46:16:@6893.4]
  assign _T_689 = 8'h76 == io_ra; // @[Mux.scala 46:19:@6894.4]
  assign _T_690 = _T_689 ? 11'h0 : _T_688; // @[Mux.scala 46:16:@6895.4]
  assign _T_691 = 8'h75 == io_ra; // @[Mux.scala 46:19:@6896.4]
  assign _T_692 = _T_691 ? 11'h0 : _T_690; // @[Mux.scala 46:16:@6897.4]
  assign _T_693 = 8'h74 == io_ra; // @[Mux.scala 46:19:@6898.4]
  assign _T_694 = _T_693 ? 11'h0 : _T_692; // @[Mux.scala 46:16:@6899.4]
  assign _T_695 = 8'h73 == io_ra; // @[Mux.scala 46:19:@6900.4]
  assign _T_696 = _T_695 ? 11'h0 : _T_694; // @[Mux.scala 46:16:@6901.4]
  assign _T_697 = 8'h72 == io_ra; // @[Mux.scala 46:19:@6902.4]
  assign _T_698 = _T_697 ? 11'h0 : _T_696; // @[Mux.scala 46:16:@6903.4]
  assign _T_699 = 8'h71 == io_ra; // @[Mux.scala 46:19:@6904.4]
  assign _T_700 = _T_699 ? 11'h0 : _T_698; // @[Mux.scala 46:16:@6905.4]
  assign _T_701 = 8'h70 == io_ra; // @[Mux.scala 46:19:@6906.4]
  assign _T_702 = _T_701 ? 11'h0 : _T_700; // @[Mux.scala 46:16:@6907.4]
  assign _T_703 = 8'h6f == io_ra; // @[Mux.scala 46:19:@6908.4]
  assign _T_704 = _T_703 ? 11'h0 : _T_702; // @[Mux.scala 46:16:@6909.4]
  assign _T_705 = 8'h6e == io_ra; // @[Mux.scala 46:19:@6910.4]
  assign _T_706 = _T_705 ? 11'h0 : _T_704; // @[Mux.scala 46:16:@6911.4]
  assign _T_707 = 8'h6d == io_ra; // @[Mux.scala 46:19:@6912.4]
  assign _T_708 = _T_707 ? 11'h0 : _T_706; // @[Mux.scala 46:16:@6913.4]
  assign _T_709 = 8'h6c == io_ra; // @[Mux.scala 46:19:@6914.4]
  assign _T_710 = _T_709 ? 11'h0 : _T_708; // @[Mux.scala 46:16:@6915.4]
  assign _T_711 = 8'h6b == io_ra; // @[Mux.scala 46:19:@6916.4]
  assign _T_712 = _T_711 ? 11'h0 : _T_710; // @[Mux.scala 46:16:@6917.4]
  assign _T_713 = 8'h6a == io_ra; // @[Mux.scala 46:19:@6918.4]
  assign _T_714 = _T_713 ? 11'h0 : _T_712; // @[Mux.scala 46:16:@6919.4]
  assign _T_715 = 8'h69 == io_ra; // @[Mux.scala 46:19:@6920.4]
  assign _T_716 = _T_715 ? 11'h0 : _T_714; // @[Mux.scala 46:16:@6921.4]
  assign _T_717 = 8'h68 == io_ra; // @[Mux.scala 46:19:@6922.4]
  assign _T_718 = _T_717 ? 11'h0 : _T_716; // @[Mux.scala 46:16:@6923.4]
  assign _T_719 = 8'h67 == io_ra; // @[Mux.scala 46:19:@6924.4]
  assign _T_720 = _T_719 ? 11'h0 : _T_718; // @[Mux.scala 46:16:@6925.4]
  assign _T_721 = 8'h66 == io_ra; // @[Mux.scala 46:19:@6926.4]
  assign _T_722 = _T_721 ? 11'h0 : _T_720; // @[Mux.scala 46:16:@6927.4]
  assign _T_723 = 8'h65 == io_ra; // @[Mux.scala 46:19:@6928.4]
  assign _T_724 = _T_723 ? 11'h0 : _T_722; // @[Mux.scala 46:16:@6929.4]
  assign _T_725 = 8'h64 == io_ra; // @[Mux.scala 46:19:@6930.4]
  assign _T_726 = _T_725 ? 11'h0 : _T_724; // @[Mux.scala 46:16:@6931.4]
  assign _T_727 = 8'h63 == io_ra; // @[Mux.scala 46:19:@6932.4]
  assign _T_728 = _T_727 ? 11'h0 : _T_726; // @[Mux.scala 46:16:@6933.4]
  assign _T_729 = 8'h62 == io_ra; // @[Mux.scala 46:19:@6934.4]
  assign _T_730 = _T_729 ? 11'h0 : _T_728; // @[Mux.scala 46:16:@6935.4]
  assign _T_731 = 8'h61 == io_ra; // @[Mux.scala 46:19:@6936.4]
  assign _T_732 = _T_731 ? 11'h0 : _T_730; // @[Mux.scala 46:16:@6937.4]
  assign _T_733 = 8'h60 == io_ra; // @[Mux.scala 46:19:@6938.4]
  assign _T_734 = _T_733 ? 11'h0 : _T_732; // @[Mux.scala 46:16:@6939.4]
  assign _T_735 = 8'h5f == io_ra; // @[Mux.scala 46:19:@6940.4]
  assign _T_736 = _T_735 ? 11'h0 : _T_734; // @[Mux.scala 46:16:@6941.4]
  assign _T_737 = 8'h5e == io_ra; // @[Mux.scala 46:19:@6942.4]
  assign _T_738 = _T_737 ? 11'h0 : _T_736; // @[Mux.scala 46:16:@6943.4]
  assign _T_739 = 8'h5d == io_ra; // @[Mux.scala 46:19:@6944.4]
  assign _T_740 = _T_739 ? 11'h0 : _T_738; // @[Mux.scala 46:16:@6945.4]
  assign _T_741 = 8'h5c == io_ra; // @[Mux.scala 46:19:@6946.4]
  assign _T_742 = _T_741 ? 11'h0 : _T_740; // @[Mux.scala 46:16:@6947.4]
  assign _T_743 = 8'h5b == io_ra; // @[Mux.scala 46:19:@6948.4]
  assign _T_744 = _T_743 ? 11'h0 : _T_742; // @[Mux.scala 46:16:@6949.4]
  assign _T_745 = 8'h5a == io_ra; // @[Mux.scala 46:19:@6950.4]
  assign _T_746 = _T_745 ? 11'h0 : _T_744; // @[Mux.scala 46:16:@6951.4]
  assign _T_747 = 8'h59 == io_ra; // @[Mux.scala 46:19:@6952.4]
  assign _T_748 = _T_747 ? 11'h0 : _T_746; // @[Mux.scala 46:16:@6953.4]
  assign _T_749 = 8'h58 == io_ra; // @[Mux.scala 46:19:@6954.4]
  assign _T_750 = _T_749 ? 11'h0 : _T_748; // @[Mux.scala 46:16:@6955.4]
  assign _T_751 = 8'h57 == io_ra; // @[Mux.scala 46:19:@6956.4]
  assign _T_752 = _T_751 ? 11'h0 : _T_750; // @[Mux.scala 46:16:@6957.4]
  assign _T_753 = 8'h56 == io_ra; // @[Mux.scala 46:19:@6958.4]
  assign _T_754 = _T_753 ? 11'h0 : _T_752; // @[Mux.scala 46:16:@6959.4]
  assign _T_755 = 8'h55 == io_ra; // @[Mux.scala 46:19:@6960.4]
  assign _T_756 = _T_755 ? 11'h0 : _T_754; // @[Mux.scala 46:16:@6961.4]
  assign _T_757 = 8'h54 == io_ra; // @[Mux.scala 46:19:@6962.4]
  assign _T_758 = _T_757 ? 11'h0 : _T_756; // @[Mux.scala 46:16:@6963.4]
  assign _T_759 = 8'h53 == io_ra; // @[Mux.scala 46:19:@6964.4]
  assign _T_760 = _T_759 ? 11'h0 : _T_758; // @[Mux.scala 46:16:@6965.4]
  assign _T_761 = 8'h52 == io_ra; // @[Mux.scala 46:19:@6966.4]
  assign _T_762 = _T_761 ? 11'h0 : _T_760; // @[Mux.scala 46:16:@6967.4]
  assign _T_763 = 8'h51 == io_ra; // @[Mux.scala 46:19:@6968.4]
  assign _T_764 = _T_763 ? 11'h0 : _T_762; // @[Mux.scala 46:16:@6969.4]
  assign _T_765 = 8'h50 == io_ra; // @[Mux.scala 46:19:@6970.4]
  assign _T_766 = _T_765 ? 11'h0 : _T_764; // @[Mux.scala 46:16:@6971.4]
  assign _T_767 = 8'h4f == io_ra; // @[Mux.scala 46:19:@6972.4]
  assign _T_768 = _T_767 ? 11'h0 : _T_766; // @[Mux.scala 46:16:@6973.4]
  assign _T_769 = 8'h4e == io_ra; // @[Mux.scala 46:19:@6974.4]
  assign _T_770 = _T_769 ? 11'h0 : _T_768; // @[Mux.scala 46:16:@6975.4]
  assign _T_771 = 8'h4d == io_ra; // @[Mux.scala 46:19:@6976.4]
  assign _T_772 = _T_771 ? 11'h0 : _T_770; // @[Mux.scala 46:16:@6977.4]
  assign _T_773 = 8'h4c == io_ra; // @[Mux.scala 46:19:@6978.4]
  assign _T_774 = _T_773 ? 11'h0 : _T_772; // @[Mux.scala 46:16:@6979.4]
  assign _T_775 = 8'h4b == io_ra; // @[Mux.scala 46:19:@6980.4]
  assign _T_776 = _T_775 ? 11'h0 : _T_774; // @[Mux.scala 46:16:@6981.4]
  assign _T_777 = 8'h4a == io_ra; // @[Mux.scala 46:19:@6982.4]
  assign _T_778 = _T_777 ? 11'h0 : _T_776; // @[Mux.scala 46:16:@6983.4]
  assign _T_779 = 8'h49 == io_ra; // @[Mux.scala 46:19:@6984.4]
  assign _T_780 = _T_779 ? 11'h0 : _T_778; // @[Mux.scala 46:16:@6985.4]
  assign _T_781 = 8'h48 == io_ra; // @[Mux.scala 46:19:@6986.4]
  assign _T_782 = _T_781 ? 11'h0 : _T_780; // @[Mux.scala 46:16:@6987.4]
  assign _T_783 = 8'h47 == io_ra; // @[Mux.scala 46:19:@6988.4]
  assign _T_784 = _T_783 ? 11'h0 : _T_782; // @[Mux.scala 46:16:@6989.4]
  assign _T_785 = 8'h46 == io_ra; // @[Mux.scala 46:19:@6990.4]
  assign _T_786 = _T_785 ? 11'h0 : _T_784; // @[Mux.scala 46:16:@6991.4]
  assign _T_787 = 8'h45 == io_ra; // @[Mux.scala 46:19:@6992.4]
  assign _T_788 = _T_787 ? 11'h0 : _T_786; // @[Mux.scala 46:16:@6993.4]
  assign _T_789 = 8'h44 == io_ra; // @[Mux.scala 46:19:@6994.4]
  assign _T_790 = _T_789 ? 11'h0 : _T_788; // @[Mux.scala 46:16:@6995.4]
  assign _T_791 = 8'h43 == io_ra; // @[Mux.scala 46:19:@6996.4]
  assign _T_792 = _T_791 ? 11'h0 : _T_790; // @[Mux.scala 46:16:@6997.4]
  assign _T_793 = 8'h42 == io_ra; // @[Mux.scala 46:19:@6998.4]
  assign _T_794 = _T_793 ? 11'h0 : _T_792; // @[Mux.scala 46:16:@6999.4]
  assign _T_795 = 8'h41 == io_ra; // @[Mux.scala 46:19:@7000.4]
  assign _T_796 = _T_795 ? 11'h0 : _T_794; // @[Mux.scala 46:16:@7001.4]
  assign _T_797 = 8'h40 == io_ra; // @[Mux.scala 46:19:@7002.4]
  assign _T_798 = _T_797 ? 11'h0 : _T_796; // @[Mux.scala 46:16:@7003.4]
  assign _T_799 = 8'h3f == io_ra; // @[Mux.scala 46:19:@7004.4]
  assign _T_800 = _T_799 ? 11'h0 : _T_798; // @[Mux.scala 46:16:@7005.4]
  assign _T_801 = 8'h3e == io_ra; // @[Mux.scala 46:19:@7006.4]
  assign _T_802 = _T_801 ? 11'h0 : _T_800; // @[Mux.scala 46:16:@7007.4]
  assign _T_803 = 8'h3d == io_ra; // @[Mux.scala 46:19:@7008.4]
  assign _T_804 = _T_803 ? 11'h0 : _T_802; // @[Mux.scala 46:16:@7009.4]
  assign _T_805 = 8'h3c == io_ra; // @[Mux.scala 46:19:@7010.4]
  assign _T_806 = _T_805 ? 11'h0 : _T_804; // @[Mux.scala 46:16:@7011.4]
  assign _T_807 = 8'h3b == io_ra; // @[Mux.scala 46:19:@7012.4]
  assign _T_808 = _T_807 ? 11'h0 : _T_806; // @[Mux.scala 46:16:@7013.4]
  assign _T_809 = 8'h3a == io_ra; // @[Mux.scala 46:19:@7014.4]
  assign _T_810 = _T_809 ? 11'h0 : _T_808; // @[Mux.scala 46:16:@7015.4]
  assign _T_811 = 8'h39 == io_ra; // @[Mux.scala 46:19:@7016.4]
  assign _T_812 = _T_811 ? 11'h0 : _T_810; // @[Mux.scala 46:16:@7017.4]
  assign _T_813 = 8'h38 == io_ra; // @[Mux.scala 46:19:@7018.4]
  assign _T_814 = _T_813 ? 11'h0 : _T_812; // @[Mux.scala 46:16:@7019.4]
  assign _T_815 = 8'h37 == io_ra; // @[Mux.scala 46:19:@7020.4]
  assign _T_816 = _T_815 ? 11'h0 : _T_814; // @[Mux.scala 46:16:@7021.4]
  assign _T_817 = 8'h36 == io_ra; // @[Mux.scala 46:19:@7022.4]
  assign _T_818 = _T_817 ? 11'h0 : _T_816; // @[Mux.scala 46:16:@7023.4]
  assign _T_819 = 8'h35 == io_ra; // @[Mux.scala 46:19:@7024.4]
  assign _T_820 = _T_819 ? 11'h0 : _T_818; // @[Mux.scala 46:16:@7025.4]
  assign _T_821 = 8'h34 == io_ra; // @[Mux.scala 46:19:@7026.4]
  assign _T_822 = _T_821 ? 11'h0 : _T_820; // @[Mux.scala 46:16:@7027.4]
  assign _T_823 = 8'h33 == io_ra; // @[Mux.scala 46:19:@7028.4]
  assign _T_824 = _T_823 ? 11'h0 : _T_822; // @[Mux.scala 46:16:@7029.4]
  assign _T_825 = 8'h32 == io_ra; // @[Mux.scala 46:19:@7030.4]
  assign _T_826 = _T_825 ? 11'h0 : _T_824; // @[Mux.scala 46:16:@7031.4]
  assign _T_827 = 8'h31 == io_ra; // @[Mux.scala 46:19:@7032.4]
  assign _T_828 = _T_827 ? 11'h0 : _T_826; // @[Mux.scala 46:16:@7033.4]
  assign _T_829 = 8'h30 == io_ra; // @[Mux.scala 46:19:@7034.4]
  assign _T_830 = _T_829 ? 11'h0 : _T_828; // @[Mux.scala 46:16:@7035.4]
  assign _T_831 = 8'h2f == io_ra; // @[Mux.scala 46:19:@7036.4]
  assign _T_832 = _T_831 ? 11'h0 : _T_830; // @[Mux.scala 46:16:@7037.4]
  assign _T_833 = 8'h2e == io_ra; // @[Mux.scala 46:19:@7038.4]
  assign _T_834 = _T_833 ? 11'h0 : _T_832; // @[Mux.scala 46:16:@7039.4]
  assign _T_835 = 8'h2d == io_ra; // @[Mux.scala 46:19:@7040.4]
  assign _T_836 = _T_835 ? 11'h0 : _T_834; // @[Mux.scala 46:16:@7041.4]
  assign _T_837 = 8'h2c == io_ra; // @[Mux.scala 46:19:@7042.4]
  assign _T_838 = _T_837 ? 11'h0 : _T_836; // @[Mux.scala 46:16:@7043.4]
  assign _T_839 = 8'h2b == io_ra; // @[Mux.scala 46:19:@7044.4]
  assign _T_840 = _T_839 ? 11'h0 : _T_838; // @[Mux.scala 46:16:@7045.4]
  assign _T_841 = 8'h2a == io_ra; // @[Mux.scala 46:19:@7046.4]
  assign _T_842 = _T_841 ? 11'h0 : _T_840; // @[Mux.scala 46:16:@7047.4]
  assign _T_843 = 8'h29 == io_ra; // @[Mux.scala 46:19:@7048.4]
  assign _T_844 = _T_843 ? 11'h0 : _T_842; // @[Mux.scala 46:16:@7049.4]
  assign _T_845 = 8'h28 == io_ra; // @[Mux.scala 46:19:@7050.4]
  assign _T_846 = _T_845 ? 11'h0 : _T_844; // @[Mux.scala 46:16:@7051.4]
  assign _T_847 = 8'h27 == io_ra; // @[Mux.scala 46:19:@7052.4]
  assign _T_848 = _T_847 ? 11'h0 : _T_846; // @[Mux.scala 46:16:@7053.4]
  assign _T_849 = 8'h26 == io_ra; // @[Mux.scala 46:19:@7054.4]
  assign _T_850 = _T_849 ? 11'h0 : _T_848; // @[Mux.scala 46:16:@7055.4]
  assign _T_851 = 8'h25 == io_ra; // @[Mux.scala 46:19:@7056.4]
  assign _T_852 = _T_851 ? 11'h0 : _T_850; // @[Mux.scala 46:16:@7057.4]
  assign _T_853 = 8'h24 == io_ra; // @[Mux.scala 46:19:@7058.4]
  assign _T_854 = _T_853 ? 11'h0 : _T_852; // @[Mux.scala 46:16:@7059.4]
  assign _T_855 = 8'h23 == io_ra; // @[Mux.scala 46:19:@7060.4]
  assign _T_856 = _T_855 ? 11'h0 : _T_854; // @[Mux.scala 46:16:@7061.4]
  assign _T_857 = 8'h22 == io_ra; // @[Mux.scala 46:19:@7062.4]
  assign _T_858 = _T_857 ? 11'h0 : _T_856; // @[Mux.scala 46:16:@7063.4]
  assign _T_859 = 8'h21 == io_ra; // @[Mux.scala 46:19:@7064.4]
  assign _T_860 = _T_859 ? 11'h0 : _T_858; // @[Mux.scala 46:16:@7065.4]
  assign _T_861 = 8'h20 == io_ra; // @[Mux.scala 46:19:@7066.4]
  assign _T_862 = _T_861 ? 11'h0 : _T_860; // @[Mux.scala 46:16:@7067.4]
  assign _T_863 = 8'h1f == io_ra; // @[Mux.scala 46:19:@7068.4]
  assign _T_864 = _T_863 ? 11'h0 : _T_862; // @[Mux.scala 46:16:@7069.4]
  assign _T_865 = 8'h1e == io_ra; // @[Mux.scala 46:19:@7070.4]
  assign _T_866 = _T_865 ? 11'h0 : _T_864; // @[Mux.scala 46:16:@7071.4]
  assign _T_867 = 8'h1d == io_ra; // @[Mux.scala 46:19:@7072.4]
  assign _T_868 = _T_867 ? 11'h0 : _T_866; // @[Mux.scala 46:16:@7073.4]
  assign _T_869 = 8'h1c == io_ra; // @[Mux.scala 46:19:@7074.4]
  assign _T_870 = _T_869 ? 11'h0 : _T_868; // @[Mux.scala 46:16:@7075.4]
  assign _T_871 = 8'h1b == io_ra; // @[Mux.scala 46:19:@7076.4]
  assign _T_872 = _T_871 ? 11'h0 : _T_870; // @[Mux.scala 46:16:@7077.4]
  assign _T_873 = 8'h1a == io_ra; // @[Mux.scala 46:19:@7078.4]
  assign _T_874 = _T_873 ? 11'h0 : _T_872; // @[Mux.scala 46:16:@7079.4]
  assign _T_875 = 8'h19 == io_ra; // @[Mux.scala 46:19:@7080.4]
  assign _T_876 = _T_875 ? 11'h0 : _T_874; // @[Mux.scala 46:16:@7081.4]
  assign _T_877 = 8'h18 == io_ra; // @[Mux.scala 46:19:@7082.4]
  assign _T_878 = _T_877 ? 11'h0 : _T_876; // @[Mux.scala 46:16:@7083.4]
  assign _T_879 = 8'h17 == io_ra; // @[Mux.scala 46:19:@7084.4]
  assign _T_880 = _T_879 ? 11'h0 : _T_878; // @[Mux.scala 46:16:@7085.4]
  assign _T_881 = 8'h16 == io_ra; // @[Mux.scala 46:19:@7086.4]
  assign _T_882 = _T_881 ? 11'h0 : _T_880; // @[Mux.scala 46:16:@7087.4]
  assign _T_883 = 8'h15 == io_ra; // @[Mux.scala 46:19:@7088.4]
  assign _T_884 = _T_883 ? 11'h0 : _T_882; // @[Mux.scala 46:16:@7089.4]
  assign _T_885 = 8'h14 == io_ra; // @[Mux.scala 46:19:@7090.4]
  assign _T_886 = _T_885 ? 11'h0 : _T_884; // @[Mux.scala 46:16:@7091.4]
  assign _T_887 = 8'h13 == io_ra; // @[Mux.scala 46:19:@7092.4]
  assign _T_888 = _T_887 ? 11'h0 : _T_886; // @[Mux.scala 46:16:@7093.4]
  assign _T_889 = 8'h12 == io_ra; // @[Mux.scala 46:19:@7094.4]
  assign _T_890 = _T_889 ? 11'h0 : _T_888; // @[Mux.scala 46:16:@7095.4]
  assign _T_891 = 8'h11 == io_ra; // @[Mux.scala 46:19:@7096.4]
  assign _T_892 = _T_891 ? 11'h0 : _T_890; // @[Mux.scala 46:16:@7097.4]
  assign _T_893 = 8'h10 == io_ra; // @[Mux.scala 46:19:@7098.4]
  assign _T_894 = _T_893 ? 11'h0 : _T_892; // @[Mux.scala 46:16:@7099.4]
  assign _T_895 = 8'hf == io_ra; // @[Mux.scala 46:19:@7100.4]
  assign _T_896 = _T_895 ? 11'h0 : _T_894; // @[Mux.scala 46:16:@7101.4]
  assign _T_897 = 8'he == io_ra; // @[Mux.scala 46:19:@7102.4]
  assign _T_898 = _T_897 ? 11'h0 : _T_896; // @[Mux.scala 46:16:@7103.4]
  assign _T_899 = 8'hd == io_ra; // @[Mux.scala 46:19:@7104.4]
  assign _T_900 = _T_899 ? 11'h0 : _T_898; // @[Mux.scala 46:16:@7105.4]
  assign _T_901 = 8'hc == io_ra; // @[Mux.scala 46:19:@7106.4]
  assign _T_902 = _T_901 ? 11'h0 : _T_900; // @[Mux.scala 46:16:@7107.4]
  assign _T_903 = 8'hb == io_ra; // @[Mux.scala 46:19:@7108.4]
  assign _T_904 = _T_903 ? 11'h0 : _T_902; // @[Mux.scala 46:16:@7109.4]
  assign _T_905 = 8'ha == io_ra; // @[Mux.scala 46:19:@7110.4]
  assign _T_906 = _T_905 ? 11'h0 : _T_904; // @[Mux.scala 46:16:@7111.4]
  assign _T_907 = 8'h9 == io_ra; // @[Mux.scala 46:19:@7112.4]
  assign _T_908 = _T_907 ? 11'h0 : _T_906; // @[Mux.scala 46:16:@7113.4]
  assign _T_909 = 8'h8 == io_ra; // @[Mux.scala 46:19:@7114.4]
  assign _T_910 = _T_909 ? 11'h0 : _T_908; // @[Mux.scala 46:16:@7115.4]
  assign _T_911 = 8'h7 == io_ra; // @[Mux.scala 46:19:@7116.4]
  assign _T_912 = _T_911 ? 11'h0 : _T_910; // @[Mux.scala 46:16:@7117.4]
  assign _T_913 = 8'h6 == io_ra; // @[Mux.scala 46:19:@7118.4]
  assign _T_914 = _T_913 ? 11'h0 : _T_912; // @[Mux.scala 46:16:@7119.4]
  assign _T_915 = 8'h5 == io_ra; // @[Mux.scala 46:19:@7120.4]
  assign _T_916 = _T_915 ? 11'h0 : _T_914; // @[Mux.scala 46:16:@7121.4]
  assign _T_917 = 8'h4 == io_ra; // @[Mux.scala 46:19:@7122.4]
  assign _T_918 = _T_917 ? 11'h0 : _T_916; // @[Mux.scala 46:16:@7123.4]
  assign _T_919 = 8'h3 == io_ra; // @[Mux.scala 46:19:@7124.4]
  assign _T_920 = _T_919 ? 11'h0 : _T_918; // @[Mux.scala 46:16:@7125.4]
  assign _T_921 = 8'h2 == io_ra; // @[Mux.scala 46:19:@7126.4]
  assign _T_922 = _T_921 ? 11'h0 : _T_920; // @[Mux.scala 46:16:@7127.4]
  assign _T_923 = 8'h1 == io_ra; // @[Mux.scala 46:19:@7128.4]
  assign _T_924 = _T_923 ? 11'h0 : _T_922; // @[Mux.scala 46:16:@7129.4]
  assign _T_925 = 8'h0 == io_ra; // @[Mux.scala 46:19:@7130.4]
  assign io_dout = _T_925 ? 11'h0 : _T_924; // @[nv_flopram.scala 81:13:@7132.4]
endmodule
module NV_NVDLA_fifo_4( // @[:@7134.2]
  input         clock, // @[:@7135.4]
  input         reset, // @[:@7136.4]
  input  [10:0] io_wr_pd, // @[:@7137.4]
  output        io_rd_pvld, // @[:@7137.4]
  input         io_rd_prdy, // @[:@7137.4]
  output [10:0] io_rd_pd // @[:@7137.4]
);
  wire [10:0] nv_flopram_io_di; // @[FIFO.scala 254:29:@7196.4]
  wire [7:0] nv_flopram_io_ra; // @[FIFO.scala 254:29:@7196.4]
  wire [10:0] nv_flopram_io_dout; // @[FIFO.scala 254:29:@7196.4]
  reg [7:0] _T_38; // @[FIFO.scala 186:53:@7154.4]
  reg [31:0] _RAND_0;
  wire [8:0] _T_40; // @[FIFO.scala 190:76:@7155.4]
  wire [8:0] _T_41; // @[FIFO.scala 190:76:@7156.4]
  wire [7:0] _T_42; // @[FIFO.scala 190:76:@7157.4]
  wire  _T_109; // @[FIFO.scala 324:38:@7228.4]
  wire [7:0] _T_48; // @[FIFO.scala 192:32:@7162.4]
  wire [7:0] _GEN_0; // @[FIFO.scala 202:40:@7173.4]
  reg [6:0] _T_71; // @[FIFO.scala 224:63:@7183.4]
  reg [31:0] _RAND_1;
  wire [7:0] _T_73; // @[FIFO.scala 225:42:@7184.4]
  wire [6:0] _T_74; // @[FIFO.scala 225:42:@7185.4]
  wire [6:0] _GEN_2; // @[FIFO.scala 227:29:@7186.4]
  wire  _T_87; // @[FIFO.scala 264:39:@7206.4]
  reg [7:0] _T_94; // @[FIFO.scala 299:53:@7212.4]
  reg [31:0] _RAND_2;
  wire [8:0] _T_96; // @[FIFO.scala 300:74:@7213.4]
  wire [8:0] _T_97; // @[FIFO.scala 300:74:@7214.4]
  wire [7:0] _T_98; // @[FIFO.scala 300:74:@7215.4]
  wire [7:0] _T_104; // @[FIFO.scala 302:32:@7220.4]
  wire [7:0] _GEN_3; // @[FIFO.scala 303:39:@7222.4]
  nv_flopram nv_flopram ( // @[FIFO.scala 254:29:@7196.4]
    .io_di(nv_flopram_io_di),
    .io_ra(nv_flopram_io_ra),
    .io_dout(nv_flopram_io_dout)
  );
  assign _T_40 = _T_38 - 8'h1; // @[FIFO.scala 190:76:@7155.4]
  assign _T_41 = $unsigned(_T_40); // @[FIFO.scala 190:76:@7156.4]
  assign _T_42 = _T_41[7:0]; // @[FIFO.scala 190:76:@7157.4]
  assign _T_109 = io_rd_pvld & io_rd_prdy; // @[FIFO.scala 324:38:@7228.4]
  assign _T_48 = _T_109 ? _T_42 : _T_38; // @[FIFO.scala 192:32:@7162.4]
  assign _GEN_0 = _T_109 ? _T_48 : _T_38; // @[FIFO.scala 202:40:@7173.4]
  assign _T_73 = _T_71 + 7'h1; // @[FIFO.scala 225:42:@7184.4]
  assign _T_74 = _T_71 + 7'h1; // @[FIFO.scala 225:42:@7185.4]
  assign _GEN_2 = _T_109 ? _T_74 : _T_71; // @[FIFO.scala 227:29:@7186.4]
  assign _T_87 = _T_38 == 8'h0; // @[FIFO.scala 264:39:@7206.4]
  assign _T_96 = _T_94 - 8'h1; // @[FIFO.scala 300:74:@7213.4]
  assign _T_97 = $unsigned(_T_96); // @[FIFO.scala 300:74:@7214.4]
  assign _T_98 = _T_97[7:0]; // @[FIFO.scala 300:74:@7215.4]
  assign _T_104 = _T_109 ? _T_98 : _T_94; // @[FIFO.scala 302:32:@7220.4]
  assign _GEN_3 = _T_109 ? _T_104 : _T_94; // @[FIFO.scala 303:39:@7222.4]
  assign io_rd_pvld = _T_94 != 8'h0; // @[FIFO.scala 326:24:@7230.4]
  assign io_rd_pd = nv_flopram_io_dout; // @[FIFO.scala 327:22:@7231.4]
  assign nv_flopram_io_di = io_wr_pd; // @[FIFO.scala 258:23:@7202.4]
  assign nv_flopram_io_ra = _T_87 ? 8'h80 : {{1'd0}, _T_71}; // @[FIFO.scala 264:23:@7208.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_38 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_71 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_94 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_38 <= 8'h0;
    end else begin
      if (_T_109) begin
        if (_T_109) begin
          _T_38 <= _T_42;
        end
      end
    end
    if (reset) begin
      _T_71 <= 7'h0;
    end else begin
      if (_T_109) begin
        _T_71 <= _T_74;
      end
    end
    if (reset) begin
      _T_94 <= 8'h0;
    end else begin
      if (_T_109) begin
        if (_T_109) begin
          _T_94 <= _T_98;
        end
      end
    end
  end
endmodule
module NV_NVDLA_CDMA_IMG_sg( // @[:@7352.2]
  input          reset, // @[:@7354.4]
  input          io_nvdla_core_clk, // @[:@7355.4]
  input          io_img_dat2mcif_rd_req_pd_ready, // @[:@7355.4]
  output         io_img_dat2mcif_rd_req_pd_valid, // @[:@7355.4]
  output [78:0]  io_img_dat2mcif_rd_req_pd_bits, // @[:@7355.4]
  output         io_mcif2img_dat_rd_rsp_pd_ready, // @[:@7355.4]
  input          io_mcif2img_dat_rd_rsp_pd_valid, // @[:@7355.4]
  input  [256:0] io_mcif2img_dat_rd_rsp_pd_bits, // @[:@7355.4]
  input          io_img_dat2cvif_rd_req_pd_ready, // @[:@7355.4]
  output         io_img_dat2cvif_rd_req_pd_valid, // @[:@7355.4]
  output [78:0]  io_img_dat2cvif_rd_req_pd_bits, // @[:@7355.4]
  output         io_cvif2img_dat_rd_rsp_pd_ready, // @[:@7355.4]
  input          io_cvif2img_dat_rd_rsp_pd_valid, // @[:@7355.4]
  input  [256:0] io_cvif2img_dat_rd_rsp_pd_bits, // @[:@7355.4]
  input  [14:0]  io_img2status_dat_entries, // @[:@7355.4]
  input          io_img2status_dat_updt, // @[:@7355.4]
  input  [14:0]  io_status2dma_free_entries, // @[:@7355.4]
  input          io_status2dma_fsm_switch, // @[:@7355.4]
  input          io_is_running, // @[:@7355.4]
  input          io_layer_st, // @[:@7355.4]
  input  [10:0]  io_pixel_order, // @[:@7355.4]
  input          io_pixel_planar, // @[:@7355.4]
  input  [3:0]   io_pixel_planar0_bundle_limit, // @[:@7355.4]
  input  [3:0]   io_pixel_planar0_bundle_limit_1st, // @[:@7355.4]
  input  [4:0]   io_pixel_planar0_byte_sft, // @[:@7355.4]
  input  [4:0]   io_pixel_planar1_byte_sft, // @[:@7355.4]
  input  [3:0]   io_pixel_planar0_lp_burst, // @[:@7355.4]
  input          io_pixel_planar0_lp_vld, // @[:@7355.4]
  input  [3:0]   io_pixel_planar0_rp_burst, // @[:@7355.4]
  input          io_pixel_planar0_rp_vld, // @[:@7355.4]
  input  [13:0]  io_pixel_planar0_width_burst, // @[:@7355.4]
  input  [4:0]   io_pixel_planar1_bundle_limit, // @[:@7355.4]
  input  [4:0]   io_pixel_planar1_bundle_limit_1st, // @[:@7355.4]
  input  [2:0]   io_pixel_planar1_lp_burst, // @[:@7355.4]
  input          io_pixel_planar1_lp_vld, // @[:@7355.4]
  input  [2:0]   io_pixel_planar1_rp_burst, // @[:@7355.4]
  input          io_pixel_planar1_rp_vld, // @[:@7355.4]
  input  [13:0]  io_pixel_planar1_width_burst, // @[:@7355.4]
  input          io_sg2pack_img_pd_ready, // @[:@7355.4]
  output         io_sg2pack_img_pd_valid, // @[:@7355.4]
  output [10:0]  io_sg2pack_img_pd_bits, // @[:@7355.4]
  output [14:0]  io_sg2pack_data_entries, // @[:@7355.4]
  output [14:0]  io_sg2pack_entry_end, // @[:@7355.4]
  output [14:0]  io_sg2pack_entry_mid, // @[:@7355.4]
  output [14:0]  io_sg2pack_entry_st, // @[:@7355.4]
  output [12:0]  io_sg2pack_height_total, // @[:@7355.4]
  output         io_sg2pack_mn_enable, // @[:@7355.4]
  output [3:0]   io_sg2pack_sub_h_end, // @[:@7355.4]
  output [3:0]   io_sg2pack_sub_h_mid, // @[:@7355.4]
  output [3:0]   io_sg2pack_sub_h_st, // @[:@7355.4]
  output         io_sg_is_done, // @[:@7355.4]
  output         io_img2sbuf_p0_wr_addr_valid, // @[:@7355.4]
  output [16:0]  io_img2sbuf_p0_wr_addr_bits, // @[:@7355.4]
  output [255:0] io_img2sbuf_p0_wr_data, // @[:@7355.4]
  input          io_reg2dp_op_en, // @[:@7355.4]
  input  [12:0]  io_reg2dp_datain_height, // @[:@7355.4]
  input          io_reg2dp_datain_ram_type, // @[:@7355.4]
  input  [31:0]  io_reg2dp_datain_addr_high_0, // @[:@7355.4]
  input  [31:0]  io_reg2dp_datain_addr_low_0, // @[:@7355.4]
  input  [31:0]  io_reg2dp_datain_addr_high_1, // @[:@7355.4]
  input  [31:0]  io_reg2dp_datain_addr_low_1, // @[:@7355.4]
  input  [31:0]  io_reg2dp_line_stride, // @[:@7355.4]
  input  [31:0]  io_reg2dp_uv_line_stride, // @[:@7355.4]
  input          io_reg2dp_mean_format, // @[:@7355.4]
  input  [13:0]  io_reg2dp_entries, // @[:@7355.4]
  input          io_reg2dp_dma_en, // @[:@7355.4]
  output [31:0]  io_dp2reg_img_rd_stall, // @[:@7355.4]
  output [31:0]  io_dp2reg_img_rd_latency // @[:@7355.4]
);
  wire  NV_NVDLA_DMAIF_rdreq_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire [78:0] NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type; // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
  wire  NV_NVDLA_DMAIF_rdrsp_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire [256:0] NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
  wire  NV_NVDLA_fifo_clock; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_io_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_io_wr_pvld; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire [10:0] NV_NVDLA_fifo_io_wr_pd; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_io_rd_prdy; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire [10:0] NV_NVDLA_fifo_io_rd_pd; // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
  wire  NV_NVDLA_fifo_1_clock; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire  NV_NVDLA_fifo_1_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire [10:0] NV_NVDLA_fifo_1_io_wr_pd; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire  NV_NVDLA_fifo_1_io_rd_pvld; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire  NV_NVDLA_fifo_1_io_rd_prdy; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire [10:0] NV_NVDLA_fifo_1_io_rd_pd; // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
  wire  NV_COUNTER_STAGE_histogram_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire  NV_COUNTER_STAGE_histogram_io_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_inc; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_clr; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire  NV_COUNTER_STAGE_histogram_io_rd_stall_cen; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire [31:0] NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
  wire  NV_COUNTER_STAGE_histogram_1_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire [8:0] NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
  wire  NV_COUNTER_STAGE_histogram_2_reset; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  wire  NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  wire [31:0] NV_COUNTER_STAGE_histogram_2_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
  reg  _T_157; // @[NV_NVDLA_CDMA_IMG_sg.scala 119:32:@7357.4]
  reg [31:0] _RAND_0;
  reg  _T_160; // @[NV_NVDLA_CDMA_IMG_sg.scala 120:31:@7358.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_163; // @[NV_NVDLA_CDMA_IMG_sg.scala 121:30:@7359.4]
  reg [31:0] _RAND_2;
  reg [12:0] _T_166; // @[NV_NVDLA_CDMA_IMG_sg.scala 122:35:@7360.4]
  reg [31:0] _RAND_3;
  reg [14:0] _T_169; // @[NV_NVDLA_CDMA_IMG_sg.scala 123:31:@7361.4]
  reg [31:0] _RAND_4;
  wire  _T_170; // @[NV_NVDLA_CDMA_IMG_sg.scala 126:44:@7362.4]
  wire  _T_171; // @[NV_NVDLA_CDMA_IMG_sg.scala 126:42:@7363.4]
  wire [13:0] _T_175; // @[NV_NVDLA_CDMA_IMG_sg.scala 131:48:@7368.6]
  wire [14:0] _T_177; // @[NV_NVDLA_CDMA_IMG_sg.scala 133:43:@7371.6]
  wire  _GEN_0; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  wire [13:0] _GEN_1; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  wire [12:0] _GEN_2; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  wire [14:0] _GEN_3; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  reg [3:0] _T_180; // @[NV_NVDLA_CDMA_IMG_sg.scala 139:34:@7374.4]
  reg [31:0] _RAND_5;
  reg [3:0] _T_183; // @[NV_NVDLA_CDMA_IMG_sg.scala 140:35:@7375.4]
  reg [31:0] _RAND_6;
  reg [3:0] _T_186; // @[NV_NVDLA_CDMA_IMG_sg.scala 141:35:@7376.4]
  reg [31:0] _RAND_7;
  reg [14:0] _T_189; // @[NV_NVDLA_CDMA_IMG_sg.scala 142:34:@7377.4]
  reg [31:0] _RAND_8;
  reg [14:0] _T_192; // @[NV_NVDLA_CDMA_IMG_sg.scala 143:35:@7378.4]
  reg [31:0] _RAND_9;
  reg [14:0] _T_195; // @[NV_NVDLA_CDMA_IMG_sg.scala 144:35:@7379.4]
  reg [31:0] _RAND_10;
  wire [9:0] _T_199; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:38:@7380.4]
  wire  _T_201; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:46:@7381.4]
  wire  _T_202; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:25:@7382.4]
  wire [3:0] _T_203; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:67:@7383.4]
  wire  _T_204; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:74:@7384.4]
  wire  _T_205; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:52:@7385.4]
  wire [3:0] _T_214; // @[NV_NVDLA_CDMA_IMG_sg.scala 153:25:@7393.4]
  wire [14:0] _GEN_58; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:38:@7396.4]
  wire [18:0] _T_217; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:38:@7396.4]
  wire [14:0] _T_218; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:53:@7397.4]
  wire [3:0] _GEN_4; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  wire [3:0] _GEN_5; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  wire [3:0] _GEN_6; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  wire [14:0] _GEN_7; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  wire [14:0] _GEN_8; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  wire [14:0] _GEN_9; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  reg [12:0] _T_226; // @[NV_NVDLA_CDMA_IMG_sg.scala 175:33:@7408.4]
  reg [31:0] _RAND_11;
  wire  _T_230; // @[NV_NVDLA_CDMA_IMG_sg.scala 177:42:@7410.4]
  wire  _T_231; // @[NV_NVDLA_CDMA_IMG_sg.scala 177:25:@7411.4]
  wire  _T_232; // @[NV_NVDLA_CDMA_IMG_sg.scala 178:42:@7412.4]
  wire [13:0] _T_235; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:83:@7414.6]
  wire [12:0] _T_236; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:83:@7415.6]
  wire [12:0] _T_237; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:30:@7416.6]
  reg  _T_433; // @[NV_NVDLA_CDMA_IMG_sg.scala 281:28:@7589.4]
  reg [31:0] _RAND_12;
  reg  _T_436; // @[NV_NVDLA_CDMA_IMG_sg.scala 282:31:@7590.4]
  reg [31:0] _RAND_13;
  wire  _T_447; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:32:@7598.4]
  wire  _T_573; // @[NV_NVDLA_CDMA_IMG_sg.scala 379:30:@7720.4 NV_NVDLA_CDMA_IMG_sg.scala 436:20:@7787.4]
  reg  _T_556; // @[NV_NVDLA_CDMA_IMG_sg.scala 348:34:@7695.4]
  reg [31:0] _RAND_14;
  wire  _T_582; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:38:@7724.4]
  wire  _T_575; // @[NV_NVDLA_CDMA_IMG_sg.scala 380:34:@7721.4 NV_NVDLA_CDMA_IMG_sg.scala 473:24:@7827.4]
  wire  _T_583; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:57:@7725.4]
  reg  _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 381:32:@7722.4]
  reg [31:0] _RAND_15;
  wire  _T_584; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:78:@7726.4]
  wire  _T_448; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:46:@7599.4]
  wire  _T_449; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:29:@7600.4]
  reg  _T_240; // @[NV_NVDLA_CDMA_IMG_sg.scala 184:37:@7419.4]
  reg [31:0] _RAND_16;
  wire  _T_417; // @[NV_NVDLA_CDMA_IMG_sg.scala 273:33:@7577.4]
  reg [13:0] _T_267; // @[NV_NVDLA_CDMA_IMG_sg.scala 206:39:@7442.4]
  reg [31:0] _RAND_17;
  reg [3:0] _T_250; // @[NV_NVDLA_CDMA_IMG_sg.scala 193:40:@7428.4]
  reg [31:0] _RAND_18;
  wire [13:0] _GEN_60; // @[NV_NVDLA_CDMA_IMG_sg.scala 213:48:@7452.4]
  wire  _T_280; // @[NV_NVDLA_CDMA_IMG_sg.scala 213:48:@7452.4]
  reg [1:0] _T_270; // @[NV_NVDLA_CDMA_IMG_sg.scala 207:37:@7443.4]
  reg [31:0] _RAND_19;
  wire  _T_293; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:66:@7463.4]
  wire  _T_294; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:44:@7464.4]
  wire  _T_295; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:77:@7465.4]
  wire  _T_296; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:75:@7466.4]
  wire  _T_298; // @[NV_NVDLA_CDMA_IMG_sg.scala 217:69:@7467.4]
  wire  _T_299; // @[NV_NVDLA_CDMA_IMG_sg.scala 217:47:@7468.4]
  wire  _T_300; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:102:@7469.4]
  reg [13:0] _T_337; // @[NV_NVDLA_CDMA_IMG_sg.scala 237:39:@7504.4]
  reg [31:0] _RAND_20;
  reg [4:0] _T_334; // @[NV_NVDLA_CDMA_IMG_sg.scala 236:40:@7503.4]
  reg [31:0] _RAND_21;
  wire [13:0] _GEN_61; // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7510.4]
  wire [14:0] _T_349; // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7510.4]
  wire [14:0] _T_350; // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7511.4]
  wire  _T_354; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:50:@7516.4]
  wire  _T_355; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:79:@7517.4]
  wire  _T_356; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:55:@7518.4]
  reg [1:0] _T_340; // @[NV_NVDLA_CDMA_IMG_sg.scala 238:37:@7505.4]
  reg [31:0] _RAND_22;
  wire  _T_369; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:69:@7529.4]
  wire  _T_370; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:47:@7530.4]
  wire  _T_371; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:80:@7531.4]
  wire  _T_372; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:78:@7532.4]
  wire  _T_374; // @[NV_NVDLA_CDMA_IMG_sg.scala 251:69:@7533.4]
  wire  _T_375; // @[NV_NVDLA_CDMA_IMG_sg.scala 251:47:@7534.4]
  wire  _T_376; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:106:@7535.4]
  wire  _T_418; // @[NV_NVDLA_CDMA_IMG_sg.scala 273:32:@7578.4]
  wire  _T_475; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:57:@7633.4]
  wire  _T_243; // @[NV_NVDLA_CDMA_IMG_sg.scala 186:50:@7421.4]
  wire  _T_476; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:77:@7634.4]
  wire  _T_477; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:39:@7635.4]
  wire [12:0] _GEN_10; // @[NV_NVDLA_CDMA_IMG_sg.scala 180:24:@7413.4]
  wire  _T_244; // @[NV_NVDLA_CDMA_IMG_sg.scala 187:54:@7422.4]
  wire  _T_247; // @[NV_NVDLA_CDMA_IMG_sg.scala 187:35:@7424.4]
  wire [14:0] _T_275; // @[NV_NVDLA_CDMA_IMG_sg.scala 211:57:@7446.4]
  wire [14:0] _T_276; // @[NV_NVDLA_CDMA_IMG_sg.scala 211:57:@7447.4]
  wire  _T_277; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:57:@7448.4]
  wire [3:0] _T_278; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:83:@7449.4]
  wire [3:0] _T_279; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:32:@7450.4]
  wire  _T_301; // @[NV_NVDLA_CDMA_IMG_sg.scala 218:47:@7471.4]
  wire  _T_302; // @[NV_NVDLA_CDMA_IMG_sg.scala 218:74:@7472.4]
  wire [4:0] _T_352; // @[NV_NVDLA_CDMA_IMG_sg.scala 245:83:@7513.4]
  wire [4:0] _T_353; // @[NV_NVDLA_CDMA_IMG_sg.scala 245:32:@7514.4]
  wire  _T_377; // @[NV_NVDLA_CDMA_IMG_sg.scala 252:50:@7536.4]
  wire  _T_378; // @[NV_NVDLA_CDMA_IMG_sg.scala 252:77:@7537.4]
  wire  _T_420; // @[NV_NVDLA_CDMA_IMG_sg.scala 274:32:@7580.4]
  wire  _T_473; // @[NV_NVDLA_CDMA_IMG_sg.scala 302:61:@7630.4]
  wire  _T_474; // @[NV_NVDLA_CDMA_IMG_sg.scala 302:43:@7631.4]
  wire  _GEN_11; // @[NV_NVDLA_CDMA_IMG_sg.scala 189:28:@7425.4]
  wire  _T_259; // @[NV_NVDLA_CDMA_IMG_sg.scala 200:55:@7434.6]
  wire [4:0] _T_260; // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7435.6]
  wire [4:0] _T_261; // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7436.6]
  wire [3:0] _T_262; // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7437.6]
  wire [3:0] _T_263; // @[NV_NVDLA_CDMA_IMG_sg.scala 201:37:@7438.6]
  wire [3:0] _T_264; // @[NV_NVDLA_CDMA_IMG_sg.scala 200:37:@7439.6]
  wire  _T_453; // @[NV_NVDLA_CDMA_IMG_sg.scala 296:63:@7606.4]
  wire  _T_454; // @[NV_NVDLA_CDMA_IMG_sg.scala 296:45:@7607.4]
  wire [3:0] _GEN_12; // @[NV_NVDLA_CDMA_IMG_sg.scala 199:30:@7433.4]
  wire [13:0] _GEN_64; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:50:@7454.4]
  wire  _T_281; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:50:@7454.4]
  wire  _T_283; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:101:@7455.4]
  wire  _T_284; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:80:@7456.4]
  wire  _T_285; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:50:@7457.4]
  wire  _T_288; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:83:@7459.4]
  wire  _T_289; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:114:@7460.4]
  wire  _T_290; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:112:@7461.4]
  wire  _T_291; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:110:@7462.4]
  wire  _T_306; // @[NV_NVDLA_CDMA_IMG_sg.scala 223:75:@7477.6]
  wire  _T_309; // @[NV_NVDLA_CDMA_IMG_sg.scala 224:75:@7480.6]
  wire  _T_312; // @[NV_NVDLA_CDMA_IMG_sg.scala 225:65:@7482.6]
  wire  _T_315; // @[NV_NVDLA_CDMA_IMG_sg.scala 226:65:@7484.6]
  wire [13:0] _T_316; // @[NV_NVDLA_CDMA_IMG_sg.scala 227:57:@7485.6]
  wire [13:0] _T_317; // @[NV_NVDLA_CDMA_IMG_sg.scala 226:36:@7486.6]
  wire [13:0] _T_318; // @[NV_NVDLA_CDMA_IMG_sg.scala 225:36:@7487.6]
  wire [13:0] _T_319; // @[NV_NVDLA_CDMA_IMG_sg.scala 224:36:@7488.6]
  wire [13:0] _T_320; // @[NV_NVDLA_CDMA_IMG_sg.scala 223:36:@7489.6]
  wire [13:0] _GEN_13; // @[NV_NVDLA_CDMA_IMG_sg.scala 222:30:@7475.4]
  wire [2:0] _T_328; // @[NV_NVDLA_CDMA_IMG_sg.scala 232:50:@7497.6]
  wire [1:0] _T_329; // @[NV_NVDLA_CDMA_IMG_sg.scala 232:50:@7498.6]
  wire [1:0] _T_330; // @[NV_NVDLA_CDMA_IMG_sg.scala 231:34:@7499.6]
  wire [1:0] _T_331; // @[NV_NVDLA_CDMA_IMG_sg.scala 230:34:@7500.6]
  wire  _T_457; // @[NV_NVDLA_CDMA_IMG_sg.scala 297:83:@7611.4]
  wire  _T_458; // @[NV_NVDLA_CDMA_IMG_sg.scala 297:43:@7612.4]
  wire [1:0] _GEN_14; // @[NV_NVDLA_CDMA_IMG_sg.scala 229:28:@7492.4]
  wire [13:0] _GEN_65; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:50:@7520.4]
  wire  _T_357; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:50:@7520.4]
  wire  _T_359; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:103:@7521.4]
  wire  _T_360; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:81:@7522.4]
  wire  _T_361; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:50:@7523.4]
  wire  _T_364; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:84:@7525.4]
  wire  _T_365; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:117:@7526.4]
  wire  _T_366; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:115:@7527.4]
  wire  _T_367; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:113:@7528.4]
  wire  _T_381; // @[NV_NVDLA_CDMA_IMG_sg.scala 256:56:@7540.6]
  wire [5:0] _T_382; // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7541.6]
  wire [5:0] _T_383; // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7542.6]
  wire [4:0] _T_384; // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7543.6]
  wire [4:0] _T_385; // @[NV_NVDLA_CDMA_IMG_sg.scala 257:37:@7544.6]
  wire [4:0] _T_386; // @[NV_NVDLA_CDMA_IMG_sg.scala 256:37:@7545.6]
  wire  _T_388; // @[NV_NVDLA_CDMA_IMG_sg.scala 259:75:@7548.6]
  wire  _T_391; // @[NV_NVDLA_CDMA_IMG_sg.scala 260:75:@7551.6]
  wire  _T_394; // @[NV_NVDLA_CDMA_IMG_sg.scala 261:66:@7553.6]
  wire  _T_397; // @[NV_NVDLA_CDMA_IMG_sg.scala 262:66:@7555.6]
  wire [13:0] _T_398; // @[NV_NVDLA_CDMA_IMG_sg.scala 263:57:@7556.6]
  wire [13:0] _T_399; // @[NV_NVDLA_CDMA_IMG_sg.scala 262:36:@7557.6]
  wire [13:0] _T_400; // @[NV_NVDLA_CDMA_IMG_sg.scala 261:36:@7558.6]
  wire [13:0] _T_401; // @[NV_NVDLA_CDMA_IMG_sg.scala 260:36:@7559.6]
  wire [13:0] _T_402; // @[NV_NVDLA_CDMA_IMG_sg.scala 259:36:@7560.6]
  wire  _T_459; // @[NV_NVDLA_CDMA_IMG_sg.scala 298:63:@7614.4]
  wire  _T_460; // @[NV_NVDLA_CDMA_IMG_sg.scala 298:45:@7615.4]
  wire [4:0] _GEN_15; // @[NV_NVDLA_CDMA_IMG_sg.scala 255:30:@7539.4]
  wire [13:0] _GEN_16; // @[NV_NVDLA_CDMA_IMG_sg.scala 255:30:@7539.4]
  wire [2:0] _T_411; // @[NV_NVDLA_CDMA_IMG_sg.scala 268:50:@7569.6]
  wire [1:0] _T_412; // @[NV_NVDLA_CDMA_IMG_sg.scala 268:50:@7570.6]
  wire [1:0] _T_413; // @[NV_NVDLA_CDMA_IMG_sg.scala 267:34:@7571.6]
  wire [1:0] _T_414; // @[NV_NVDLA_CDMA_IMG_sg.scala 266:34:@7572.6]
  wire  _T_462; // @[NV_NVDLA_CDMA_IMG_sg.scala 299:82:@7618.4]
  wire  _T_463; // @[NV_NVDLA_CDMA_IMG_sg.scala 299:43:@7619.4]
  wire [1:0] _GEN_17; // @[NV_NVDLA_CDMA_IMG_sg.scala 265:28:@7563.4]
  wire  _T_416; // @[NV_NVDLA_CDMA_IMG_sg.scala 272:31:@7576.4]
  wire [4:0] _T_422; // @[NV_NVDLA_CDMA_IMG_sg.scala 275:33:@7582.4]
  wire  _T_424; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:49:@7584.4]
  wire  _T_425; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:66:@7585.4]
  wire  _T_426; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:27:@7586.4]
  wire  _T_439; // @[NV_NVDLA_CDMA_IMG_sg.scala 285:27:@7592.4]
  wire  _T_450; // @[NV_NVDLA_CDMA_IMG_sg.scala 293:39:@7601.4]
  wire  _T_451; // @[NV_NVDLA_CDMA_IMG_sg.scala 293:60:@7602.4]
  wire  _T_442; // @[NV_NVDLA_CDMA_IMG_sg.scala 287:38:@7593.4]
  wire  _T_444; // @[NV_NVDLA_CDMA_IMG_sg.scala 287:26:@7594.4]
  wire  _T_445; // @[NV_NVDLA_CDMA_IMG_sg.scala 286:26:@7595.4]
  wire  _T_446; // @[NV_NVDLA_CDMA_IMG_sg.scala 285:26:@7596.4]
  wire  _T_466; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:113:@7623.4]
  wire  _T_467; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:95:@7624.4]
  wire  _T_468; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:55:@7625.4]
  wire  _T_470; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:112:@7627.4]
  wire  _T_471; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:94:@7628.4]
  wire  _T_472; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:55:@7629.4]
  reg [31:0] _T_480; // @[NV_NVDLA_CDMA_IMG_sg.scala 306:41:@7637.4]
  reg [31:0] _RAND_23;
  reg [31:0] _T_483; // @[NV_NVDLA_CDMA_IMG_sg.scala 307:41:@7638.4]
  reg [31:0] _RAND_24;
  wire [32:0] _T_485; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:99:@7640.6]
  wire [31:0] _T_486; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:99:@7641.6]
  wire [31:0] _T_487; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:38:@7642.6]
  wire [31:0] _GEN_18; // @[NV_NVDLA_CDMA_IMG_sg.scala 309:24:@7639.4]
  wire  _T_488; // @[NV_NVDLA_CDMA_IMG_sg.scala 312:24:@7645.4]
  wire [32:0] _T_490; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:99:@7647.6]
  wire [31:0] _T_491; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:99:@7648.6]
  wire [31:0] _T_492; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:38:@7649.6]
  wire [31:0] _GEN_19; // @[NV_NVDLA_CDMA_IMG_sg.scala 312:41:@7646.4]
  reg [26:0] _T_495; // @[NV_NVDLA_CDMA_IMG_sg.scala 316:42:@7652.4]
  reg [31:0] _RAND_25;
  reg [26:0] _T_498; // @[NV_NVDLA_CDMA_IMG_sg.scala 317:42:@7653.4]
  reg [31:0] _RAND_26;
  wire [26:0] _GEN_66; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7656.6]
  wire [27:0] _T_501; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7656.6]
  wire [26:0] _T_502; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7657.6]
  wire [26:0] _T_503; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:39:@7658.6]
  wire [26:0] _GEN_20; // @[NV_NVDLA_CDMA_IMG_sg.scala 319:37:@7654.4]
  wire [26:0] _GEN_67; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7663.6]
  wire [27:0] _T_506; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7663.6]
  wire [26:0] _T_507; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7664.6]
  wire [26:0] _T_508; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:39:@7665.6]
  wire [26:0] _GEN_21; // @[NV_NVDLA_CDMA_IMG_sg.scala 322:37:@7661.4]
  reg [63:0] _T_510; // @[NV_NVDLA_CDMA_IMG_sg.scala 327:35:@7668.4]
  reg [63:0] _RAND_27;
  reg [63:0] _T_512; // @[NV_NVDLA_CDMA_IMG_sg.scala 328:35:@7669.4]
  reg [63:0] _RAND_28;
  wire [63:0] _GEN_68; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7670.4]
  wire [64:0] _T_513; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7670.4]
  wire [63:0] _T_514; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7671.4]
  wire [27:0] _T_516; // @[Cat.scala 30:58:@7672.4]
  wire [63:0] _GEN_69; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7673.4]
  wire [64:0] _T_517; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7673.4]
  wire [63:0] _T_518; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7674.4]
  wire [63:0] _GEN_70; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7675.4]
  wire [64:0] _T_519; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7675.4]
  wire [63:0] _T_520; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7676.4]
  wire [27:0] _T_522; // @[Cat.scala 30:58:@7677.4]
  wire [63:0] _GEN_71; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7678.4]
  wire [64:0] _T_523; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7678.4]
  wire [63:0] _T_524; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7679.4]
  wire [63:0] _T_525; // @[Cat.scala 30:58:@7681.6]
  wire [63:0] _T_526; // @[Cat.scala 30:58:@7683.6]
  reg [63:0] _T_529; // @[NV_NVDLA_CDMA_IMG_sg.scala 339:30:@7686.4]
  reg [63:0] _RAND_29;
  reg [4:0] _T_532; // @[NV_NVDLA_CDMA_IMG_sg.scala 340:30:@7687.4]
  reg [31:0] _RAND_30;
  reg [4:0] _T_535; // @[NV_NVDLA_CDMA_IMG_sg.scala 341:34:@7688.4]
  reg [31:0] _RAND_31;
  reg  _T_538; // @[NV_NVDLA_CDMA_IMG_sg.scala 342:33:@7689.4]
  reg [31:0] _RAND_32;
  reg  _T_541; // @[NV_NVDLA_CDMA_IMG_sg.scala 343:36:@7690.4]
  reg [31:0] _RAND_33;
  reg  _T_544; // @[NV_NVDLA_CDMA_IMG_sg.scala 344:34:@7691.4]
  reg [31:0] _RAND_34;
  reg  _T_547; // @[NV_NVDLA_CDMA_IMG_sg.scala 345:35:@7692.4]
  reg [31:0] _RAND_35;
  reg  _T_550; // @[NV_NVDLA_CDMA_IMG_sg.scala 346:29:@7693.4]
  reg [31:0] _RAND_36;
  reg  _T_553; // @[NV_NVDLA_CDMA_IMG_sg.scala 347:32:@7694.4]
  reg [31:0] _RAND_37;
  wire  _T_561; // @[NV_NVDLA_CDMA_IMG_sg.scala 352:29:@7697.4]
  wire  _T_562; // @[NV_NVDLA_CDMA_IMG_sg.scala 351:29:@7698.4]
  wire  _T_563; // @[NV_NVDLA_CDMA_IMG_sg.scala 350:29:@7699.4]
  wire [63:0] _T_564; // @[NV_NVDLA_CDMA_IMG_sg.scala 353:23:@7700.4]
  wire [5:0] _T_566; // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7701.4]
  wire [5:0] _T_567; // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7702.4]
  wire [4:0] _T_568; // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7703.4]
  wire  _T_569; // @[NV_NVDLA_CDMA_IMG_sg.scala 357:45:@7704.4]
  wire [63:0] _GEN_24; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire [4:0] _GEN_26; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_27; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_28; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_29; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_30; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_31; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_32; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  wire  _GEN_33; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  reg  _T_581; // @[NV_NVDLA_CDMA_IMG_sg.scala 382:30:@7723.4]
  reg [31:0] _RAND_38;
  wire  _T_586; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:43:@7728.4]
  wire  _T_587; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:58:@7729.4]
  wire  _T_589; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:28:@7730.4]
  wire  _T_590; // @[NV_NVDLA_CDMA_IMG_sg.scala 385:28:@7731.4]
  reg  _T_593; // @[NV_NVDLA_CDMA_IMG_sg.scala 392:34:@7733.4]
  reg [31:0] _RAND_39;
  wire  _T_594; // @[NV_NVDLA_CDMA_IMG_sg.scala 394:49:@7734.4]
  wire [14:0] _T_596; // @[NV_NVDLA_CDMA_IMG_sg.scala 396:33:@7735.4]
  wire [14:0] _T_597; // @[NV_NVDLA_CDMA_IMG_sg.scala 395:33:@7736.4]
  wire [14:0] _T_598; // @[NV_NVDLA_CDMA_IMG_sg.scala 394:33:@7737.4]
  wire [14:0] _GEN_72; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7738.4]
  wire [15:0] _T_599; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7738.4]
  wire [14:0] _T_600; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7739.4]
  wire  _T_601; // @[NV_NVDLA_CDMA_IMG_sg.scala 399:53:@7740.4]
  wire  _T_603; // @[NV_NVDLA_CDMA_IMG_sg.scala 400:46:@7742.4]
  wire  _T_606; // @[NV_NVDLA_CDMA_IMG_sg.scala 401:59:@7744.4]
  wire  _T_608; // @[NV_NVDLA_CDMA_IMG_sg.scala 402:31:@7745.4]
  wire  _T_609; // @[NV_NVDLA_CDMA_IMG_sg.scala 402:30:@7746.4]
  wire  _T_610; // @[NV_NVDLA_CDMA_IMG_sg.scala 401:30:@7747.4]
  wire  _T_611; // @[NV_NVDLA_CDMA_IMG_sg.scala 400:30:@7748.4]
  wire [14:0] _T_613; // @[NV_NVDLA_CDMA_IMG_sg.scala 404:34:@7749.4]
  wire  _T_614; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:35:@7750.4]
  wire  _T_615; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:48:@7751.4]
  wire  _T_617; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:65:@7753.4]
  wire [14:0] _T_619; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:34:@7754.4]
  wire [15:0] _T_620; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:45:@7755.4]
  wire [14:0] _T_621; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:45:@7756.4]
  wire [15:0] _T_622; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7757.4]
  wire [15:0] _T_623; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7758.4]
  wire [14:0] _T_624; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7759.4]
  wire  _T_629; // @[NV_NVDLA_CDMA_IMG_sg.scala 407:79:@7764.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CDMA_IMG_sg.scala 410:29:@7766.4]
  wire [14:0] _T_641; // @[NV_NVDLA_CDMA_IMG_sg.scala 452:31:@7801.4 NV_NVDLA_CDMA_IMG_sg.scala 459:21:@7814.4]
  wire  _T_650; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:36:@7808.4]
  wire  _T_651; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:57:@7809.4]
  wire  _T_652; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:75:@7810.4]
  wire  _T_653; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:73:@7811.4]
  wire  _T_682; // @[NV_NVDLA_CDMA_IMG_sg.scala 498:42:@7850.4]
  wire  _T_684; // @[NV_NVDLA_CDMA_IMG_sg.scala 501:43:@7852.4]
  wire  _T_661; // @[NV_NVDLA_CDMA_IMG_sg.scala 480:38:@7830.4]
  wire [6:0] _T_665; // @[Cat.scala 30:58:@7835.4]
  wire [3:0] _T_668; // @[Cat.scala 30:58:@7838.4]
  wire [256:0] _T_635; // @[NV_NVDLA_CDMA_IMG_sg.scala 422:29:@7771.4 NV_NVDLA_CDMA_IMG_sg.scala 445:19:@7798.4]
  wire [255:0] _T_670; // @[NV_NVDLA_CDMA_IMG_sg.scala 488:40:@7841.4]
  wire  _T_671; // @[NV_NVDLA_CDMA_IMG_sg.scala 489:40:@7842.4]
  reg [4:0] _T_674; // @[NV_NVDLA_CDMA_IMG_sg.scala 490:35:@7843.4]
  reg [31:0] _RAND_40;
  wire  _T_677; // @[NV_NVDLA_CDMA_IMG_sg.scala 493:43:@7845.4]
  wire  _T_678; // @[NV_NVDLA_CDMA_IMG_sg.scala 494:40:@7846.4]
  wire  _T_679; // @[NV_NVDLA_CDMA_IMG_sg.scala 495:45:@7847.4]
  wire  _T_681; // @[NV_NVDLA_CDMA_IMG_sg.scala 497:44:@7849.4]
  wire [4:0] _T_683; // @[NV_NVDLA_CDMA_IMG_sg.scala 499:41:@7851.4]
  wire  _T_685; // @[NV_NVDLA_CDMA_IMG_sg.scala 503:28:@7854.4]
  wire  _T_687; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:27:@7855.4]
  wire  _T_637; // @[NV_NVDLA_CDMA_IMG_sg.scala 423:30:@7772.4 NV_NVDLA_CDMA_IMG_sg.scala 446:20:@7799.4]
  wire  _T_689; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:58:@7857.4]
  wire  _T_691; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:26:@7858.4]
  wire  _T_692; // @[NV_NVDLA_CDMA_IMG_sg.scala 503:27:@7859.4]
  wire [4:0] _GEN_74; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7860.4]
  wire [5:0] _T_693; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7860.4]
  wire [4:0] _T_694; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7861.4]
  wire  _T_695; // @[NV_NVDLA_CDMA_IMG_sg.scala 508:55:@7862.4]
  wire [4:0] _T_697; // @[NV_NVDLA_CDMA_IMG_sg.scala 508:33:@7863.4]
  wire  _T_698; // @[NV_NVDLA_CDMA_IMG_sg.scala 513:54:@7867.4]
  wire  _T_699; // @[NV_NVDLA_CDMA_IMG_sg.scala 513:37:@7868.4]
  wire [4:0] _GEN_35; // @[NV_NVDLA_CDMA_IMG_sg.scala 510:22:@7864.4]
  wire  _T_701; // @[NV_NVDLA_CDMA_IMG_sg.scala 514:40:@7871.4]
  reg  _T_710; // @[NV_NVDLA_CDMA_IMG_sg.scala 523:33:@7876.4]
  reg [31:0] _RAND_41;
  reg [255:0] _T_712; // @[NV_NVDLA_CDMA_IMG_sg.scala 524:30:@7877.4]
  reg [255:0] _RAND_42;
  wire  _T_713; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:41:@7882.4]
  wire  _T_714; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:45:@7883.4]
  wire  _T_715; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:76:@7884.4]
  wire  _T_716; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:79:@7885.4]
  wire [7:0] _T_717; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:110:@7886.4]
  wire  _T_718; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:39:@7887.4]
  wire  _T_719; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:44:@7888.4]
  wire  _T_720; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:60:@7889.4]
  wire  _T_721; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:42:@7890.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@7893.4]
  wire  _T_1041; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:67:@8190.4]
  wire [255:0] _T_1045; // @[Bitwise.scala 72:12:@8192.4]
  wire [255:0] _T_1046; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:72:@8193.4]
  wire  _T_1047; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:66:@8194.4]
  wire [255:0] _T_1051; // @[Bitwise.scala 72:12:@8196.4]
  wire [7:0] _T_774; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7943.4]
  wire [7:0] _T_775; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7944.4]
  wire [7:0] _T_776; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7945.4]
  wire [7:0] _T_777; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7946.4]
  wire [7:0] _T_767; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7936.4]
  wire [7:0] _T_768; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7937.4]
  wire [7:0] _T_769; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7938.4]
  wire [7:0] _T_770; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7939.4]
  wire [7:0] _T_760; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7929.4]
  wire [7:0] _T_761; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7930.4]
  wire [7:0] _T_762; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7931.4]
  wire [7:0] _T_763; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7932.4]
  wire [7:0] _T_753; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7922.4]
  wire [7:0] _T_754; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7923.4]
  wire [7:0] _T_755; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7924.4]
  wire [7:0] _T_756; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7925.4]
  wire [63:0] _T_798; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7962.4]
  wire [7:0] _T_746; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7915.4]
  wire [7:0] _T_747; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7916.4]
  wire [7:0] _T_748; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7917.4]
  wire [7:0] _T_749; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7918.4]
  wire [7:0] _T_739; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7908.4]
  wire [7:0] _T_740; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7909.4]
  wire [7:0] _T_741; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7910.4]
  wire [7:0] _T_742; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7911.4]
  wire [7:0] _T_732; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7901.4]
  wire [7:0] _T_733; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7902.4]
  wire [7:0] _T_734; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7903.4]
  wire [7:0] _T_735; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7904.4]
  wire [7:0] _T_725; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7894.4]
  wire [7:0] _T_726; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7895.4]
  wire [7:0] _T_727; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7896.4]
  wire [7:0] _T_728; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7897.4]
  wire [63:0] _T_795; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7959.4]
  wire [127:0] _T_797; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7961.4]
  wire [255:0] _T_801; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7965.4]
  wire [255:0] _T_1052; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:71:@8197.4]
  wire [255:0] _T_1053; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:94:@8198.4]
  wire  _T_1054; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:66:@8199.4]
  wire [255:0] _T_1058; // @[Bitwise.scala 72:12:@8201.4]
  wire [63:0] _T_875; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8034.4]
  wire [63:0] _T_872; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8031.4]
  wire [127:0] _T_874; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8033.4]
  wire [255:0] _T_878; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8037.4]
  wire [255:0] _T_1059; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:71:@8202.4]
  wire [255:0] _T_1060; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:93:@8203.4]
  wire  _T_1061; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:66:@8204.4]
  wire [255:0] _T_1065; // @[Bitwise.scala 72:12:@8206.4]
  wire [63:0] _T_952; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8106.4]
  wire [63:0] _T_949; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8103.4]
  wire [127:0] _T_951; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8105.4]
  wire [255:0] _T_955; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8109.4]
  wire [255:0] _T_1066; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:71:@8207.4]
  wire [255:0] _T_1067; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:93:@8208.4]
  wire  _T_1068; // @[NV_NVDLA_CDMA_IMG_sg.scala 563:66:@8209.4]
  wire [255:0] _T_1072; // @[Bitwise.scala 72:12:@8211.4]
  wire [63:0] _T_1035; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8184.4]
  wire [63:0] _T_1028; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8177.4]
  wire [127:0] _T_1032; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8181.4]
  wire [255:0] _T_1040; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8189.4]
  wire [255:0] _T_1073; // @[NV_NVDLA_CDMA_IMG_sg.scala 563:71:@8212.4]
  wire [255:0] _T_1074; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:93:@8213.4]
  wire  _T_1076; // @[NV_NVDLA_CDMA_IMG_sg.scala 566:67:@8215.4]
  wire  _T_1077; // @[NV_NVDLA_CDMA_IMG_sg.scala 566:47:@8216.4]
  reg  _T_1080; // @[NV_NVDLA_CDMA_IMG_sg.scala 568:33:@8217.4]
  reg [31:0] _RAND_43;
  reg  _T_1083; // @[NV_NVDLA_CDMA_IMG_sg.scala 569:36:@8218.4]
  reg [31:0] _RAND_44;
  reg  _T_1086; // @[NV_NVDLA_CDMA_IMG_sg.scala 570:34:@8219.4]
  reg [31:0] _RAND_45;
  wire  _GEN_37; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  wire  _GEN_38; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  wire  _GEN_39; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  reg [4:0] _T_1092; // @[NV_NVDLA_CDMA_IMG_sg.scala 579:39:@8227.4]
  reg [31:0] _RAND_46;
  reg  _T_1095; // @[NV_NVDLA_CDMA_IMG_sg.scala 580:35:@8228.4]
  reg [31:0] _RAND_47;
  reg  _T_1101; // @[NV_NVDLA_CDMA_IMG_sg.scala 582:30:@8230.4]
  reg [31:0] _RAND_48;
  wire  _T_1102; // @[NV_NVDLA_CDMA_IMG_sg.scala 583:24:@8231.4]
  wire [4:0] _GEN_40; // @[NV_NVDLA_CDMA_IMG_sg.scala 583:45:@8232.4]
  wire  _T_1103; // @[NV_NVDLA_CDMA_IMG_sg.scala 587:46:@8236.6]
  wire  _T_1105; // @[NV_NVDLA_CDMA_IMG_sg.scala 589:36:@8240.6]
  wire  _GEN_41; // @[NV_NVDLA_CDMA_IMG_sg.scala 586:24:@8235.4]
  wire  _GEN_43; // @[NV_NVDLA_CDMA_IMG_sg.scala 586:24:@8235.4]
  wire  _T_1106; // @[NV_NVDLA_CDMA_IMG_sg.scala 596:49:@8243.4]
  wire  _T_1107; // @[NV_NVDLA_CDMA_IMG_sg.scala 596:46:@8244.4]
  wire  _T_1108; // @[NV_NVDLA_CDMA_IMG_sg.scala 597:46:@8245.4]
  reg [255:0] _T_1111; // @[NV_NVDLA_CDMA_IMG_sg.scala 600:40:@8246.4]
  reg [255:0] _RAND_49;
  reg [255:0] _T_1114; // @[NV_NVDLA_CDMA_IMG_sg.scala 601:40:@8247.4]
  reg [255:0] _RAND_50;
  wire [255:0] _GEN_44; // @[NV_NVDLA_CDMA_IMG_sg.scala 603:29:@8248.4]
  wire [255:0] _GEN_45; // @[NV_NVDLA_CDMA_IMG_sg.scala 606:29:@8251.4]
  reg  _T_1117; // @[NV_NVDLA_CDMA_IMG_sg.scala 611:36:@8254.4]
  reg [31:0] _RAND_51;
  reg [255:0] _T_1119; // @[NV_NVDLA_CDMA_IMG_sg.scala 612:33:@8255.4]
  reg [255:0] _RAND_52;
  wire  _T_1122; // @[NV_NVDLA_CDMA_IMG_sg.scala 615:49:@8257.4]
  wire  _T_1123; // @[NV_NVDLA_CDMA_IMG_sg.scala 615:46:@8258.4]
  wire [255:0] _T_1124; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:62:@8259.4]
  wire [4:0] _T_1131; // @[NV_NVDLA_CDMA_IMG_sg.scala 624:23:@8268.4]
  wire [7:0] _T_1126; // @[Cat.scala 30:58:@8260.4]
  wire [255:0] _T_1127; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:128:@8261.4]
  wire [511:0] _T_1128; // @[Cat.scala 30:58:@8262.4]
  wire [255:0] _T_1129; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:165:@8263.4]
  reg [6:0] _T_1134; // @[NV_NVDLA_CDMA_IMG_sg.scala 627:41:@8270.4]
  reg [31:0] _RAND_53;
  reg [6:0] _T_1137; // @[NV_NVDLA_CDMA_IMG_sg.scala 628:41:@8271.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_1140; // @[NV_NVDLA_CDMA_IMG_sg.scala 629:37:@8272.4]
  reg [31:0] _RAND_55;
  wire [7:0] _T_1141; // @[NV_NVDLA_CDMA_IMG_sg.scala 631:61:@8273.4]
  wire [6:0] _T_1142; // @[NV_NVDLA_CDMA_IMG_sg.scala 631:61:@8274.4]
  wire [7:0] _T_1143; // @[NV_NVDLA_CDMA_IMG_sg.scala 632:61:@8275.4]
  wire [6:0] _T_1144; // @[NV_NVDLA_CDMA_IMG_sg.scala 632:61:@8276.4]
  wire [6:0] _T_1146; // @[NV_NVDLA_CDMA_IMG_sg.scala 633:39:@8277.4]
  wire [6:0] _T_1148; // @[NV_NVDLA_CDMA_IMG_sg.scala 634:39:@8278.4]
  wire  _T_1150; // @[NV_NVDLA_CDMA_IMG_sg.scala 635:73:@8280.4]
  wire  _T_1151; // @[NV_NVDLA_CDMA_IMG_sg.scala 635:50:@8281.4]
  wire  _T_1152; // @[NV_NVDLA_CDMA_IMG_sg.scala 636:73:@8282.4]
  wire  _T_1153; // @[NV_NVDLA_CDMA_IMG_sg.scala 636:50:@8283.4]
  wire  _T_1156; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:83:@8285.4]
  wire [5:0] _T_1157; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:110:@8286.4]
  wire [7:0] _T_1159; // @[Cat.scala 30:58:@8288.4]
  wire  _T_1161; // @[NV_NVDLA_CDMA_IMG_sg.scala 638:60:@8289.4]
  wire [5:0] _T_1162; // @[NV_NVDLA_CDMA_IMG_sg.scala 638:87:@8290.4]
  wire [7:0] _T_1164; // @[Cat.scala 30:58:@8292.4]
  wire [7:0] _T_1165; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:30:@8293.4]
  wire [6:0] _GEN_47; // @[NV_NVDLA_CDMA_IMG_sg.scala 640:32:@8294.4]
  wire [6:0] _GEN_48; // @[NV_NVDLA_CDMA_IMG_sg.scala 643:32:@8297.4]
  wire [7:0] _GEN_49; // @[NV_NVDLA_CDMA_IMG_sg.scala 646:30:@8300.4]
  reg [3:0] _T_1168; // @[NV_NVDLA_CDMA_IMG_sg.scala 651:39:@8303.4]
  reg [31:0] _RAND_56;
  reg [4:0] _T_1171; // @[NV_NVDLA_CDMA_IMG_sg.scala 652:39:@8304.4]
  reg [31:0] _RAND_57;
  reg [3:0] _T_1174; // @[NV_NVDLA_CDMA_IMG_sg.scala 653:43:@8305.4]
  reg [31:0] _RAND_58;
  reg [4:0] _T_1177; // @[NV_NVDLA_CDMA_IMG_sg.scala 654:43:@8306.4]
  reg [31:0] _RAND_59;
  wire [3:0] _T_1187; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:79:@8310.4]
  wire [4:0] _T_1188; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:57:@8311.4]
  wire [3:0] _T_1189; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:57:@8312.4]
  wire [3:0] _GEN_75; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8313.4]
  wire [4:0] _T_1190; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8313.4]
  wire [4:0] _T_1191; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8314.4]
  wire [3:0] _T_1192; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8315.4]
  wire [5:0] _T_1193; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:57:@8316.4]
  wire [4:0] _T_1194; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:57:@8317.4]
  wire [4:0] _GEN_76; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8318.4]
  wire [5:0] _T_1195; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8318.4]
  wire [5:0] _T_1196; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8319.4]
  wire [4:0] _T_1197; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8320.4]
  wire [3:0] _T_1202; // @[NV_NVDLA_CDMA_IMG_sg.scala 663:37:@8323.4]
  wire [3:0] _T_1204; // @[NV_NVDLA_CDMA_IMG_sg.scala 661:37:@8325.4]
  wire [4:0] _T_1208; // @[NV_NVDLA_CDMA_IMG_sg.scala 667:37:@8327.4]
  wire [4:0] _T_1210; // @[NV_NVDLA_CDMA_IMG_sg.scala 665:37:@8329.4]
  wire [3:0] _GEN_50; // @[NV_NVDLA_CDMA_IMG_sg.scala 677:34:@8343.4]
  wire [4:0] _GEN_51; // @[NV_NVDLA_CDMA_IMG_sg.scala 680:34:@8346.4]
  wire [3:0] _GEN_52; // @[NV_NVDLA_CDMA_IMG_sg.scala 683:35:@8349.4]
  wire [4:0] _GEN_53; // @[NV_NVDLA_CDMA_IMG_sg.scala 686:35:@8352.4]
  reg  _T_1226; // @[NV_NVDLA_CDMA_IMG_sg.scala 695:34:@8360.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[NV_NVDLA_CDMA_IMG_sg.scala 698:45:@8361.4]
  wire  _T_1230; // @[NV_NVDLA_CDMA_IMG_sg.scala 698:32:@8362.4]
  wire  _T_1231; // @[NV_NVDLA_CDMA_IMG_sg.scala 697:32:@8363.4]
  wire  _GEN_56; // @[NV_NVDLA_CDMA_IMG_sg.scala 700:24:@8364.4]
  wire [8:0] _T_1234; // @[Cat.scala 30:58:@8372.4]
  reg  _T_1243; // @[NV_NVDLA_CDMA_IMG_sg.scala 756:33:@8398.4]
  reg [31:0] _RAND_61;
  wire  _T_1244; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:24:@8399.4]
  wire  _T_1245; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:42:@8400.4]
  wire  _T_1246; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:56:@8401.4]
  wire  _GEN_57; // @[NV_NVDLA_CDMA_IMG_sg.scala 760:24:@8402.4]
  wire  _T_1247; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:53:@8406.4]
  wire  _T_1248; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:51:@8407.4]
  wire  _T_1249; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:69:@8408.4]
  reg  _T_1252; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:35:@8409.4]
  reg [31:0] _RAND_62;
  wire  _T_1253; // @[NV_NVDLA_CDMA_IMG_sg.scala 770:61:@8411.4]
  reg  _T_1256; // @[NV_NVDLA_CDMA_IMG_sg.scala 770:35:@8412.4]
  reg [31:0] _RAND_63;
  wire  _T_1257; // @[NV_NVDLA_CDMA_IMG_sg.scala 771:52:@8414.4]
  reg  _T_1260; // @[NV_NVDLA_CDMA_IMG_sg.scala 771:35:@8415.4]
  reg [31:0] _RAND_64;
  reg  _T_1267; // @[NV_NVDLA_CDMA_IMG_sg.scala 784:37:@8429.4]
  reg [31:0] _RAND_65;
  wire  _T_1269; // @[NV_NVDLA_CDMA_IMG_sg.scala 785:57:@8432.4]
  wire  _T_1270; // @[NV_NVDLA_CDMA_IMG_sg.scala 785:74:@8433.4]
  reg  _T_1273; // @[NV_NVDLA_CDMA_IMG_sg.scala 785:37:@8434.4]
  reg [31:0] _RAND_66;
  reg  _T_1276; // @[NV_NVDLA_CDMA_IMG_sg.scala 786:37:@8436.4]
  reg [31:0] _RAND_67;
  reg  _T_1280; // @[NV_NVDLA_CDMA_IMG_sg.scala 787:37:@8439.4]
  reg [31:0] _RAND_68;
  wire [8:0] _T_1282; // @[NV_NVDLA_CDMA_IMG_sg.scala 789:42:@8441.4 NV_NVDLA_CDMA_IMG_sg.scala 799:32:@8454.4]
  wire  _T_1284; // @[NV_NVDLA_CDMA_IMG_sg.scala 790:49:@8442.4]
  wire [31:0] _T_1289; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:48:@8455.4]
  wire  _T_1291; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:48:@8456.4]
  wire  _T_1292; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:22:@8457.4]
  wire  _T_1294; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:84:@8458.4]
  NV_soDLA_DMAIF_rdreq NV_soDLA_DMAIF_rdreq ( // @[NV_NVDLA_CDMA_IMG_sg.scala 426:41:@7774.4]
    .reset(NV_NVDLA_DMAIF_rdreq_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk),
    .io_dmaif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready),
    .io_dmaif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid),
    .io_dmaif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits),
    .io_mcif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready),
    .io_mcif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid),
    .io_mcif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits),
    .io_cvif_rd_req_pd_ready(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready),
    .io_cvif_rd_req_pd_valid(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid),
    .io_cvif_rd_req_pd_bits(NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits),
    .io_reg2dp_src_ram_type(NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type)
  );
  NV_soDLA_DMAIF_rdrsp NV_soDLA_DMAIF_rdrsp ( // @[NV_NVDLA_CDMA_IMG_sg.scala 438:41:@7788.4]
    .reset(NV_NVDLA_DMAIF_rdrsp_reset),
    .io_nvdla_core_clk(NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk),
    .io_mcif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready),
    .io_mcif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid),
    .io_mcif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits),
    .io_cvif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready),
    .io_cvif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid),
    .io_cvif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits),
    .io_dmaif_rd_rsp_pd_ready(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready),
    .io_dmaif_rd_rsp_pd_valid(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid),
    .io_dmaif_rd_rsp_pd_bits(NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits)
  );
  NV_NVDLA_fifo_3 NV_NVDLA_fifo ( // @[NV_NVDLA_CDMA_IMG_sg.scala 467:42:@7821.4]
    .clock(NV_NVDLA_fifo_clock),
    .reset(NV_NVDLA_fifo_reset),
    .io_clk(NV_NVDLA_fifo_io_clk),
    .io_wr_pvld(NV_NVDLA_fifo_io_wr_pvld),
    .io_wr_prdy(NV_NVDLA_fifo_io_wr_prdy),
    .io_wr_pd(NV_NVDLA_fifo_io_wr_pd),
    .io_rd_pvld(NV_NVDLA_fifo_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_io_rd_pd)
  );
  NV_NVDLA_fifo_4 NV_NVDLA_fifo_1 ( // @[NV_NVDLA_CDMA_IMG_sg.scala 729:50:@8379.4]
    .clock(NV_NVDLA_fifo_1_clock),
    .reset(NV_NVDLA_fifo_1_reset),
    .io_wr_pd(NV_NVDLA_fifo_1_io_wr_pd),
    .io_rd_pvld(NV_NVDLA_fifo_1_io_rd_pvld),
    .io_rd_prdy(NV_NVDLA_fifo_1_io_rd_prdy),
    .io_rd_pd(NV_NVDLA_fifo_1_io_rd_pd)
  );
  NV_COUNTER_STAGE_histogram NV_COUNTER_STAGE_histogram ( // @[NV_NVDLA_CDMA_IMG_sg.scala 775:21:@8417.4]
    .reset(NV_COUNTER_STAGE_histogram_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_io_rd_stall_inc),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_io_cnt_cur)
  );
  NV_COUNTER_STAGE_histogram_1 NV_COUNTER_STAGE_histogram_1 ( // @[NV_NVDLA_CDMA_IMG_sg.scala 793:23:@8446.4]
    .reset(NV_COUNTER_STAGE_histogram_1_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_1_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc),
    .io_rd_stall_dec(NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_1_io_cnt_cur)
  );
  NV_COUNTER_STAGE_histogram NV_COUNTER_STAGE_histogram_2 ( // @[NV_NVDLA_CDMA_IMG_sg.scala 805:23:@8460.4]
    .reset(NV_COUNTER_STAGE_histogram_2_reset),
    .io_clk(NV_COUNTER_STAGE_histogram_2_io_clk),
    .io_rd_stall_inc(NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc),
    .io_rd_stall_clr(NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr),
    .io_rd_stall_cen(NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen),
    .io_cnt_cur(NV_COUNTER_STAGE_histogram_2_io_cnt_cur)
  );
  assign _T_170 = ~ _T_157; // @[NV_NVDLA_CDMA_IMG_sg.scala 126:44:@7362.4]
  assign _T_171 = io_is_running & _T_170; // @[NV_NVDLA_CDMA_IMG_sg.scala 126:42:@7363.4]
  assign _T_175 = io_reg2dp_datain_height + 13'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 131:48:@7368.6]
  assign _T_177 = io_reg2dp_entries + 14'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 133:43:@7371.6]
  assign _GEN_0 = io_layer_st ? io_reg2dp_mean_format : _T_160; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  assign _GEN_1 = io_layer_st ? _T_175 : _T_163; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  assign _GEN_2 = io_layer_st ? io_reg2dp_datain_height : _T_166; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  assign _GEN_3 = io_layer_st ? _T_177 : _T_169; // @[NV_NVDLA_CDMA_IMG_sg.scala 129:22:@7365.4]
  assign _T_199 = _T_163[13:4]; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:38:@7380.4]
  assign _T_201 = _T_199 != 10'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:46:@7381.4]
  assign _T_202 = ~ _T_201; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:25:@7382.4]
  assign _T_203 = _T_163[3:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:67:@7383.4]
  assign _T_204 = _T_203 <= 4'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:74:@7384.4]
  assign _T_205 = _T_202 & _T_204; // @[NV_NVDLA_CDMA_IMG_sg.scala 150:52:@7385.4]
  assign _T_214 = _T_205 ? _T_203 : 4'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 153:25:@7393.4]
  assign _GEN_58 = {{11'd0}, _T_214}; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:38:@7396.4]
  assign _T_217 = _GEN_58 * _T_169; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:38:@7396.4]
  assign _T_218 = _T_217[14:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 155:53:@7397.4]
  assign _GEN_4 = _T_171 ? _T_214 : _T_180; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _GEN_5 = _T_171 ? 4'h1 : _T_183; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _GEN_6 = _T_171 ? _T_214 : _T_186; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _GEN_7 = _T_171 ? _T_218 : _T_189; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _GEN_8 = _T_171 ? _T_169 : _T_192; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _GEN_9 = _T_171 ? _T_218 : _T_195; // @[NV_NVDLA_CDMA_IMG_sg.scala 158:27:@7400.4]
  assign _T_230 = _T_226 != 13'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 177:42:@7410.4]
  assign _T_231 = ~ _T_230; // @[NV_NVDLA_CDMA_IMG_sg.scala 177:25:@7411.4]
  assign _T_232 = _T_226 == _T_166; // @[NV_NVDLA_CDMA_IMG_sg.scala 178:42:@7412.4]
  assign _T_235 = _T_226 + 13'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:83:@7414.6]
  assign _T_236 = _T_226 + 13'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:83:@7415.6]
  assign _T_237 = _T_171 ? 13'h0 : _T_236; // @[NV_NVDLA_CDMA_IMG_sg.scala 181:30:@7416.6]
  assign _T_447 = ~ _T_436; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:32:@7598.4]
  assign _T_573 = NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 379:30:@7720.4 NV_NVDLA_CDMA_IMG_sg.scala 436:20:@7787.4]
  assign _T_582 = _T_573 | _T_556; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:38:@7724.4]
  assign _T_575 = NV_NVDLA_fifo_io_wr_prdy; // @[NV_NVDLA_CDMA_IMG_sg.scala 380:34:@7721.4 NV_NVDLA_CDMA_IMG_sg.scala 473:24:@7827.4]
  assign _T_583 = _T_582 & _T_575; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:57:@7725.4]
  assign _T_584 = _T_583 & _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 384:78:@7726.4]
  assign _T_448 = _T_447 | _T_584; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:46:@7599.4]
  assign _T_449 = _T_433 & _T_448; // @[NV_NVDLA_CDMA_IMG_sg.scala 292:29:@7600.4]
  assign _T_417 = ~ _T_240; // @[NV_NVDLA_CDMA_IMG_sg.scala 273:33:@7577.4]
  assign _GEN_60 = {{10'd0}, _T_250}; // @[NV_NVDLA_CDMA_IMG_sg.scala 213:48:@7452.4]
  assign _T_280 = _T_267 <= _GEN_60; // @[NV_NVDLA_CDMA_IMG_sg.scala 213:48:@7452.4]
  assign _T_293 = _T_270 == 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:66:@7463.4]
  assign _T_294 = _T_280 & _T_293; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:44:@7464.4]
  assign _T_295 = ~ io_pixel_planar0_rp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:77:@7465.4]
  assign _T_296 = _T_294 & _T_295; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:75:@7466.4]
  assign _T_298 = _T_270 == 2'h2; // @[NV_NVDLA_CDMA_IMG_sg.scala 217:69:@7467.4]
  assign _T_299 = _T_280 & _T_298; // @[NV_NVDLA_CDMA_IMG_sg.scala 217:47:@7468.4]
  assign _T_300 = _T_296 | _T_299; // @[NV_NVDLA_CDMA_IMG_sg.scala 216:102:@7469.4]
  assign _GEN_61 = {{9'd0}, _T_334}; // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7510.4]
  assign _T_349 = _T_337 - _GEN_61; // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7510.4]
  assign _T_350 = $unsigned(_T_349); // @[NV_NVDLA_CDMA_IMG_sg.scala 244:57:@7511.4]
  assign _T_354 = _T_350[14]; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:50:@7516.4]
  assign _T_355 = _T_337 == _GEN_61; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:79:@7517.4]
  assign _T_356 = _T_354 | _T_355; // @[NV_NVDLA_CDMA_IMG_sg.scala 247:55:@7518.4]
  assign _T_369 = _T_340 == 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:69:@7529.4]
  assign _T_370 = _T_356 & _T_369; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:47:@7530.4]
  assign _T_371 = ~ io_pixel_planar1_rp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:80:@7531.4]
  assign _T_372 = _T_370 & _T_371; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:78:@7532.4]
  assign _T_374 = _T_340 == 2'h2; // @[NV_NVDLA_CDMA_IMG_sg.scala 251:69:@7533.4]
  assign _T_375 = _T_356 & _T_374; // @[NV_NVDLA_CDMA_IMG_sg.scala 251:47:@7534.4]
  assign _T_376 = _T_372 | _T_375; // @[NV_NVDLA_CDMA_IMG_sg.scala 250:106:@7535.4]
  assign _T_418 = _T_417 ? _T_300 : _T_376; // @[NV_NVDLA_CDMA_IMG_sg.scala 273:32:@7578.4]
  assign _T_475 = _T_449 & _T_418; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:57:@7633.4]
  assign _T_243 = _T_240 == io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_sg.scala 186:50:@7421.4]
  assign _T_476 = _T_475 & _T_243; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:77:@7634.4]
  assign _T_477 = _T_171 | _T_476; // @[NV_NVDLA_CDMA_IMG_sg.scala 303:39:@7635.4]
  assign _GEN_10 = _T_477 ? _T_237 : _T_226; // @[NV_NVDLA_CDMA_IMG_sg.scala 180:24:@7413.4]
  assign _T_244 = _T_171 | _T_243; // @[NV_NVDLA_CDMA_IMG_sg.scala 187:54:@7422.4]
  assign _T_247 = _T_244 ? 1'h0 : _T_417; // @[NV_NVDLA_CDMA_IMG_sg.scala 187:35:@7424.4]
  assign _T_275 = _T_267 - _GEN_60; // @[NV_NVDLA_CDMA_IMG_sg.scala 211:57:@7446.4]
  assign _T_276 = $unsigned(_T_275); // @[NV_NVDLA_CDMA_IMG_sg.scala 211:57:@7447.4]
  assign _T_277 = _T_276[14]; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:57:@7448.4]
  assign _T_278 = _T_267[3:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:83:@7449.4]
  assign _T_279 = _T_277 ? _T_278 : _T_250; // @[NV_NVDLA_CDMA_IMG_sg.scala 212:32:@7450.4]
  assign _T_301 = _T_279 == _T_250; // @[NV_NVDLA_CDMA_IMG_sg.scala 218:47:@7471.4]
  assign _T_302 = _T_301 | _T_300; // @[NV_NVDLA_CDMA_IMG_sg.scala 218:74:@7472.4]
  assign _T_352 = _T_337[4:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 245:83:@7513.4]
  assign _T_353 = _T_354 ? _T_352 : _T_334; // @[NV_NVDLA_CDMA_IMG_sg.scala 245:32:@7514.4]
  assign _T_377 = _T_353 == _T_334; // @[NV_NVDLA_CDMA_IMG_sg.scala 252:50:@7536.4]
  assign _T_378 = _T_377 | _T_376; // @[NV_NVDLA_CDMA_IMG_sg.scala 252:77:@7537.4]
  assign _T_420 = _T_417 ? _T_302 : _T_378; // @[NV_NVDLA_CDMA_IMG_sg.scala 274:32:@7580.4]
  assign _T_473 = _T_449 & _T_420; // @[NV_NVDLA_CDMA_IMG_sg.scala 302:61:@7630.4]
  assign _T_474 = _T_171 | _T_473; // @[NV_NVDLA_CDMA_IMG_sg.scala 302:43:@7631.4]
  assign _GEN_11 = _T_474 ? _T_247 : _T_240; // @[NV_NVDLA_CDMA_IMG_sg.scala 189:28:@7425.4]
  assign _T_259 = _T_171 | _T_300; // @[NV_NVDLA_CDMA_IMG_sg.scala 200:55:@7434.6]
  assign _T_260 = _T_250 - _T_279; // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7435.6]
  assign _T_261 = $unsigned(_T_260); // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7436.6]
  assign _T_262 = _T_261[3:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 202:56:@7437.6]
  assign _T_263 = _T_302 ? io_pixel_planar0_bundle_limit : _T_262; // @[NV_NVDLA_CDMA_IMG_sg.scala 201:37:@7438.6]
  assign _T_264 = _T_259 ? io_pixel_planar0_bundle_limit_1st : _T_263; // @[NV_NVDLA_CDMA_IMG_sg.scala 200:37:@7439.6]
  assign _T_453 = _T_449 & _T_417; // @[NV_NVDLA_CDMA_IMG_sg.scala 296:63:@7606.4]
  assign _T_454 = _T_171 | _T_453; // @[NV_NVDLA_CDMA_IMG_sg.scala 296:45:@7607.4]
  assign _GEN_12 = _T_454 ? _T_264 : _T_250; // @[NV_NVDLA_CDMA_IMG_sg.scala 199:30:@7433.4]
  assign _GEN_64 = {{10'd0}, io_pixel_planar0_lp_burst}; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:50:@7454.4]
  assign _T_281 = _T_267 == _GEN_64; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:50:@7454.4]
  assign _T_283 = _T_270 == 2'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:101:@7455.4]
  assign _T_284 = _T_281 & _T_283; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:80:@7456.4]
  assign _T_285 = _T_267 == io_pixel_planar0_width_burst; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:50:@7457.4]
  assign _T_288 = _T_285 & _T_293; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:83:@7459.4]
  assign _T_289 = ~ io_pixel_planar0_lp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:114:@7460.4]
  assign _T_290 = _T_288 & _T_289; // @[NV_NVDLA_CDMA_IMG_sg.scala 215:112:@7461.4]
  assign _T_291 = _T_284 | _T_290; // @[NV_NVDLA_CDMA_IMG_sg.scala 214:110:@7462.4]
  assign _T_306 = _T_259 & io_pixel_planar0_lp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 223:75:@7477.6]
  assign _T_309 = _T_259 & _T_289; // @[NV_NVDLA_CDMA_IMG_sg.scala 224:75:@7480.6]
  assign _T_312 = _T_283 & _T_280; // @[NV_NVDLA_CDMA_IMG_sg.scala 225:65:@7482.6]
  assign _T_315 = _T_293 & _T_280; // @[NV_NVDLA_CDMA_IMG_sg.scala 226:65:@7484.6]
  assign _T_316 = _T_276[13:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 227:57:@7485.6]
  assign _T_317 = _T_315 ? {{10'd0}, io_pixel_planar0_rp_burst} : _T_316; // @[NV_NVDLA_CDMA_IMG_sg.scala 226:36:@7486.6]
  assign _T_318 = _T_312 ? io_pixel_planar0_width_burst : _T_317; // @[NV_NVDLA_CDMA_IMG_sg.scala 225:36:@7487.6]
  assign _T_319 = _T_309 ? io_pixel_planar0_width_burst : _T_318; // @[NV_NVDLA_CDMA_IMG_sg.scala 224:36:@7488.6]
  assign _T_320 = _T_306 ? {{10'd0}, io_pixel_planar0_lp_burst} : _T_319; // @[NV_NVDLA_CDMA_IMG_sg.scala 223:36:@7489.6]
  assign _GEN_13 = _T_454 ? _T_320 : _T_267; // @[NV_NVDLA_CDMA_IMG_sg.scala 222:30:@7475.4]
  assign _T_328 = _T_270 + 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 232:50:@7497.6]
  assign _T_329 = _T_270 + 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 232:50:@7498.6]
  assign _T_330 = _T_306 ? 2'h1 : _T_329; // @[NV_NVDLA_CDMA_IMG_sg.scala 231:34:@7499.6]
  assign _T_331 = _T_306 ? 2'h0 : _T_330; // @[NV_NVDLA_CDMA_IMG_sg.scala 230:34:@7500.6]
  assign _T_457 = _T_453 & _T_280; // @[NV_NVDLA_CDMA_IMG_sg.scala 297:83:@7611.4]
  assign _T_458 = _T_171 | _T_457; // @[NV_NVDLA_CDMA_IMG_sg.scala 297:43:@7612.4]
  assign _GEN_14 = _T_458 ? _T_331 : _T_270; // @[NV_NVDLA_CDMA_IMG_sg.scala 229:28:@7492.4]
  assign _GEN_65 = {{11'd0}, io_pixel_planar1_lp_burst}; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:50:@7520.4]
  assign _T_357 = _T_337 == _GEN_65; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:50:@7520.4]
  assign _T_359 = _T_340 == 2'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:103:@7521.4]
  assign _T_360 = _T_357 & _T_359; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:81:@7522.4]
  assign _T_361 = _T_337 == io_pixel_planar1_width_burst; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:50:@7523.4]
  assign _T_364 = _T_361 & _T_369; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:84:@7525.4]
  assign _T_365 = ~ io_pixel_planar1_lp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:117:@7526.4]
  assign _T_366 = _T_364 & _T_365; // @[NV_NVDLA_CDMA_IMG_sg.scala 249:115:@7527.4]
  assign _T_367 = _T_360 | _T_366; // @[NV_NVDLA_CDMA_IMG_sg.scala 248:113:@7528.4]
  assign _T_381 = _T_171 | _T_376; // @[NV_NVDLA_CDMA_IMG_sg.scala 256:56:@7540.6]
  assign _T_382 = _T_334 - _T_353; // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7541.6]
  assign _T_383 = $unsigned(_T_382); // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7542.6]
  assign _T_384 = _T_383[4:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 258:55:@7543.6]
  assign _T_385 = _T_378 ? io_pixel_planar1_bundle_limit : _T_384; // @[NV_NVDLA_CDMA_IMG_sg.scala 257:37:@7544.6]
  assign _T_386 = _T_381 ? io_pixel_planar1_bundle_limit_1st : _T_385; // @[NV_NVDLA_CDMA_IMG_sg.scala 256:37:@7545.6]
  assign _T_388 = _T_381 & io_pixel_planar1_lp_vld; // @[NV_NVDLA_CDMA_IMG_sg.scala 259:75:@7548.6]
  assign _T_391 = _T_381 & _T_365; // @[NV_NVDLA_CDMA_IMG_sg.scala 260:75:@7551.6]
  assign _T_394 = _T_359 & _T_356; // @[NV_NVDLA_CDMA_IMG_sg.scala 261:66:@7553.6]
  assign _T_397 = _T_369 & _T_356; // @[NV_NVDLA_CDMA_IMG_sg.scala 262:66:@7555.6]
  assign _T_398 = _T_350[13:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 263:57:@7556.6]
  assign _T_399 = _T_397 ? {{11'd0}, io_pixel_planar1_rp_burst} : _T_398; // @[NV_NVDLA_CDMA_IMG_sg.scala 262:36:@7557.6]
  assign _T_400 = _T_394 ? io_pixel_planar1_width_burst : _T_399; // @[NV_NVDLA_CDMA_IMG_sg.scala 261:36:@7558.6]
  assign _T_401 = _T_391 ? io_pixel_planar1_width_burst : _T_400; // @[NV_NVDLA_CDMA_IMG_sg.scala 260:36:@7559.6]
  assign _T_402 = _T_388 ? {{11'd0}, io_pixel_planar1_lp_burst} : _T_401; // @[NV_NVDLA_CDMA_IMG_sg.scala 259:36:@7560.6]
  assign _T_459 = _T_449 & _T_240; // @[NV_NVDLA_CDMA_IMG_sg.scala 298:63:@7614.4]
  assign _T_460 = _T_171 | _T_459; // @[NV_NVDLA_CDMA_IMG_sg.scala 298:45:@7615.4]
  assign _GEN_15 = _T_460 ? _T_386 : _T_334; // @[NV_NVDLA_CDMA_IMG_sg.scala 255:30:@7539.4]
  assign _GEN_16 = _T_460 ? _T_402 : _T_337; // @[NV_NVDLA_CDMA_IMG_sg.scala 255:30:@7539.4]
  assign _T_411 = _T_340 + 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 268:50:@7569.6]
  assign _T_412 = _T_340 + 2'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 268:50:@7570.6]
  assign _T_413 = _T_391 ? 2'h1 : _T_412; // @[NV_NVDLA_CDMA_IMG_sg.scala 267:34:@7571.6]
  assign _T_414 = _T_388 ? 2'h0 : _T_413; // @[NV_NVDLA_CDMA_IMG_sg.scala 266:34:@7572.6]
  assign _T_462 = _T_459 & _T_356; // @[NV_NVDLA_CDMA_IMG_sg.scala 299:82:@7618.4]
  assign _T_463 = _T_171 | _T_462; // @[NV_NVDLA_CDMA_IMG_sg.scala 299:43:@7619.4]
  assign _GEN_17 = _T_463 ? _T_414 : _T_340; // @[NV_NVDLA_CDMA_IMG_sg.scala 265:28:@7563.4]
  assign _T_416 = _T_417 ? _T_291 : _T_367; // @[NV_NVDLA_CDMA_IMG_sg.scala 272:31:@7576.4]
  assign _T_422 = _T_417 ? {{1'd0}, _T_279} : _T_353; // @[NV_NVDLA_CDMA_IMG_sg.scala 275:33:@7582.4]
  assign _T_424 = ~ _T_293; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:49:@7584.4]
  assign _T_425 = ~ _T_369; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:66:@7585.4]
  assign _T_426 = _T_417 ? _T_424 : _T_425; // @[NV_NVDLA_CDMA_IMG_sg.scala 276:27:@7586.4]
  assign _T_439 = ~ io_is_running; // @[NV_NVDLA_CDMA_IMG_sg.scala 285:27:@7592.4]
  assign _T_450 = _T_418 & _T_243; // @[NV_NVDLA_CDMA_IMG_sg.scala 293:39:@7601.4]
  assign _T_451 = _T_450 & _T_232; // @[NV_NVDLA_CDMA_IMG_sg.scala 293:60:@7602.4]
  assign _T_442 = _T_449 & _T_451; // @[NV_NVDLA_CDMA_IMG_sg.scala 287:38:@7593.4]
  assign _T_444 = _T_442 ? 1'h0 : _T_433; // @[NV_NVDLA_CDMA_IMG_sg.scala 287:26:@7594.4]
  assign _T_445 = _T_171 ? 1'h1 : _T_444; // @[NV_NVDLA_CDMA_IMG_sg.scala 286:26:@7595.4]
  assign _T_446 = _T_439 ? 1'h0 : _T_445; // @[NV_NVDLA_CDMA_IMG_sg.scala 285:26:@7596.4]
  assign _T_466 = _T_293 | _T_300; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:113:@7623.4]
  assign _T_467 = _T_453 & _T_466; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:95:@7624.4]
  assign _T_468 = _T_171 | _T_467; // @[NV_NVDLA_CDMA_IMG_sg.scala 300:55:@7625.4]
  assign _T_470 = _T_369 | _T_376; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:112:@7627.4]
  assign _T_471 = _T_459 & _T_470; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:94:@7628.4]
  assign _T_472 = _T_171 | _T_471; // @[NV_NVDLA_CDMA_IMG_sg.scala 301:55:@7629.4]
  assign _T_485 = _T_480 + io_reg2dp_line_stride; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:99:@7640.6]
  assign _T_486 = _T_480 + io_reg2dp_line_stride; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:99:@7641.6]
  assign _T_487 = _T_171 ? 32'h0 : _T_486; // @[NV_NVDLA_CDMA_IMG_sg.scala 310:38:@7642.6]
  assign _GEN_18 = _T_477 ? _T_487 : _T_480; // @[NV_NVDLA_CDMA_IMG_sg.scala 309:24:@7639.4]
  assign _T_488 = _T_477 & io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_sg.scala 312:24:@7645.4]
  assign _T_490 = _T_480 + io_reg2dp_uv_line_stride; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:99:@7647.6]
  assign _T_491 = _T_480 + io_reg2dp_uv_line_stride; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:99:@7648.6]
  assign _T_492 = _T_171 ? 32'h0 : _T_491; // @[NV_NVDLA_CDMA_IMG_sg.scala 313:38:@7649.6]
  assign _GEN_19 = _T_488 ? _T_492 : _T_483; // @[NV_NVDLA_CDMA_IMG_sg.scala 312:41:@7646.4]
  assign _GEN_66 = {{23'd0}, _T_279}; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7656.6]
  assign _T_501 = _T_495 + _GEN_66; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7656.6]
  assign _T_502 = _T_495 + _GEN_66; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:134:@7657.6]
  assign _T_503 = _T_259 ? 27'h0 : _T_502; // @[NV_NVDLA_CDMA_IMG_sg.scala 320:39:@7658.6]
  assign _GEN_20 = _T_468 ? _T_503 : _T_495; // @[NV_NVDLA_CDMA_IMG_sg.scala 319:37:@7654.4]
  assign _GEN_67 = {{22'd0}, _T_353}; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7663.6]
  assign _T_506 = _T_498 + _GEN_67; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7663.6]
  assign _T_507 = _T_498 + _GEN_67; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:134:@7664.6]
  assign _T_508 = _T_381 ? 27'h0 : _T_507; // @[NV_NVDLA_CDMA_IMG_sg.scala 323:39:@7665.6]
  assign _GEN_21 = _T_472 ? _T_508 : _T_498; // @[NV_NVDLA_CDMA_IMG_sg.scala 322:37:@7661.4]
  assign _GEN_68 = {{32'd0}, _T_480}; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7670.4]
  assign _T_513 = _T_510 + _GEN_68; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7670.4]
  assign _T_514 = _T_510 + _GEN_68; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:48:@7671.4]
  assign _T_516 = {_T_495,1'h0}; // @[Cat.scala 30:58:@7672.4]
  assign _GEN_69 = {{36'd0}, _T_516}; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7673.4]
  assign _T_517 = _T_514 + _GEN_69; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7673.4]
  assign _T_518 = _T_514 + _GEN_69; // @[NV_NVDLA_CDMA_IMG_sg.scala 330:73:@7674.4]
  assign _GEN_70 = {{32'd0}, _T_483}; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7675.4]
  assign _T_519 = _T_512 + _GEN_70; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7675.4]
  assign _T_520 = _T_512 + _GEN_70; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:48:@7676.4]
  assign _T_522 = {_T_498,1'h0}; // @[Cat.scala 30:58:@7677.4]
  assign _GEN_71 = {{36'd0}, _T_522}; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7678.4]
  assign _T_523 = _T_520 + _GEN_71; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7678.4]
  assign _T_524 = _T_520 + _GEN_71; // @[NV_NVDLA_CDMA_IMG_sg.scala 331:73:@7679.4]
  assign _T_525 = {io_reg2dp_datain_addr_high_0,io_reg2dp_datain_addr_low_0}; // @[Cat.scala 30:58:@7681.6]
  assign _T_526 = {io_reg2dp_datain_addr_high_1,io_reg2dp_datain_addr_low_1}; // @[Cat.scala 30:58:@7683.6]
  assign _T_561 = _T_584 ? 1'h0 : _T_436; // @[NV_NVDLA_CDMA_IMG_sg.scala 352:29:@7697.4]
  assign _T_562 = _T_433 ? 1'h1 : _T_561; // @[NV_NVDLA_CDMA_IMG_sg.scala 351:29:@7698.4]
  assign _T_563 = _T_439 ? 1'h0 : _T_562; // @[NV_NVDLA_CDMA_IMG_sg.scala 350:29:@7699.4]
  assign _T_564 = _T_240 ? _T_524 : _T_518; // @[NV_NVDLA_CDMA_IMG_sg.scala 353:23:@7700.4]
  assign _T_566 = _T_422 - 5'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7701.4]
  assign _T_567 = $unsigned(_T_566); // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7702.4]
  assign _T_568 = _T_567[4:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 355:33:@7703.4]
  assign _T_569 = _T_420 & _T_243; // @[NV_NVDLA_CDMA_IMG_sg.scala 357:45:@7704.4]
  assign _GEN_24 = _T_449 ? _T_564 : _T_529; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_25 = _T_449 ? _T_422 : _T_532; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_26 = _T_449 ? _T_568 : _T_535; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_27 = _T_449 ? _T_416 : _T_538; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_28 = _T_449 ? _T_569 : _T_541; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_29 = _T_449 ? _T_450 : _T_544; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_30 = _T_449 ? _T_450 : _T_547; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_31 = _T_449 ? _T_451 : _T_550; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_32 = _T_449 ? _T_240 : _T_553; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _GEN_33 = _T_449 ? _T_426 : _T_556; // @[NV_NVDLA_CDMA_IMG_sg.scala 363:21:@7708.4]
  assign _T_586 = _T_436 & _T_584; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:43:@7728.4]
  assign _T_587 = _T_586 & _T_550; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:58:@7729.4]
  assign _T_589 = _T_587 ? 1'h1 : _T_581; // @[NV_NVDLA_CDMA_IMG_sg.scala 386:28:@7730.4]
  assign _T_590 = _T_171 ? 1'h0 : _T_589; // @[NV_NVDLA_CDMA_IMG_sg.scala 385:28:@7731.4]
  assign _T_594 = _T_578 | _T_581; // @[NV_NVDLA_CDMA_IMG_sg.scala 394:49:@7734.4]
  assign _T_596 = _T_231 ? _T_189 : _T_192; // @[NV_NVDLA_CDMA_IMG_sg.scala 396:33:@7735.4]
  assign _T_597 = _T_232 ? _T_195 : _T_596; // @[NV_NVDLA_CDMA_IMG_sg.scala 395:33:@7736.4]
  assign _T_598 = _T_594 ? 15'h0 : _T_597; // @[NV_NVDLA_CDMA_IMG_sg.scala 394:33:@7737.4]
  assign _GEN_72 = {{14'd0}, _T_593}; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7738.4]
  assign _T_599 = _T_598 + _GEN_72; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7738.4]
  assign _T_600 = _T_598 + _GEN_72; // @[NV_NVDLA_CDMA_IMG_sg.scala 398:51:@7739.4]
  assign _T_601 = io_status2dma_free_entries >= _T_600; // @[NV_NVDLA_CDMA_IMG_sg.scala 399:53:@7740.4]
  assign _T_603 = _T_439 | _T_171; // @[NV_NVDLA_CDMA_IMG_sg.scala 400:46:@7742.4]
  assign _T_606 = _T_586 & _T_547; // @[NV_NVDLA_CDMA_IMG_sg.scala 401:59:@7744.4]
  assign _T_608 = ~ _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 402:31:@7745.4]
  assign _T_609 = _T_608 ? _T_601 : _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 402:30:@7746.4]
  assign _T_610 = _T_606 ? 1'h0 : _T_609; // @[NV_NVDLA_CDMA_IMG_sg.scala 401:30:@7747.4]
  assign _T_611 = _T_603 ? 1'h0 : _T_610; // @[NV_NVDLA_CDMA_IMG_sg.scala 400:30:@7748.4]
  assign _T_613 = io_img2status_dat_updt ? io_img2status_dat_entries : 15'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 404:34:@7749.4]
  assign _T_614 = ~ _T_581; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:35:@7750.4]
  assign _T_615 = _T_614 & _T_601; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:48:@7751.4]
  assign _T_617 = _T_615 & _T_608; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:65:@7753.4]
  assign _T_619 = _T_617 ? _T_598 : 15'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 405:34:@7754.4]
  assign _T_620 = _GEN_72 + _T_619; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:45:@7755.4]
  assign _T_621 = _GEN_72 + _T_619; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:45:@7756.4]
  assign _T_622 = _T_621 - _T_613; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7757.4]
  assign _T_623 = $unsigned(_T_622); // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7758.4]
  assign _T_624 = _T_623[14:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 406:67:@7759.4]
  assign _T_629 = _T_617 | io_img2status_dat_updt; // @[NV_NVDLA_CDMA_IMG_sg.scala 407:79:@7764.4]
  assign _GEN_34 = _T_629 ? _T_624 : {{14'd0}, _T_593}; // @[NV_NVDLA_CDMA_IMG_sg.scala 410:29:@7766.4]
  assign _T_641 = {{10'd0}, _T_535}; // @[NV_NVDLA_CDMA_IMG_sg.scala 452:31:@7801.4 NV_NVDLA_CDMA_IMG_sg.scala 459:21:@7814.4]
  assign _T_650 = _T_436 & _T_575; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:36:@7808.4]
  assign _T_651 = _T_650 & _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:57:@7809.4]
  assign _T_652 = ~ _T_556; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:75:@7810.4]
  assign _T_653 = _T_651 & _T_652; // @[NV_NVDLA_CDMA_IMG_sg.scala 457:73:@7811.4]
  assign _T_682 = NV_NVDLA_fifo_io_rd_pd[5]; // @[NV_NVDLA_CDMA_IMG_sg.scala 498:42:@7850.4]
  assign _T_684 = NV_NVDLA_fifo_io_rd_pvld & _T_682; // @[NV_NVDLA_CDMA_IMG_sg.scala 501:43:@7852.4]
  assign _T_661 = _T_436 & _T_578; // @[NV_NVDLA_CDMA_IMG_sg.scala 480:38:@7830.4]
  assign _T_665 = {_T_538,_T_556,_T_532}; // @[Cat.scala 30:58:@7835.4]
  assign _T_668 = {_T_553,_T_550,_T_544,_T_541}; // @[Cat.scala 30:58:@7838.4]
  assign _T_635 = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 422:29:@7771.4 NV_NVDLA_CDMA_IMG_sg.scala 445:19:@7798.4]
  assign _T_670 = _T_635[255:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 488:40:@7841.4]
  assign _T_671 = _T_635[256]; // @[NV_NVDLA_CDMA_IMG_sg.scala 489:40:@7842.4]
  assign _T_677 = NV_NVDLA_fifo_io_rd_pd[10]; // @[NV_NVDLA_CDMA_IMG_sg.scala 493:43:@7845.4]
  assign _T_678 = NV_NVDLA_fifo_io_rd_pd[9]; // @[NV_NVDLA_CDMA_IMG_sg.scala 494:40:@7846.4]
  assign _T_679 = NV_NVDLA_fifo_io_rd_pd[8]; // @[NV_NVDLA_CDMA_IMG_sg.scala 495:45:@7847.4]
  assign _T_681 = NV_NVDLA_fifo_io_rd_pd[6]; // @[NV_NVDLA_CDMA_IMG_sg.scala 497:44:@7849.4]
  assign _T_683 = NV_NVDLA_fifo_io_rd_pd[4:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 499:41:@7851.4]
  assign _T_685 = ~ NV_NVDLA_fifo_io_rd_pvld; // @[NV_NVDLA_CDMA_IMG_sg.scala 503:28:@7854.4]
  assign _T_687 = ~ _T_682; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:27:@7855.4]
  assign _T_637 = NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 423:30:@7772.4 NV_NVDLA_CDMA_IMG_sg.scala 446:20:@7799.4]
  assign _T_689 = _T_637 & _T_671; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:58:@7857.4]
  assign _T_691 = _T_687 ? _T_689 : 1'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 504:26:@7858.4]
  assign _T_692 = _T_685 ? 1'h0 : _T_691; // @[NV_NVDLA_CDMA_IMG_sg.scala 503:27:@7859.4]
  assign _GEN_74 = {{4'd0}, _T_692}; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7860.4]
  assign _T_693 = _T_674 + _GEN_74; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7860.4]
  assign _T_694 = _T_674 + _GEN_74; // @[NV_NVDLA_CDMA_IMG_sg.scala 507:49:@7861.4]
  assign _T_695 = _T_694 == _T_683; // @[NV_NVDLA_CDMA_IMG_sg.scala 508:55:@7862.4]
  assign _T_697 = _T_695 ? 5'h0 : _T_694; // @[NV_NVDLA_CDMA_IMG_sg.scala 508:33:@7863.4]
  assign _T_698 = _T_682 | _T_637; // @[NV_NVDLA_CDMA_IMG_sg.scala 513:54:@7867.4]
  assign _T_699 = NV_NVDLA_fifo_io_rd_pvld & _T_698; // @[NV_NVDLA_CDMA_IMG_sg.scala 513:37:@7868.4]
  assign _GEN_35 = _T_699 ? _T_697 : _T_674; // @[NV_NVDLA_CDMA_IMG_sg.scala 510:22:@7864.4]
  assign _T_701 = _T_699 & _T_695; // @[NV_NVDLA_CDMA_IMG_sg.scala 514:40:@7871.4]
  assign _T_713 = io_pixel_order[10]; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:41:@7882.4]
  assign _T_714 = _T_713 & _T_677; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:45:@7883.4]
  assign _T_715 = io_pixel_order[9]; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:76:@7884.4]
  assign _T_716 = _T_715 & _T_677; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:79:@7885.4]
  assign _T_717 = io_pixel_order[8:1]; // @[NV_NVDLA_CDMA_IMG_sg.scala 545:110:@7886.4]
  assign _T_718 = io_pixel_order[0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:39:@7887.4]
  assign _T_719 = ~ _T_677; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:44:@7888.4]
  assign _T_720 = _T_719 & io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:60:@7889.4]
  assign _T_721 = _T_718 | _T_720; // @[NV_NVDLA_CDMA_IMG_sg.scala 546:42:@7890.4]
  assign _T_724 = {_T_714,_T_716,_T_717,_T_721}; // @[Cat.scala 30:58:@7893.4]
  assign _T_1041 = _T_724[0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:67:@8190.4]
  assign _T_1045 = _T_1041 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@8192.4]
  assign _T_1046 = _T_1045 & _T_670; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:72:@8193.4]
  assign _T_1047 = _T_724[1]; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:66:@8194.4]
  assign _T_1051 = _T_1047 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@8196.4]
  assign _T_774 = _T_670[255:248]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7943.4]
  assign _T_775 = _T_670[231:224]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7944.4]
  assign _T_776 = _T_670[239:232]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7945.4]
  assign _T_777 = _T_670[247:240]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7946.4]
  assign _T_767 = _T_670[223:216]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7936.4]
  assign _T_768 = _T_670[199:192]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7937.4]
  assign _T_769 = _T_670[207:200]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7938.4]
  assign _T_770 = _T_670[215:208]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7939.4]
  assign _T_760 = _T_670[191:184]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7929.4]
  assign _T_761 = _T_670[167:160]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7930.4]
  assign _T_762 = _T_670[175:168]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7931.4]
  assign _T_763 = _T_670[183:176]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7932.4]
  assign _T_753 = _T_670[159:152]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7922.4]
  assign _T_754 = _T_670[135:128]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7923.4]
  assign _T_755 = _T_670[143:136]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7924.4]
  assign _T_756 = _T_670[151:144]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7925.4]
  assign _T_798 = {_T_760,_T_761,_T_762,_T_763,_T_753,_T_754,_T_755,_T_756}; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7962.4]
  assign _T_746 = _T_670[127:120]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7915.4]
  assign _T_747 = _T_670[103:96]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7916.4]
  assign _T_748 = _T_670[111:104]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7917.4]
  assign _T_749 = _T_670[119:112]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7918.4]
  assign _T_739 = _T_670[95:88]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7908.4]
  assign _T_740 = _T_670[71:64]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7909.4]
  assign _T_741 = _T_670[79:72]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7910.4]
  assign _T_742 = _T_670[87:80]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7911.4]
  assign _T_732 = _T_670[63:56]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7901.4]
  assign _T_733 = _T_670[39:32]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7902.4]
  assign _T_734 = _T_670[47:40]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7903.4]
  assign _T_735 = _T_670[55:48]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7904.4]
  assign _T_725 = _T_670[31:24]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:26:@7894.4]
  assign _T_726 = _T_670[7:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:53:@7895.4]
  assign _T_727 = _T_670[15:8]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:76:@7896.4]
  assign _T_728 = _T_670[23:16]; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:102:@7897.4]
  assign _T_795 = {_T_732,_T_733,_T_734,_T_735,_T_725,_T_726,_T_727,_T_728}; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7959.4]
  assign _T_797 = {_T_746,_T_747,_T_748,_T_749,_T_739,_T_740,_T_741,_T_742,_T_795}; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7961.4]
  assign _T_801 = {_T_774,_T_775,_T_776,_T_777,_T_767,_T_768,_T_769,_T_770,_T_798,_T_797}; // @[NV_NVDLA_CDMA_IMG_sg.scala 551:124:@7965.4]
  assign _T_1052 = _T_1051 & _T_801; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:71:@8197.4]
  assign _T_1053 = _T_1046 | _T_1052; // @[NV_NVDLA_CDMA_IMG_sg.scala 559:94:@8198.4]
  assign _T_1054 = _T_724[3]; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:66:@8199.4]
  assign _T_1058 = _T_1054 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@8201.4]
  assign _T_875 = {_T_761,_T_760,_T_763,_T_762,_T_754,_T_753,_T_756,_T_755}; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8034.4]
  assign _T_872 = {_T_733,_T_732,_T_735,_T_734,_T_726,_T_725,_T_728,_T_727}; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8031.4]
  assign _T_874 = {_T_747,_T_746,_T_749,_T_748,_T_740,_T_739,_T_742,_T_741,_T_872}; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8033.4]
  assign _T_878 = {_T_775,_T_774,_T_777,_T_776,_T_768,_T_767,_T_770,_T_769,_T_875,_T_874}; // @[NV_NVDLA_CDMA_IMG_sg.scala 553:124:@8037.4]
  assign _T_1059 = _T_1058 & _T_878; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:71:@8202.4]
  assign _T_1060 = _T_1053 | _T_1059; // @[NV_NVDLA_CDMA_IMG_sg.scala 560:93:@8203.4]
  assign _T_1061 = _T_724[5]; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:66:@8204.4]
  assign _T_1065 = _T_1061 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@8206.4]
  assign _T_952 = {_T_761,_T_762,_T_763,_T_760,_T_754,_T_755,_T_756,_T_753}; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8106.4]
  assign _T_949 = {_T_733,_T_734,_T_735,_T_732,_T_726,_T_727,_T_728,_T_725}; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8103.4]
  assign _T_951 = {_T_747,_T_748,_T_749,_T_746,_T_740,_T_741,_T_742,_T_739,_T_949}; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8105.4]
  assign _T_955 = {_T_775,_T_776,_T_777,_T_774,_T_768,_T_769,_T_770,_T_767,_T_952,_T_951}; // @[NV_NVDLA_CDMA_IMG_sg.scala 555:124:@8109.4]
  assign _T_1066 = _T_1065 & _T_955; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:71:@8207.4]
  assign _T_1067 = _T_1060 | _T_1066; // @[NV_NVDLA_CDMA_IMG_sg.scala 561:93:@8208.4]
  assign _T_1068 = _T_724[9]; // @[NV_NVDLA_CDMA_IMG_sg.scala 563:66:@8209.4]
  assign _T_1072 = _T_1068 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@8211.4]
  assign _T_1035 = {_T_763,_T_760,_T_761,_T_762,_T_756,_T_753,_T_754,_T_755}; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8184.4]
  assign _T_1028 = {_T_735,_T_732,_T_733,_T_734,_T_728,_T_725,_T_726,_T_727}; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8177.4]
  assign _T_1032 = {_T_749,_T_746,_T_747,_T_748,_T_742,_T_739,_T_740,_T_741,_T_1028}; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8181.4]
  assign _T_1040 = {_T_777,_T_774,_T_775,_T_776,_T_770,_T_767,_T_768,_T_769,_T_1035,_T_1032}; // @[NV_NVDLA_CDMA_IMG_sg.scala 557:70:@8189.4]
  assign _T_1073 = _T_1072 & _T_1040; // @[NV_NVDLA_CDMA_IMG_sg.scala 563:71:@8212.4]
  assign _T_1074 = _T_1067 | _T_1073; // @[NV_NVDLA_CDMA_IMG_sg.scala 562:93:@8213.4]
  assign _T_1076 = _T_674 == 5'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 566:67:@8215.4]
  assign _T_1077 = _T_681 & _T_1076; // @[NV_NVDLA_CDMA_IMG_sg.scala 566:47:@8216.4]
  assign _GEN_37 = _T_699 ? _T_677 : _T_1080; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  assign _GEN_38 = _T_699 ? _T_1077 : _T_1083; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  assign _GEN_39 = _T_699 ? _T_701 : _T_1086; // @[NV_NVDLA_CDMA_IMG_sg.scala 572:24:@8221.4]
  assign _T_1102 = _T_699 & _T_701; // @[NV_NVDLA_CDMA_IMG_sg.scala 583:24:@8231.4]
  assign _GEN_40 = _T_1102 ? _T_683 : _T_1092; // @[NV_NVDLA_CDMA_IMG_sg.scala 583:45:@8232.4]
  assign _T_1103 = _T_679 & _T_701; // @[NV_NVDLA_CDMA_IMG_sg.scala 587:46:@8236.6]
  assign _T_1105 = _T_678 & _T_701; // @[NV_NVDLA_CDMA_IMG_sg.scala 589:36:@8240.6]
  assign _GEN_41 = _T_699 ? _T_1103 : _T_1095; // @[NV_NVDLA_CDMA_IMG_sg.scala 586:24:@8235.4]
  assign _GEN_43 = _T_699 ? _T_1105 : _T_1101; // @[NV_NVDLA_CDMA_IMG_sg.scala 586:24:@8235.4]
  assign _T_1106 = ~ _T_1080; // @[NV_NVDLA_CDMA_IMG_sg.scala 596:49:@8243.4]
  assign _T_1107 = _T_710 & _T_1106; // @[NV_NVDLA_CDMA_IMG_sg.scala 596:46:@8244.4]
  assign _T_1108 = _T_710 & _T_1080; // @[NV_NVDLA_CDMA_IMG_sg.scala 597:46:@8245.4]
  assign _GEN_44 = _T_1107 ? _T_712 : _T_1111; // @[NV_NVDLA_CDMA_IMG_sg.scala 603:29:@8248.4]
  assign _GEN_45 = _T_1108 ? _T_712 : _T_1114; // @[NV_NVDLA_CDMA_IMG_sg.scala 606:29:@8251.4]
  assign _T_1122 = ~ _T_1083; // @[NV_NVDLA_CDMA_IMG_sg.scala 615:49:@8257.4]
  assign _T_1123 = _T_710 & _T_1122; // @[NV_NVDLA_CDMA_IMG_sg.scala 615:46:@8258.4]
  assign _T_1124 = _T_1107 ? _T_1111 : _T_1114; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:62:@8259.4]
  assign _T_1131 = _T_1080 ? io_pixel_planar1_byte_sft : io_pixel_planar0_byte_sft; // @[NV_NVDLA_CDMA_IMG_sg.scala 624:23:@8268.4]
  assign _T_1126 = {_T_1131,3'h0}; // @[Cat.scala 30:58:@8260.4]
  assign _T_1127 = _T_1124 >> _T_1126; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:128:@8261.4]
  assign _T_1128 = {_T_712,_T_1127}; // @[Cat.scala 30:58:@8262.4]
  assign _T_1129 = _T_1128[255:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 617:165:@8263.4]
  assign _T_1141 = _T_1134 + 7'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 631:61:@8273.4]
  assign _T_1142 = _T_1134 + 7'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 631:61:@8274.4]
  assign _T_1143 = _T_1137 + 7'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 632:61:@8275.4]
  assign _T_1144 = _T_1137 + 7'h1; // @[NV_NVDLA_CDMA_IMG_sg.scala 632:61:@8276.4]
  assign _T_1146 = _T_171 ? 7'h0 : _T_1142; // @[NV_NVDLA_CDMA_IMG_sg.scala 633:39:@8277.4]
  assign _T_1148 = _T_171 ? 7'h0 : _T_1144; // @[NV_NVDLA_CDMA_IMG_sg.scala 634:39:@8278.4]
  assign _T_1150 = _T_1123 & _T_1106; // @[NV_NVDLA_CDMA_IMG_sg.scala 635:73:@8280.4]
  assign _T_1151 = _T_171 | _T_1150; // @[NV_NVDLA_CDMA_IMG_sg.scala 635:50:@8281.4]
  assign _T_1152 = _T_1123 & _T_1080; // @[NV_NVDLA_CDMA_IMG_sg.scala 636:73:@8282.4]
  assign _T_1153 = _T_171 | _T_1152; // @[NV_NVDLA_CDMA_IMG_sg.scala 636:50:@8283.4]
  assign _T_1156 = _T_1134[0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:83:@8285.4]
  assign _T_1157 = _T_1134[6:1]; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:110:@8286.4]
  assign _T_1159 = {1'h0,_T_1156,_T_1157}; // @[Cat.scala 30:58:@8288.4]
  assign _T_1161 = _T_1137[0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 638:60:@8289.4]
  assign _T_1162 = _T_1137[6:1]; // @[NV_NVDLA_CDMA_IMG_sg.scala 638:87:@8290.4]
  assign _T_1164 = {1'h1,_T_1161,_T_1162}; // @[Cat.scala 30:58:@8292.4]
  assign _T_1165 = _T_1106 ? _T_1159 : _T_1164; // @[NV_NVDLA_CDMA_IMG_sg.scala 637:30:@8293.4]
  assign _GEN_47 = _T_1151 ? _T_1146 : _T_1134; // @[NV_NVDLA_CDMA_IMG_sg.scala 640:32:@8294.4]
  assign _GEN_48 = _T_1153 ? _T_1148 : _T_1137; // @[NV_NVDLA_CDMA_IMG_sg.scala 643:32:@8297.4]
  assign _GEN_49 = _T_1123 ? _T_1165 : _T_1140; // @[NV_NVDLA_CDMA_IMG_sg.scala 646:30:@8300.4]
  assign _T_1187 = _T_1092[3:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:79:@8310.4]
  assign _T_1188 = _T_1168 + _T_1187; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:57:@8311.4]
  assign _T_1189 = _T_1168 + _T_1187; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:57:@8312.4]
  assign _GEN_75 = {{3'd0}, _T_1086}; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8313.4]
  assign _T_1190 = _T_1189 - _GEN_75; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8313.4]
  assign _T_1191 = $unsigned(_T_1190); // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8314.4]
  assign _T_1192 = _T_1191[3:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 659:86:@8315.4]
  assign _T_1193 = _T_1171 + _T_1092; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:57:@8316.4]
  assign _T_1194 = _T_1171 + _T_1092; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:57:@8317.4]
  assign _GEN_76 = {{4'd0}, _T_1086}; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8318.4]
  assign _T_1195 = _T_1194 - _GEN_76; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8318.4]
  assign _T_1196 = $unsigned(_T_1195); // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8319.4]
  assign _T_1197 = _T_1196[4:0]; // @[NV_NVDLA_CDMA_IMG_sg.scala 660:80:@8320.4]
  assign _T_1202 = _T_1106 ? _T_1192 : _T_1168; // @[NV_NVDLA_CDMA_IMG_sg.scala 663:37:@8323.4]
  assign _T_1204 = _T_171 ? 4'h0 : _T_1202; // @[NV_NVDLA_CDMA_IMG_sg.scala 661:37:@8325.4]
  assign _T_1208 = _T_1080 ? _T_1197 : _T_1171; // @[NV_NVDLA_CDMA_IMG_sg.scala 667:37:@8327.4]
  assign _T_1210 = _T_171 ? 5'h0 : _T_1208; // @[NV_NVDLA_CDMA_IMG_sg.scala 665:37:@8329.4]
  assign _GEN_50 = _T_171 ? _T_1204 : _T_1168; // @[NV_NVDLA_CDMA_IMG_sg.scala 677:34:@8343.4]
  assign _GEN_51 = _T_171 ? _T_1210 : _T_1171; // @[NV_NVDLA_CDMA_IMG_sg.scala 680:34:@8346.4]
  assign _GEN_52 = _T_171 ? _T_1202 : _T_1174; // @[NV_NVDLA_CDMA_IMG_sg.scala 683:35:@8349.4]
  assign _GEN_53 = _T_171 ? _T_1197 : _T_1177; // @[NV_NVDLA_CDMA_IMG_sg.scala 686:35:@8352.4]
  assign _T_1228 = _T_1101 & _T_1095; // @[NV_NVDLA_CDMA_IMG_sg.scala 698:45:@8361.4]
  assign _T_1230 = _T_1228 ? 1'h1 : _T_1226; // @[NV_NVDLA_CDMA_IMG_sg.scala 698:32:@8362.4]
  assign _T_1231 = _T_171 ? 1'h0 : _T_1230; // @[NV_NVDLA_CDMA_IMG_sg.scala 697:32:@8363.4]
  assign _GEN_56 = io_is_running ? _T_1231 : _T_1226; // @[NV_NVDLA_CDMA_IMG_sg.scala 700:24:@8364.4]
  assign _T_1234 = {_T_1177,_T_1174}; // @[Cat.scala 30:58:@8372.4]
  assign _T_1244 = ~ _T_171; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:24:@8399.4]
  assign _T_1245 = _T_1244 & _T_581; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:42:@8400.4]
  assign _T_1246 = _T_1245 & _T_1226; // @[NV_NVDLA_CDMA_IMG_sg.scala 758:56:@8401.4]
  assign _GEN_57 = io_is_running ? _T_1246 : _T_1243; // @[NV_NVDLA_CDMA_IMG_sg.scala 760:24:@8402.4]
  assign _T_1247 = ~ _T_573; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:53:@8406.4]
  assign _T_1248 = _T_653 & _T_1247; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:51:@8407.4]
  assign _T_1249 = _T_1248 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_IMG_sg.scala 769:69:@8408.4]
  assign _T_1253 = io_status2dma_fsm_switch & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_IMG_sg.scala 770:61:@8411.4]
  assign _T_1257 = io_reg2dp_op_en & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_IMG_sg.scala 771:52:@8414.4]
  assign _T_1269 = _T_701 & _T_687; // @[NV_NVDLA_CDMA_IMG_sg.scala 785:57:@8432.4]
  assign _T_1270 = _T_1269 & io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_IMG_sg.scala 785:74:@8433.4]
  assign _T_1282 = NV_COUNTER_STAGE_histogram_1_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 789:42:@8441.4 NV_NVDLA_CDMA_IMG_sg.scala 799:32:@8454.4]
  assign _T_1284 = _T_1282 != 9'h1ff; // @[NV_NVDLA_CDMA_IMG_sg.scala 790:49:@8442.4]
  assign _T_1289 = ~ io_dp2reg_img_rd_latency; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:48:@8455.4]
  assign _T_1291 = _T_1289 == 32'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:48:@8456.4]
  assign _T_1292 = ~ _T_1291; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:22:@8457.4]
  assign _T_1294 = _T_1282 != 9'h0; // @[NV_NVDLA_CDMA_IMG_sg.scala 802:84:@8458.4]
  assign io_img_dat2mcif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 432:31:@7783.4]
  assign io_img_dat2mcif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 432:31:@7782.4]
  assign io_mcif2img_dat_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 443:47:@7797.4]
  assign io_img_dat2cvif_rd_req_pd_valid = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 430:39:@7780.4]
  assign io_img_dat2cvif_rd_req_pd_bits = NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 430:39:@7779.4]
  assign io_cvif2img_dat_rd_rsp_pd_ready = NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 441:55:@7794.4]
  assign io_sg2pack_img_pd_valid = NV_NVDLA_fifo_1_io_rd_pvld; // @[NV_NVDLA_CDMA_IMG_sg.scala 725:29:@8377.4]
  assign io_sg2pack_img_pd_bits = NV_NVDLA_fifo_1_io_rd_pd; // @[NV_NVDLA_CDMA_IMG_sg.scala 726:28:@8378.4]
  assign io_sg2pack_data_entries = _T_169; // @[NV_NVDLA_CDMA_IMG_sg.scala 745:29:@8391.4]
  assign io_sg2pack_entry_end = _T_195; // @[NV_NVDLA_CDMA_IMG_sg.scala 748:26:@8394.4]
  assign io_sg2pack_entry_mid = _T_192; // @[NV_NVDLA_CDMA_IMG_sg.scala 747:26:@8393.4]
  assign io_sg2pack_entry_st = _T_189; // @[NV_NVDLA_CDMA_IMG_sg.scala 746:25:@8392.4]
  assign io_sg2pack_height_total = _T_166; // @[NV_NVDLA_CDMA_IMG_sg.scala 743:29:@8389.4]
  assign io_sg2pack_mn_enable = _T_160; // @[NV_NVDLA_CDMA_IMG_sg.scala 744:26:@8390.4]
  assign io_sg2pack_sub_h_end = _T_186; // @[NV_NVDLA_CDMA_IMG_sg.scala 751:26:@8397.4]
  assign io_sg2pack_sub_h_mid = _T_183; // @[NV_NVDLA_CDMA_IMG_sg.scala 750:26:@8396.4]
  assign io_sg2pack_sub_h_st = _T_180; // @[NV_NVDLA_CDMA_IMG_sg.scala 749:25:@8395.4]
  assign io_sg_is_done = _T_1243; // @[NV_NVDLA_CDMA_IMG_sg.scala 763:19:@8405.4]
  assign io_img2sbuf_p0_wr_addr_valid = _T_1117; // @[NV_NVDLA_CDMA_IMG_sg.scala 706:34:@8367.4]
  assign io_img2sbuf_p0_wr_addr_bits = {{9'd0}, _T_1140}; // @[NV_NVDLA_CDMA_IMG_sg.scala 707:33:@8368.4]
  assign io_img2sbuf_p0_wr_data = _T_1119; // @[NV_NVDLA_CDMA_IMG_sg.scala 708:28:@8369.4]
  assign io_dp2reg_img_rd_stall = NV_COUNTER_STAGE_histogram_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 781:28:@8425.4]
  assign io_dp2reg_img_rd_latency = NV_COUNTER_STAGE_histogram_2_io_cnt_cur; // @[NV_NVDLA_CDMA_IMG_sg.scala 811:30:@8468.4]
  assign NV_NVDLA_DMAIF_rdreq_reset = reset; // @[:@7776.4]
  assign NV_NVDLA_DMAIF_rdreq_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 427:47:@7777.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_valid = _T_651 & _T_652; // @[NV_NVDLA_CDMA_IMG_sg.scala 435:54:@7786.4]
  assign NV_NVDLA_DMAIF_rdreq_io_dmaif_rd_req_pd_bits = {_T_641,_T_529}; // @[NV_NVDLA_CDMA_IMG_sg.scala 434:53:@7785.4]
  assign NV_NVDLA_DMAIF_rdreq_io_mcif_rd_req_pd_ready = io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 432:31:@7784.4]
  assign NV_NVDLA_DMAIF_rdreq_io_cvif_rd_req_pd_ready = io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 430:39:@7781.4]
  assign NV_NVDLA_DMAIF_rdreq_io_reg2dp_src_ram_type = io_reg2dp_datain_ram_type; // @[NV_NVDLA_CDMA_IMG_sg.scala 428:52:@7778.4]
  assign NV_NVDLA_DMAIF_rdrsp_reset = reset; // @[:@7790.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 439:47:@7791.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_valid = io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 443:47:@7796.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_mcif_rd_rsp_pd_bits = io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 443:47:@7795.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_valid = io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_IMG_sg.scala 441:55:@7793.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_cvif_rd_rsp_pd_bits = io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_IMG_sg.scala 441:55:@7792.4]
  assign NV_NVDLA_DMAIF_rdrsp_io_dmaif_rd_rsp_pd_ready = ~ _T_684; // @[NV_NVDLA_CDMA_IMG_sg.scala 447:54:@7800.4]
  assign NV_NVDLA_fifo_clock = io_nvdla_core_clk; // @[:@7822.4]
  assign NV_NVDLA_fifo_reset = reset; // @[:@7823.4]
  assign NV_NVDLA_fifo_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 470:37:@7824.4]
  assign NV_NVDLA_fifo_io_wr_pvld = _T_661 & _T_582; // @[NV_NVDLA_CDMA_IMG_sg.scala 472:41:@7826.4]
  assign NV_NVDLA_fifo_io_wr_pd = {_T_668,_T_665}; // @[NV_NVDLA_CDMA_IMG_sg.scala 474:39:@7828.4]
  assign NV_NVDLA_fifo_io_rd_prdy = _T_699 & _T_695; // @[NV_NVDLA_CDMA_IMG_sg.scala 476:41:@7829.4]
  assign NV_NVDLA_fifo_1_clock = io_nvdla_core_clk; // @[:@8380.4]
  assign NV_NVDLA_fifo_1_reset = reset; // @[:@8381.4]
  assign NV_NVDLA_fifo_1_io_wr_pd = {2'h0,_T_1234}; // @[NV_NVDLA_CDMA_IMG_sg.scala 737:47:@8385.4]
  assign NV_NVDLA_fifo_1_io_rd_prdy = io_sg2pack_img_pd_ready; // @[NV_NVDLA_CDMA_IMG_sg.scala 739:49:@8387.4]
  assign NV_COUNTER_STAGE_histogram_reset = reset; // @[:@8419.4]
  assign NV_COUNTER_STAGE_histogram_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 776:16:@8420.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_inc = _T_1252; // @[NV_NVDLA_CDMA_IMG_sg.scala 777:25:@8421.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_clr = _T_1256; // @[NV_NVDLA_CDMA_IMG_sg.scala 779:25:@8423.4]
  assign NV_COUNTER_STAGE_histogram_io_rd_stall_cen = _T_1260; // @[NV_NVDLA_CDMA_IMG_sg.scala 780:25:@8424.4]
  assign NV_COUNTER_STAGE_histogram_1_reset = reset; // @[:@8448.4]
  assign NV_COUNTER_STAGE_histogram_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 794:18:@8449.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_inc = _T_1284 & _T_1267; // @[NV_NVDLA_CDMA_IMG_sg.scala 795:27:@8450.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_dec = _T_1284 & _T_1273; // @[NV_NVDLA_CDMA_IMG_sg.scala 796:27:@8451.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_clr = _T_1276; // @[NV_NVDLA_CDMA_IMG_sg.scala 797:27:@8452.4]
  assign NV_COUNTER_STAGE_histogram_1_io_rd_stall_cen = _T_1280; // @[NV_NVDLA_CDMA_IMG_sg.scala 798:27:@8453.4]
  assign NV_COUNTER_STAGE_histogram_2_reset = reset; // @[:@8462.4]
  assign NV_COUNTER_STAGE_histogram_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_IMG_sg.scala 806:18:@8463.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_inc = _T_1292 & _T_1294; // @[NV_NVDLA_CDMA_IMG_sg.scala 807:27:@8464.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_clr = _T_1276; // @[NV_NVDLA_CDMA_IMG_sg.scala 809:27:@8466.4]
  assign NV_COUNTER_STAGE_histogram_2_io_rd_stall_cen = _T_1280; // @[NV_NVDLA_CDMA_IMG_sg.scala 810:27:@8467.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_157 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_160 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_163 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_166 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_169 = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_180 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_183 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_186 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_189 = _RAND_8[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_192 = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_195 = _RAND_10[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_226 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_433 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_436 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_556 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_578 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_240 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_267 = _RAND_17[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_250 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_270 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_337 = _RAND_20[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_334 = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_340 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_480 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_483 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_495 = _RAND_25[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_498 = _RAND_26[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_510 = _RAND_27[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_512 = _RAND_28[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_529 = _RAND_29[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_532 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_535 = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_538 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_541 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_544 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_547 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_550 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_553 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_581 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_593 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_674 = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_710 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {8{`RANDOM}};
  _T_712 = _RAND_42[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1080 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1083 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1086 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1092 = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1095 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1101 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {8{`RANDOM}};
  _T_1111 = _RAND_49[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {8{`RANDOM}};
  _T_1114 = _RAND_50[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1117 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {8{`RANDOM}};
  _T_1119 = _RAND_52[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1134 = _RAND_53[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1137 = _RAND_54[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1140 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1168 = _RAND_56[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1171 = _RAND_57[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1174 = _RAND_58[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1177 = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1226 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1243 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1252 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1256 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1260 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1267 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1273 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1276 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1280 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_157 <= 1'h0;
    end else begin
      _T_157 <= io_is_running;
    end
    if (reset) begin
      _T_160 <= 1'h0;
    end else begin
      if (io_layer_st) begin
        _T_160 <= io_reg2dp_mean_format;
      end
    end
    if (reset) begin
      _T_163 <= 14'h0;
    end else begin
      if (io_layer_st) begin
        _T_163 <= _T_175;
      end
    end
    if (reset) begin
      _T_166 <= 13'h0;
    end else begin
      if (io_layer_st) begin
        _T_166 <= io_reg2dp_datain_height;
      end
    end
    if (reset) begin
      _T_169 <= 15'h0;
    end else begin
      if (io_layer_st) begin
        _T_169 <= _T_177;
      end
    end
    if (reset) begin
      _T_180 <= 4'h0;
    end else begin
      if (_T_171) begin
        if (_T_205) begin
          _T_180 <= _T_203;
        end else begin
          _T_180 <= 4'h1;
        end
      end
    end
    if (reset) begin
      _T_183 <= 4'h0;
    end else begin
      if (_T_171) begin
        _T_183 <= 4'h1;
      end
    end
    if (reset) begin
      _T_186 <= 4'h0;
    end else begin
      if (_T_171) begin
        if (_T_205) begin
          _T_186 <= _T_203;
        end else begin
          _T_186 <= 4'h1;
        end
      end
    end
    if (reset) begin
      _T_189 <= 15'h0;
    end else begin
      if (_T_171) begin
        _T_189 <= _T_218;
      end
    end
    if (reset) begin
      _T_192 <= 15'h0;
    end else begin
      if (_T_171) begin
        _T_192 <= _T_169;
      end
    end
    if (reset) begin
      _T_195 <= 15'h0;
    end else begin
      if (_T_171) begin
        _T_195 <= _T_218;
      end
    end
    if (reset) begin
      _T_226 <= 13'h0;
    end else begin
      if (_T_477) begin
        if (_T_171) begin
          _T_226 <= 13'h0;
        end else begin
          _T_226 <= _T_236;
        end
      end
    end
    if (reset) begin
      _T_433 <= 1'h0;
    end else begin
      if (_T_439) begin
        _T_433 <= 1'h0;
      end else begin
        if (_T_171) begin
          _T_433 <= 1'h1;
        end else begin
          if (_T_442) begin
            _T_433 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_436 <= 1'h0;
    end else begin
      if (_T_439) begin
        _T_436 <= 1'h0;
      end else begin
        if (_T_433) begin
          _T_436 <= 1'h1;
        end else begin
          if (_T_584) begin
            _T_436 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_556 <= 1'h0;
    end else begin
      if (_T_449) begin
        if (_T_417) begin
          _T_556 <= _T_424;
        end else begin
          _T_556 <= _T_425;
        end
      end
    end
    if (reset) begin
      _T_578 <= 1'h1;
    end else begin
      if (_T_603) begin
        _T_578 <= 1'h0;
      end else begin
        if (_T_606) begin
          _T_578 <= 1'h0;
        end else begin
          if (_T_608) begin
            _T_578 <= _T_601;
          end
        end
      end
    end
    if (reset) begin
      _T_240 <= 1'h0;
    end else begin
      if (_T_474) begin
        if (_T_244) begin
          _T_240 <= 1'h0;
        end else begin
          _T_240 <= _T_417;
        end
      end
    end
    if (reset) begin
      _T_267 <= 14'h0;
    end else begin
      if (_T_454) begin
        if (_T_306) begin
          _T_267 <= {{10'd0}, io_pixel_planar0_lp_burst};
        end else begin
          if (_T_309) begin
            _T_267 <= io_pixel_planar0_width_burst;
          end else begin
            if (_T_312) begin
              _T_267 <= io_pixel_planar0_width_burst;
            end else begin
              if (_T_315) begin
                _T_267 <= {{10'd0}, io_pixel_planar0_rp_burst};
              end else begin
                _T_267 <= _T_316;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_250 <= 4'h0;
    end else begin
      if (_T_454) begin
        if (_T_259) begin
          _T_250 <= io_pixel_planar0_bundle_limit_1st;
        end else begin
          if (_T_302) begin
            _T_250 <= io_pixel_planar0_bundle_limit;
          end else begin
            _T_250 <= _T_262;
          end
        end
      end
    end
    if (reset) begin
      _T_270 <= 2'h0;
    end else begin
      if (_T_458) begin
        if (_T_306) begin
          _T_270 <= 2'h0;
        end else begin
          if (_T_306) begin
            _T_270 <= 2'h1;
          end else begin
            _T_270 <= _T_329;
          end
        end
      end
    end
    if (reset) begin
      _T_337 <= 14'h0;
    end else begin
      if (_T_460) begin
        if (_T_388) begin
          _T_337 <= {{11'd0}, io_pixel_planar1_lp_burst};
        end else begin
          if (_T_391) begin
            _T_337 <= io_pixel_planar1_width_burst;
          end else begin
            if (_T_394) begin
              _T_337 <= io_pixel_planar1_width_burst;
            end else begin
              if (_T_397) begin
                _T_337 <= {{11'd0}, io_pixel_planar1_rp_burst};
              end else begin
                _T_337 <= _T_398;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_334 <= 5'h0;
    end else begin
      if (_T_460) begin
        if (_T_381) begin
          _T_334 <= io_pixel_planar1_bundle_limit_1st;
        end else begin
          if (_T_378) begin
            _T_334 <= io_pixel_planar1_bundle_limit;
          end else begin
            _T_334 <= _T_384;
          end
        end
      end
    end
    if (reset) begin
      _T_340 <= 2'h0;
    end else begin
      if (_T_463) begin
        if (_T_388) begin
          _T_340 <= 2'h0;
        end else begin
          if (_T_391) begin
            _T_340 <= 2'h1;
          end else begin
            _T_340 <= _T_412;
          end
        end
      end
    end
    if (reset) begin
      _T_480 <= 32'h0;
    end else begin
      if (_T_477) begin
        if (_T_171) begin
          _T_480 <= 32'h0;
        end else begin
          _T_480 <= _T_486;
        end
      end
    end
    if (reset) begin
      _T_483 <= 32'h0;
    end else begin
      if (_T_488) begin
        if (_T_171) begin
          _T_483 <= 32'h0;
        end else begin
          _T_483 <= _T_491;
        end
      end
    end
    if (reset) begin
      _T_495 <= 27'h0;
    end else begin
      if (_T_468) begin
        if (_T_259) begin
          _T_495 <= 27'h0;
        end else begin
          _T_495 <= _T_502;
        end
      end
    end
    if (reset) begin
      _T_498 <= 27'h0;
    end else begin
      if (_T_472) begin
        if (_T_381) begin
          _T_498 <= 27'h0;
        end else begin
          _T_498 <= _T_507;
        end
      end
    end
    if (io_layer_st) begin
      _T_510 <= _T_525;
    end
    if (io_layer_st) begin
      _T_512 <= _T_526;
    end
    if (reset) begin
      _T_529 <= 64'h0;
    end else begin
      if (_T_449) begin
        if (_T_240) begin
          _T_529 <= _T_524;
        end else begin
          _T_529 <= _T_518;
        end
      end
    end
    if (reset) begin
      _T_532 <= 5'h0;
    end else begin
      if (_T_449) begin
        if (_T_417) begin
          _T_532 <= {{1'd0}, _T_279};
        end else begin
          if (_T_354) begin
            _T_532 <= _T_352;
          end else begin
            _T_532 <= _T_334;
          end
        end
      end
    end
    if (reset) begin
      _T_535 <= 5'h0;
    end else begin
      if (_T_449) begin
        _T_535 <= _T_568;
      end
    end
    if (reset) begin
      _T_538 <= 1'h0;
    end else begin
      if (_T_449) begin
        if (_T_417) begin
          _T_538 <= _T_291;
        end else begin
          _T_538 <= _T_367;
        end
      end
    end
    if (reset) begin
      _T_541 <= 1'h0;
    end else begin
      if (_T_449) begin
        _T_541 <= _T_569;
      end
    end
    if (reset) begin
      _T_544 <= 1'h0;
    end else begin
      if (_T_449) begin
        _T_544 <= _T_450;
      end
    end
    if (reset) begin
      _T_547 <= 1'h0;
    end else begin
      if (_T_449) begin
        _T_547 <= _T_450;
      end
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      if (_T_449) begin
        _T_550 <= _T_451;
      end
    end
    if (reset) begin
      _T_553 <= 1'h0;
    end else begin
      if (_T_449) begin
        _T_553 <= _T_240;
      end
    end
    if (reset) begin
      _T_581 <= 1'h1;
    end else begin
      if (_T_171) begin
        _T_581 <= 1'h0;
      end else begin
        if (_T_587) begin
          _T_581 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_593 <= 1'h0;
    end else begin
      _T_593 <= _GEN_34[0];
    end
    if (reset) begin
      _T_674 <= 5'h0;
    end else begin
      if (_T_699) begin
        if (_T_695) begin
          _T_674 <= 5'h0;
        end else begin
          _T_674 <= _T_694;
        end
      end
    end
    if (reset) begin
      _T_710 <= 1'h0;
    end else begin
      if (_T_685) begin
        _T_710 <= 1'h0;
      end else begin
        if (_T_687) begin
          _T_710 <= _T_689;
        end else begin
          _T_710 <= 1'h1;
        end
      end
    end
    if (_T_692) begin
      _T_712 <= _T_1074;
    end
    if (reset) begin
      _T_1080 <= 1'h0;
    end else begin
      if (_T_699) begin
        _T_1080 <= _T_677;
      end
    end
    if (reset) begin
      _T_1083 <= 1'h0;
    end else begin
      if (_T_699) begin
        _T_1083 <= _T_1077;
      end
    end
    if (reset) begin
      _T_1086 <= 1'h0;
    end else begin
      if (_T_699) begin
        _T_1086 <= _T_701;
      end
    end
    if (reset) begin
      _T_1092 <= 5'h0;
    end else begin
      if (_T_1102) begin
        _T_1092 <= _T_683;
      end
    end
    if (reset) begin
      _T_1095 <= 1'h0;
    end else begin
      if (_T_699) begin
        _T_1095 <= _T_1103;
      end
    end
    if (reset) begin
      _T_1101 <= 1'h0;
    end else begin
      if (_T_699) begin
        _T_1101 <= _T_1105;
      end
    end
    if (reset) begin
      _T_1111 <= 256'h0;
    end else begin
      if (_T_1107) begin
        _T_1111 <= _T_712;
      end
    end
    if (reset) begin
      _T_1114 <= 256'h0;
    end else begin
      if (_T_1108) begin
        _T_1114 <= _T_712;
      end
    end
    if (reset) begin
      _T_1117 <= 1'h0;
    end else begin
      _T_1117 <= _T_1123;
    end
    if (_T_1123) begin
      _T_1119 <= _T_1129;
    end
    if (reset) begin
      _T_1134 <= 7'h0;
    end else begin
      if (_T_1151) begin
        if (_T_171) begin
          _T_1134 <= 7'h0;
        end else begin
          _T_1134 <= _T_1142;
        end
      end
    end
    if (reset) begin
      _T_1137 <= 7'h0;
    end else begin
      if (_T_1153) begin
        if (_T_171) begin
          _T_1137 <= 7'h0;
        end else begin
          _T_1137 <= _T_1144;
        end
      end
    end
    if (reset) begin
      _T_1140 <= 8'h0;
    end else begin
      if (_T_1123) begin
        if (_T_1106) begin
          _T_1140 <= _T_1159;
        end else begin
          _T_1140 <= _T_1164;
        end
      end
    end
    if (reset) begin
      _T_1168 <= 4'h0;
    end else begin
      if (_T_171) begin
        if (_T_171) begin
          _T_1168 <= 4'h0;
        end else begin
          if (_T_1106) begin
            _T_1168 <= _T_1192;
          end
        end
      end
    end
    if (reset) begin
      _T_1171 <= 5'h0;
    end else begin
      if (_T_171) begin
        if (_T_171) begin
          _T_1171 <= 5'h0;
        end else begin
          if (_T_1080) begin
            _T_1171 <= _T_1197;
          end
        end
      end
    end
    if (reset) begin
      _T_1174 <= 4'h0;
    end else begin
      if (_T_171) begin
        if (_T_1106) begin
          _T_1174 <= _T_1192;
        end else begin
          _T_1174 <= _T_1168;
        end
      end
    end
    if (reset) begin
      _T_1177 <= 5'h0;
    end else begin
      if (_T_171) begin
        _T_1177 <= _T_1197;
      end
    end
    if (reset) begin
      _T_1226 <= 1'h1;
    end else begin
      if (io_is_running) begin
        if (_T_171) begin
          _T_1226 <= 1'h0;
        end else begin
          if (_T_1228) begin
            _T_1226 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_1243 <= 1'h1;
    end else begin
      if (io_is_running) begin
        _T_1243 <= _T_1246;
      end
    end
    if (reset) begin
      _T_1252 <= 1'h0;
    end else begin
      _T_1252 <= _T_1249;
    end
    if (reset) begin
      _T_1256 <= 1'h0;
    end else begin
      _T_1256 <= _T_1253;
    end
    if (reset) begin
      _T_1260 <= 1'h0;
    end else begin
      _T_1260 <= _T_1257;
    end
    if (reset) begin
      _T_1267 <= 1'h0;
    end else begin
      _T_1267 <= _T_1249;
    end
    if (reset) begin
      _T_1273 <= 1'h0;
    end else begin
      _T_1273 <= _T_1270;
    end
    if (reset) begin
      _T_1276 <= 1'h0;
    end else begin
      _T_1276 <= io_status2dma_fsm_switch;
    end
    if (reset) begin
      _T_1280 <= 1'h0;
    end else begin
      _T_1280 <= _T_1257;
    end
  end
endmodule
module NV_NVDLA_CDMA_IMG_pack( // @[:@8470.2]
  input          reset, // @[:@8472.4]
  input          io_nvdla_core_clk, // @[:@8473.4]
  output         io_img2sbuf_p0_rd_addr_valid, // @[:@8473.4]
  output [7:0]   io_img2sbuf_p0_rd_addr_bits, // @[:@8473.4]
  input  [255:0] io_img2sbuf_p0_rd_data, // @[:@8473.4]
  input          io_is_running, // @[:@8473.4]
  input          io_layer_st, // @[:@8473.4]
  input  [5:0]   io_pixel_bank, // @[:@8473.4]
  input          io_pixel_early_end, // @[:@8473.4]
  input          io_pixel_packed_10b, // @[:@8473.4]
  input          io_pixel_planar, // @[:@8473.4]
  input  [2:0]   io_pixel_planar0_sft, // @[:@8473.4]
  input  [2:0]   io_pixel_planar1_sft, // @[:@8473.4]
  input  [1:0]   io_pixel_precision, // @[:@8473.4]
  input          io_pixel_uint, // @[:@8473.4]
  output         io_sg2pack_img_pd_ready, // @[:@8473.4]
  input          io_sg2pack_img_pd_valid, // @[:@8473.4]
  input  [10:0]  io_sg2pack_img_pd_bits, // @[:@8473.4]
  input  [14:0]  io_sg2pack_data_entries, // @[:@8473.4]
  input  [14:0]  io_sg2pack_entry_end, // @[:@8473.4]
  input  [14:0]  io_sg2pack_entry_mid, // @[:@8473.4]
  input  [14:0]  io_sg2pack_entry_st, // @[:@8473.4]
  input  [12:0]  io_sg2pack_height_total, // @[:@8473.4]
  input          io_sg2pack_mn_enable, // @[:@8473.4]
  input  [3:0]   io_sg2pack_sub_h_end, // @[:@8473.4]
  input  [3:0]   io_sg2pack_sub_h_mid, // @[:@8473.4]
  input  [3:0]   io_sg2pack_sub_h_st, // @[:@8473.4]
  input  [14:0]  io_status2dma_wr_idx, // @[:@8473.4]
  output         io_img2cvt_dat_wr_sel, // @[:@8473.4]
  output         io_img2cvt_dat_wr_addr_valid, // @[:@8473.4]
  output [16:0]  io_img2cvt_dat_wr_addr_bits, // @[:@8473.4]
  output [255:0] io_img2cvt_dat_wr_data, // @[:@8473.4]
  output [511:0] io_img2cvt_mn_wr_data, // @[:@8473.4]
  output [31:0]  io_img2cvt_dat_wr_pad_mask, // @[:@8473.4]
  output [11:0]  io_img2cvt_dat_wr_info_pd, // @[:@8473.4]
  output         io_img2status_dat_updt_valid, // @[:@8473.4]
  output [14:0]  io_img2status_dat_updt_bits_entries, // @[:@8473.4]
  output [13:0]  io_img2status_dat_updt_bits_slices, // @[:@8473.4]
  output         io_pack_is_done, // @[:@8473.4]
  input  [12:0]  io_reg2dp_datain_width, // @[:@8473.4]
  input  [12:0]  io_reg2dp_datain_channel, // @[:@8473.4]
  input  [15:0]  io_reg2dp_mean_ry, // @[:@8473.4]
  input  [15:0]  io_reg2dp_mean_gu, // @[:@8473.4]
  input  [15:0]  io_reg2dp_mean_bv, // @[:@8473.4]
  input  [15:0]  io_reg2dp_mean_ax, // @[:@8473.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@8473.4]
  input  [5:0]   io_reg2dp_pad_right // @[:@8473.4]
);
  reg  _T_115; // @[NV_NVDLA_CDMA_IMG_pack.scala 91:28:@8475.4]
  reg [31:0] _RAND_0;
  wire [10:0] _T_117; // @[NV_NVDLA_CDMA_IMG_pack.scala 93:17:@8476.4]
  wire [3:0] _T_118; // @[NV_NVDLA_CDMA_IMG_pack.scala 95:26:@8477.4]
  wire [4:0] _T_119; // @[NV_NVDLA_CDMA_IMG_pack.scala 96:26:@8478.4]
  wire  _T_120; // @[NV_NVDLA_CDMA_IMG_pack.scala 97:26:@8479.4]
  wire  _T_121; // @[NV_NVDLA_CDMA_IMG_pack.scala 98:27:@8480.4]
  wire  _T_122; // @[NV_NVDLA_CDMA_IMG_pack.scala 100:24:@8481.4]
  wire  _T_123; // @[NV_NVDLA_CDMA_IMG_pack.scala 100:39:@8482.4]
  reg [13:0] _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 106:32:@8484.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_129; // @[NV_NVDLA_CDMA_IMG_pack.scala 107:32:@8485.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_132; // @[NV_NVDLA_CDMA_IMG_pack.scala 108:32:@8486.4]
  reg [31:0] _RAND_3;
  wire [12:0] _GEN_82; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:45:@8489.6]
  wire [13:0] _T_133; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:45:@8489.6]
  wire [14:0] _T_135; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:71:@8490.6]
  wire [14:0] _GEN_84; // @[NV_NVDLA_CDMA_IMG_pack.scala 113:78:@8494.6]
  wire [15:0] _T_139; // @[NV_NVDLA_CDMA_IMG_pack.scala 113:78:@8494.6]
  wire [13:0] _GEN_0; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  wire [14:0] _GEN_1; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  wire [15:0] _GEN_2; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  reg [4:0] _T_142; // @[NV_NVDLA_CDMA_IMG_pack.scala 116:34:@8497.4]
  reg [31:0] _RAND_4;
  reg [4:0] _T_145; // @[NV_NVDLA_CDMA_IMG_pack.scala 117:34:@8498.4]
  reg [31:0] _RAND_5;
  reg [4:0] _T_148; // @[NV_NVDLA_CDMA_IMG_pack.scala 118:34:@8499.4]
  reg [31:0] _RAND_6;
  reg [4:0] _T_151; // @[NV_NVDLA_CDMA_IMG_pack.scala 119:34:@8500.4]
  reg [31:0] _RAND_7;
  reg [4:0] _T_154; // @[NV_NVDLA_CDMA_IMG_pack.scala 120:36:@8501.4]
  reg [31:0] _RAND_8;
  reg [4:0] _T_157; // @[NV_NVDLA_CDMA_IMG_pack.scala 121:36:@8502.4]
  reg [31:0] _RAND_9;
  reg [5:0] _T_160; // @[NV_NVDLA_CDMA_IMG_pack.scala 122:31:@8503.4]
  reg [31:0] _RAND_10;
  reg [5:0] _T_163; // @[NV_NVDLA_CDMA_IMG_pack.scala 123:31:@8504.4]
  reg [31:0] _RAND_11;
  wire [4:0] _T_164; // @[NV_NVDLA_CDMA_IMG_pack.scala 126:49:@8506.6]
  wire [9:0] _T_170; // @[Cat.scala 30:58:@8508.6]
  wire [9:0] _T_171; // @[NV_NVDLA_CDMA_IMG_pack.scala 126:97:@8509.6]
  wire [9:0] _T_179; // @[NV_NVDLA_CDMA_IMG_pack.scala 127:97:@8514.6]
  wire [4:0] _T_180; // @[NV_NVDLA_CDMA_IMG_pack.scala 128:49:@8516.6]
  wire [9:0] _T_186; // @[Cat.scala 30:58:@8518.6]
  wire [9:0] _T_187; // @[NV_NVDLA_CDMA_IMG_pack.scala 128:97:@8519.6]
  wire [9:0] _T_195; // @[NV_NVDLA_CDMA_IMG_pack.scala 129:97:@8524.6]
  wire [4:0] _T_196; // @[NV_NVDLA_CDMA_IMG_pack.scala 130:51:@8526.6]
  wire [9:0] _T_202; // @[Cat.scala 30:58:@8528.6]
  wire [9:0] _T_203; // @[NV_NVDLA_CDMA_IMG_pack.scala 130:99:@8529.6]
  wire [9:0] _T_211; // @[NV_NVDLA_CDMA_IMG_pack.scala 131:99:@8534.6]
  wire [7:0] _T_213; // @[NV_NVDLA_CDMA_IMG_pack.scala 132:29:@8536.6]
  wire [7:0] _T_215; // @[NV_NVDLA_CDMA_IMG_pack.scala 133:29:@8538.6]
  wire [9:0] _GEN_3; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [9:0] _GEN_4; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [9:0] _GEN_5; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [9:0] _GEN_6; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [9:0] _GEN_7; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [9:0] _GEN_8; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [7:0] _GEN_9; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  wire [7:0] _GEN_10; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  reg [12:0] _T_218; // @[NV_NVDLA_CDMA_IMG_pack.scala 139:28:@8541.4]
  reg [31:0] _RAND_12;
  wire  _T_222; // @[NV_NVDLA_CDMA_IMG_pack.scala 142:37:@8543.4]
  wire  _T_223; // @[NV_NVDLA_CDMA_IMG_pack.scala 142:21:@8544.4]
  wire  _T_224; // @[NV_NVDLA_CDMA_IMG_pack.scala 143:37:@8545.4]
  wire [13:0] _T_226; // @[NV_NVDLA_CDMA_IMG_pack.scala 144:39:@8546.4]
  wire [12:0] _T_227; // @[NV_NVDLA_CDMA_IMG_pack.scala 144:39:@8547.4]
  wire [12:0] _T_229; // @[NV_NVDLA_CDMA_IMG_pack.scala 145:26:@8548.4]
  reg  _T_281; // @[NV_NVDLA_CDMA_IMG_pack.scala 193:27:@8590.4]
  reg [31:0] _RAND_13;
  wire  _T_283; // @[NV_NVDLA_CDMA_IMG_pack.scala 196:36:@8593.4]
  reg [1:0] _T_257; // @[NV_NVDLA_CDMA_IMG_pack.scala 179:28:@8572.4]
  reg [31:0] _RAND_14;
  reg  _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 170:28:@8562.4]
  reg [31:0] _RAND_15;
  reg [3:0] _T_234; // @[NV_NVDLA_CDMA_IMG_pack.scala 157:26:@8552.4]
  reg [31:0] _RAND_16;
  wire [4:0] _T_238; // @[NV_NVDLA_CDMA_IMG_pack.scala 162:35:@8554.4]
  wire [3:0] _T_239; // @[NV_NVDLA_CDMA_IMG_pack.scala 162:35:@8555.4]
  wire  _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 163:37:@8556.4]
  wire  _T_260; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:45:@8574.4]
  wire  _T_261; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:74:@8575.4]
  wire  _T_262; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:61:@8576.4]
  wire  _T_263; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:59:@8577.4]
  wire  _T_264; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:42:@8578.4]
  wire [1:0] _T_267; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:26:@8579.4]
  wire  _T_268; // @[NV_NVDLA_CDMA_IMG_pack.scala 184:37:@8580.4]
  wire  _T_301; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:28:@8610.4]
  wire  _T_249; // @[NV_NVDLA_CDMA_IMG_pack.scala 172:22:@8564.4]
  wire  _T_250; // @[NV_NVDLA_CDMA_IMG_pack.scala 172:39:@8565.4]
  wire  _T_302; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:45:@8611.4]
  wire  _T_303; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:62:@8612.4]
  wire  _T_305; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:93:@8614.4]
  wire  _T_316; // @[NV_NVDLA_CDMA_IMG_pack.scala 210:38:@8628.4]
  wire [12:0] _GEN_11; // @[NV_NVDLA_CDMA_IMG_pack.scala 147:19:@8549.4]
  wire  _T_241; // @[NV_NVDLA_CDMA_IMG_pack.scala 166:41:@8558.6]
  wire [3:0] _T_243; // @[NV_NVDLA_CDMA_IMG_pack.scala 166:23:@8559.6]
  wire  _T_315; // @[NV_NVDLA_CDMA_IMG_pack.scala 209:38:@8626.4]
  wire [3:0] _GEN_12; // @[NV_NVDLA_CDMA_IMG_pack.scala 165:17:@8557.4]
  wire  _T_251; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:43:@8567.6]
  wire  _T_253; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:70:@8568.6]
  wire  _T_254; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:25:@8569.6]
  wire  _T_313; // @[NV_NVDLA_CDMA_IMG_pack.scala 208:55:@8623.4]
  wire  _T_314; // @[NV_NVDLA_CDMA_IMG_pack.scala 208:38:@8624.4]
  wire  _GEN_13; // @[NV_NVDLA_CDMA_IMG_pack.scala 174:19:@8566.4]
  wire  _T_269; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:43:@8582.6]
  wire [2:0] _T_272; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:93:@8583.6]
  wire [1:0] _T_273; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:93:@8584.6]
  wire [1:0] _T_274; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:25:@8585.6]
  wire  _T_312; // @[NV_NVDLA_CDMA_IMG_pack.scala 207:38:@8621.4]
  wire [1:0] _GEN_14; // @[NV_NVDLA_CDMA_IMG_pack.scala 186:19:@8581.4]
  wire  _T_284; // @[NV_NVDLA_CDMA_IMG_pack.scala 197:26:@8595.4]
  wire  _T_288; // @[NV_NVDLA_CDMA_IMG_pack.scala 199:25:@8596.4]
  wire  _T_289; // @[NV_NVDLA_CDMA_IMG_pack.scala 198:25:@8597.4]
  wire  _T_290; // @[NV_NVDLA_CDMA_IMG_pack.scala 197:25:@8598.4]
  wire  _T_311; // @[NV_NVDLA_CDMA_IMG_pack.scala 206:108:@8620.4]
  wire  _T_319; // @[NV_NVDLA_CDMA_IMG_pack.scala 212:52:@8632.4]
  wire  _T_320; // @[NV_NVDLA_CDMA_IMG_pack.scala 212:69:@8633.4]
  wire  _T_322; // @[NV_NVDLA_CDMA_IMG_pack.scala 213:52:@8635.4]
  wire  _T_323; // @[NV_NVDLA_CDMA_IMG_pack.scala 213:68:@8636.4]
  wire  _T_329; // @[NV_NVDLA_CDMA_IMG_pack.scala 215:99:@8642.4]
  wire  _T_334; // @[NV_NVDLA_CDMA_IMG_pack.scala 216:98:@8647.4]
  reg  _T_337; // @[NV_NVDLA_CDMA_IMG_pack.scala 219:24:@8649.4]
  reg [31:0] _RAND_17;
  reg  _T_354; // @[NV_NVDLA_CDMA_IMG_pack.scala 237:27:@8661.4]
  reg [31:0] _RAND_18;
  reg [6:0] _T_358; // @[NV_NVDLA_CDMA_IMG_pack.scala 242:32:@8665.4]
  reg [31:0] _RAND_19;
  reg [6:0] _T_361; // @[NV_NVDLA_CDMA_IMG_pack.scala 243:32:@8666.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_370; // @[NV_NVDLA_CDMA_IMG_pack.scala 246:25:@8669.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_373; // @[NV_NVDLA_CDMA_IMG_pack.scala 247:28:@8670.4]
  reg [31:0] _RAND_22;
  wire [7:0] _T_382; // @[NV_NVDLA_CDMA_IMG_pack.scala 254:47:@8675.4]
  wire [6:0] _T_383; // @[NV_NVDLA_CDMA_IMG_pack.scala 254:47:@8676.4]
  wire [7:0] _T_384; // @[NV_NVDLA_CDMA_IMG_pack.scala 255:47:@8677.4]
  wire [6:0] _T_385; // @[NV_NVDLA_CDMA_IMG_pack.scala 255:47:@8678.4]
  wire [6:0] _T_387; // @[NV_NVDLA_CDMA_IMG_pack.scala 256:30:@8679.4]
  wire [6:0] _T_389; // @[NV_NVDLA_CDMA_IMG_pack.scala 257:30:@8680.4]
  wire  _T_392; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:65:@8682.4]
  wire [5:0] _T_393; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:87:@8683.4]
  wire [7:0] _T_395; // @[Cat.scala 30:58:@8685.4]
  wire  _T_397; // @[NV_NVDLA_CDMA_IMG_pack.scala 259:43:@8686.4]
  wire [5:0] _T_398; // @[NV_NVDLA_CDMA_IMG_pack.scala 259:65:@8687.4]
  wire [7:0] _T_400; // @[Cat.scala 30:58:@8689.4]
  wire [7:0] _T_401; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:18:@8690.4]
  wire  _T_403; // @[NV_NVDLA_CDMA_IMG_pack.scala 279:45:@8708.4]
  wire  _T_404; // @[NV_NVDLA_CDMA_IMG_pack.scala 279:35:@8709.4]
  wire [6:0] _GEN_15; // @[NV_NVDLA_CDMA_IMG_pack.scala 262:20:@8692.4]
  wire  _T_405; // @[NV_NVDLA_CDMA_IMG_pack.scala 280:45:@8711.4]
  wire  _T_406; // @[NV_NVDLA_CDMA_IMG_pack.scala 280:35:@8712.4]
  wire [6:0] _GEN_16; // @[NV_NVDLA_CDMA_IMG_pack.scala 265:20:@8695.4]
  wire [7:0] _GEN_19; // @[NV_NVDLA_CDMA_IMG_pack.scala 274:16:@8704.4]
  reg [13:0] _T_409; // @[NV_NVDLA_CDMA_IMG_pack.scala 286:35:@8716.4]
  reg [31:0] _RAND_23;
  reg [13:0] _T_412; // @[NV_NVDLA_CDMA_IMG_pack.scala 287:35:@8717.4]
  reg [31:0] _RAND_24;
  wire [13:0] _GEN_85; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8718.4]
  wire [14:0] _T_413; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8718.4]
  wire [13:0] _T_414; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8719.4]
  wire [13:0] _GEN_86; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8720.4]
  wire [14:0] _T_415; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8720.4]
  wire [13:0] _T_416; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8721.4]
  wire  _T_417; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:57:@8722.4]
  wire  _T_418; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:98:@8723.4]
  wire  _T_419; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:139:@8724.4]
  wire [2:0] _T_421; // @[Cat.scala 30:58:@8726.4]
  wire  _T_422; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:57:@8727.4]
  wire  _T_423; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:98:@8728.4]
  wire  _T_424; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:139:@8729.4]
  wire [2:0] _T_426; // @[Cat.scala 30:58:@8731.4]
  wire  _T_431; // @[NV_NVDLA_CDMA_IMG_pack.scala 298:50:@8735.6]
  wire [13:0] _T_433; // @[NV_NVDLA_CDMA_IMG_pack.scala 298:32:@8736.6]
  wire [13:0] _GEN_20; // @[NV_NVDLA_CDMA_IMG_pack.scala 297:22:@8734.4]
  wire  _T_434; // @[NV_NVDLA_CDMA_IMG_pack.scala 301:50:@8740.6]
  wire [13:0] _T_436; // @[NV_NVDLA_CDMA_IMG_pack.scala 301:32:@8741.6]
  wire [13:0] _GEN_21; // @[NV_NVDLA_CDMA_IMG_pack.scala 300:22:@8739.4]
  reg [31:0] _T_450; // @[NV_NVDLA_CDMA_IMG_pack.scala 312:29:@8750.4]
  reg [31:0] _RAND_25;
  reg [31:0] _T_452; // @[NV_NVDLA_CDMA_IMG_pack.scala 313:28:@8751.4]
  reg [31:0] _RAND_26;
  wire [14:0] _T_453; // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8752.4]
  wire [14:0] _T_454; // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8753.4]
  wire [13:0] _T_455; // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8754.4]
  wire  _T_456; // @[NV_NVDLA_CDMA_IMG_pack.scala 317:57:@8755.4]
  wire  _T_457; // @[NV_NVDLA_CDMA_IMG_pack.scala 317:99:@8756.4]
  wire [1:0] _T_458; // @[Cat.scala 30:58:@8757.4]
  wire  _T_459; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:60:@8758.4]
  wire  _T_460; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:35:@8759.4]
  wire  _T_466; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:62:@8761.4]
  wire  _T_467; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:37:@8762.4]
  wire [286:0] _T_473; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:93:@8764.4]
  wire [286:0] _T_474; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:67:@8765.4]
  wire [286:0] _T_480; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:36:@8767.4]
  wire [286:0] _T_481; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:34:@8768.4]
  wire  _T_482; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:60:@8769.4]
  wire  _T_483; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:35:@8770.4]
  wire  _T_489; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:62:@8772.4]
  wire  _T_490; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:37:@8773.4]
  wire [286:0] _T_496; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:92:@8775.4]
  wire [286:0] _T_502; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:36:@8777.4]
  wire [286:0] _T_503; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:34:@8778.4]
  wire  _T_504; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:59:@8779.4]
  wire  _T_505; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:34:@8780.4]
  wire [286:0] _T_516; // @[NV_NVDLA_CDMA_IMG_pack.scala 325:58:@8783.4]
  wire [286:0] _T_517; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:33:@8784.4]
  wire [286:0] _T_518; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:55:@8786.4]
  wire [31:0] _T_438; // @[NV_NVDLA_CDMA_IMG_pack.scala 306:37:@8744.4 NV_NVDLA_CDMA_IMG_pack.scala 324:27:@8785.4]
  wire [31:0] _T_519; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:84:@8787.4]
  wire [286:0] _GEN_88; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:82:@8788.4]
  wire [286:0] _T_520; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:82:@8788.4]
  wire [14:0] _T_521; // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8790.4]
  wire [14:0] _T_522; // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8791.4]
  wire [13:0] _T_523; // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8792.4]
  wire  _T_524; // @[NV_NVDLA_CDMA_IMG_pack.scala 329:57:@8793.4]
  wire  _T_525; // @[NV_NVDLA_CDMA_IMG_pack.scala 329:99:@8794.4]
  wire [1:0] _T_526; // @[Cat.scala 30:58:@8795.4]
  wire  _T_527; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:60:@8796.4]
  wire  _T_528; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:35:@8797.4]
  wire  _T_534; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:62:@8799.4]
  wire  _T_535; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:37:@8800.4]
  wire [286:0] _T_541; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:93:@8802.4]
  wire [286:0] _T_542; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:67:@8803.4]
  wire [286:0] _T_548; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:36:@8805.4]
  wire [286:0] _T_549; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:34:@8806.4]
  wire  _T_550; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:60:@8807.4]
  wire  _T_551; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:35:@8808.4]
  wire  _T_557; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:62:@8810.4]
  wire  _T_558; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:37:@8811.4]
  wire [286:0] _T_564; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:92:@8813.4]
  wire [286:0] _T_570; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:36:@8815.4]
  wire [286:0] _T_571; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:34:@8816.4]
  wire  _T_572; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:59:@8817.4]
  wire  _T_573; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:34:@8818.4]
  wire [286:0] _T_584; // @[NV_NVDLA_CDMA_IMG_pack.scala 337:58:@8821.4]
  wire [286:0] _T_585; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:33:@8822.4]
  wire [286:0] _T_586; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:55:@8824.4]
  wire [31:0] _T_442; // @[NV_NVDLA_CDMA_IMG_pack.scala 308:37:@8746.4 NV_NVDLA_CDMA_IMG_pack.scala 336:27:@8823.4]
  wire [31:0] _T_587; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:84:@8825.4]
  wire [286:0] _GEN_90; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:82:@8826.4]
  wire [286:0] _T_588; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:82:@8826.4]
  wire [31:0] _T_440; // @[NV_NVDLA_CDMA_IMG_pack.scala 307:36:@8745.4 NV_NVDLA_CDMA_IMG_pack.scala 326:26:@8789.4]
  wire [31:0] _T_444; // @[NV_NVDLA_CDMA_IMG_pack.scala 309:36:@8747.4 NV_NVDLA_CDMA_IMG_pack.scala 338:26:@8827.4]
  wire [31:0] _T_590; // @[NV_NVDLA_CDMA_IMG_pack.scala 340:22:@8829.4]
  reg  _T_604; // @[NV_NVDLA_CDMA_IMG_pack.scala 351:27:@8849.4]
  reg [31:0] _RAND_27;
  reg [2:0] _T_607; // @[NV_NVDLA_CDMA_IMG_pack.scala 352:26:@8850.4]
  reg [31:0] _RAND_28;
  reg  _T_610; // @[NV_NVDLA_CDMA_IMG_pack.scala 353:30:@8851.4]
  reg [31:0] _RAND_29;
  reg  _T_613; // @[NV_NVDLA_CDMA_IMG_pack.scala 354:29:@8852.4]
  reg [31:0] _RAND_30;
  reg  _T_616; // @[NV_NVDLA_CDMA_IMG_pack.scala 355:33:@8853.4]
  reg [31:0] _RAND_31;
  reg  _T_619; // @[NV_NVDLA_CDMA_IMG_pack.scala 356:31:@8854.4]
  reg [31:0] _RAND_32;
  reg  _T_622; // @[NV_NVDLA_CDMA_IMG_pack.scala 357:30:@8855.4]
  reg [31:0] _RAND_33;
  wire  _T_623; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:41:@8861.6]
  wire  _T_624; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:58:@8862.6]
  wire  _T_625; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:73:@8863.6]
  wire  _T_626; // @[NV_NVDLA_CDMA_IMG_pack.scala 366:37:@8866.6]
  wire  _GEN_24; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire [2:0] _GEN_25; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire  _GEN_26; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire  _GEN_27; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire  _GEN_28; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire  _GEN_29; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  wire  _GEN_30; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  reg  _T_631; // @[NV_NVDLA_CDMA_IMG_pack.scala 380:59:@8872.4]
  reg [31:0] _RAND_34;
  reg  _T_634; // @[NV_NVDLA_CDMA_IMG_pack.scala 380:59:@8873.4]
  reg [31:0] _RAND_35;
  reg  _T_639; // @[NV_NVDLA_CDMA_IMG_pack.scala 382:62:@8875.4]
  reg [31:0] _RAND_36;
  reg  _T_642; // @[NV_NVDLA_CDMA_IMG_pack.scala 382:62:@8876.4]
  reg [31:0] _RAND_37;
  reg [2:0] _T_647; // @[NV_NVDLA_CDMA_IMG_pack.scala 384:62:@8878.4]
  reg [31:0] _RAND_38;
  reg [2:0] _T_650; // @[NV_NVDLA_CDMA_IMG_pack.scala 384:62:@8879.4]
  reg [31:0] _RAND_39;
  reg  _T_655; // @[NV_NVDLA_CDMA_IMG_pack.scala 386:59:@8881.4]
  reg [31:0] _RAND_40;
  reg  _T_658; // @[NV_NVDLA_CDMA_IMG_pack.scala 386:59:@8882.4]
  reg [31:0] _RAND_41;
  reg  _T_663; // @[NV_NVDLA_CDMA_IMG_pack.scala 388:62:@8884.4]
  reg [31:0] _RAND_42;
  reg  _T_666; // @[NV_NVDLA_CDMA_IMG_pack.scala 388:62:@8885.4]
  reg [31:0] _RAND_43;
  reg  _T_671; // @[NV_NVDLA_CDMA_IMG_pack.scala 390:59:@8887.4]
  reg [31:0] _RAND_44;
  reg  _T_674; // @[NV_NVDLA_CDMA_IMG_pack.scala 390:59:@8888.4]
  reg [31:0] _RAND_45;
  reg  _T_679; // @[NV_NVDLA_CDMA_IMG_pack.scala 392:62:@8890.4]
  reg [31:0] _RAND_46;
  reg  _T_682; // @[NV_NVDLA_CDMA_IMG_pack.scala 392:62:@8891.4]
  reg [31:0] _RAND_47;
  reg  _T_687; // @[NV_NVDLA_CDMA_IMG_pack.scala 394:59:@8893.4]
  reg [31:0] _RAND_48;
  reg  _T_690; // @[NV_NVDLA_CDMA_IMG_pack.scala 394:59:@8894.4]
  reg [31:0] _RAND_49;
  reg [31:0] _T_694; // @[NV_NVDLA_CDMA_IMG_pack.scala 397:64:@8896.4]
  reg [31:0] _RAND_50;
  reg [31:0] _T_696; // @[NV_NVDLA_CDMA_IMG_pack.scala 397:64:@8897.4]
  reg [31:0] _RAND_51;
  reg [31:0] _T_700; // @[NV_NVDLA_CDMA_IMG_pack.scala 399:64:@8899.4]
  reg [31:0] _RAND_52;
  reg [31:0] _T_702; // @[NV_NVDLA_CDMA_IMG_pack.scala 399:64:@8900.4]
  reg [31:0] _RAND_53;
  wire  _GEN_32; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire [2:0] _GEN_33; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_34; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_35; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_36; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_37; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_38; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  wire  _GEN_42; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire [2:0] _GEN_43; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _GEN_44; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _GEN_45; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _GEN_46; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _GEN_47; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _GEN_48; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  wire  _T_703; // @[NV_NVDLA_CDMA_IMG_pack.scala 437:43:@8937.4]
  wire  _T_704; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:34:@8938.4]
  wire  _T_705; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:54:@8939.4]
  wire  _T_706; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:52:@8940.4]
  reg  _T_709; // @[NV_NVDLA_CDMA_IMG_pack.scala 440:28:@8941.4]
  reg [31:0] _RAND_54;
  reg [2:0] _T_712; // @[NV_NVDLA_CDMA_IMG_pack.scala 441:30:@8942.4]
  reg [31:0] _RAND_55;
  reg  _T_715; // @[NV_NVDLA_CDMA_IMG_pack.scala 442:34:@8943.4]
  reg [31:0] _RAND_56;
  reg  _T_718; // @[NV_NVDLA_CDMA_IMG_pack.scala 443:33:@8944.4]
  reg [31:0] _RAND_57;
  reg  _T_721; // @[NV_NVDLA_CDMA_IMG_pack.scala 444:37:@8945.4]
  reg [31:0] _RAND_58;
  reg  _T_724; // @[NV_NVDLA_CDMA_IMG_pack.scala 445:35:@8946.4]
  reg [31:0] _RAND_59;
  reg  _T_727; // @[NV_NVDLA_CDMA_IMG_pack.scala 446:34:@8947.4]
  reg [31:0] _RAND_60;
  wire [2:0] _GEN_51; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  wire  _GEN_52; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  wire  _GEN_53; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  wire  _GEN_54; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  wire  _GEN_55; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  wire  _GEN_56; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  reg [1:0] _T_730; // @[NV_NVDLA_CDMA_IMG_pack.scala 466:28:@8957.4]
  reg [31:0] _RAND_61;
  wire  _T_732; // @[NV_NVDLA_CDMA_IMG_pack.scala 468:55:@8959.4]
  wire  _T_733; // @[NV_NVDLA_CDMA_IMG_pack.scala 468:41:@8960.4]
  wire  _T_734; // @[NV_NVDLA_CDMA_IMG_pack.scala 470:25:@8961.4]
  wire [2:0] _T_735; // @[NV_NVDLA_CDMA_IMG_pack.scala 471:27:@8962.4]
  wire  _T_736; // @[NV_NVDLA_CDMA_IMG_pack.scala 472:31:@8963.4]
  wire  _T_737; // @[NV_NVDLA_CDMA_IMG_pack.scala 473:30:@8964.4]
  wire  _T_738; // @[NV_NVDLA_CDMA_IMG_pack.scala 474:34:@8965.4]
  wire  _T_739; // @[NV_NVDLA_CDMA_IMG_pack.scala 475:32:@8966.4]
  wire  _T_740; // @[NV_NVDLA_CDMA_IMG_pack.scala 476:31:@8967.4]
  wire  _T_741; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:46:@8968.4]
  wire  _T_742; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:44:@8969.4]
  wire [2:0] _T_745; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:94:@8970.4]
  wire [1:0] _T_746; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:94:@8971.4]
  wire [1:0] _T_747; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:26:@8972.4]
  wire [1:0] _GEN_57; // @[NV_NVDLA_CDMA_IMG_pack.scala 481:17:@8973.4]
  reg  _T_758; // @[NV_NVDLA_CDMA_IMG_pack.scala 488:25:@8978.4]
  reg [31:0] _RAND_62;
  reg [2:0] _T_761; // @[NV_NVDLA_CDMA_IMG_pack.scala 489:27:@8979.4]
  reg [31:0] _RAND_63;
  reg [3:0] _T_764; // @[NV_NVDLA_CDMA_IMG_pack.scala 490:26:@8980.4]
  reg [31:0] _RAND_64;
  reg  _T_767; // @[NV_NVDLA_CDMA_IMG_pack.scala 491:26:@8981.4]
  reg [31:0] _RAND_65;
  reg  _T_770; // @[NV_NVDLA_CDMA_IMG_pack.scala 492:26:@8982.4]
  reg [31:0] _RAND_66;
  wire [2:0] _GEN_58; // @[NV_NVDLA_CDMA_IMG_pack.scala 495:20:@8984.4]
  wire [3:0] _GEN_59; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  wire  _GEN_60; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  wire  _GEN_61; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  wire [5:0] _T_775; // @[Cat.scala 30:58:@8993.4]
  wire [5:0] _T_778; // @[Cat.scala 30:58:@8996.4]
  reg [255:0] _T_782; // @[NV_NVDLA_CDMA_IMG_pack.scala 509:35:@8998.4]
  reg [255:0] _RAND_67;
  reg [255:0] _T_785; // @[NV_NVDLA_CDMA_IMG_pack.scala 510:35:@8999.4]
  reg [255:0] _RAND_68;
  reg [255:0] _T_788; // @[NV_NVDLA_CDMA_IMG_pack.scala 511:35:@9000.4]
  reg [255:0] _RAND_69;
  reg [31:0] _T_791; // @[NV_NVDLA_CDMA_IMG_pack.scala 512:37:@9001.4]
  reg [31:0] _RAND_70;
  reg [31:0] _T_794; // @[NV_NVDLA_CDMA_IMG_pack.scala 513:37:@9002.4]
  reg [31:0] _RAND_71;
  reg [31:0] _T_797; // @[NV_NVDLA_CDMA_IMG_pack.scala 514:37:@9003.4]
  reg [31:0] _RAND_72;
  reg [255:0] _T_799; // @[NV_NVDLA_CDMA_IMG_pack.scala 515:25:@9004.4]
  reg [255:0] _RAND_73;
  reg [31:0] _T_802; // @[NV_NVDLA_CDMA_IMG_pack.scala 516:33:@9005.4]
  reg [31:0] _RAND_74;
  wire  _T_813; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9014.4]
  wire  _T_814; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9015.4]
  wire  _T_815; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9016.4]
  wire  _T_816; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9017.4]
  wire [7:0] _T_818; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9018.4]
  wire [7:0] _T_819; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9019.4]
  wire  _T_820; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9020.4]
  wire  _T_821; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9021.4]
  wire  _T_822; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9022.4]
  wire  _T_823; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9023.4]
  wire [7:0] _T_825; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9024.4]
  wire [7:0] _T_826; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9025.4]
  wire  _T_827; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9026.4]
  wire  _T_828; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9027.4]
  wire  _T_829; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9028.4]
  wire  _T_830; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9029.4]
  wire [7:0] _T_832; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9030.4]
  wire [7:0] _T_833; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9031.4]
  wire  _T_834; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9032.4]
  wire  _T_835; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9033.4]
  wire  _T_836; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9034.4]
  wire  _T_837; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9035.4]
  wire [7:0] _T_839; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9036.4]
  wire [7:0] _T_840; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9037.4]
  wire  _T_841; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9038.4]
  wire  _T_842; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9039.4]
  wire  _T_843; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9040.4]
  wire  _T_844; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9041.4]
  wire [7:0] _T_846; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9042.4]
  wire [7:0] _T_847; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9043.4]
  wire  _T_848; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9044.4]
  wire  _T_849; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9045.4]
  wire  _T_850; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9046.4]
  wire  _T_851; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9047.4]
  wire [7:0] _T_853; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9048.4]
  wire [7:0] _T_854; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9049.4]
  wire  _T_855; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9050.4]
  wire  _T_856; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9051.4]
  wire  _T_857; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9052.4]
  wire  _T_858; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9053.4]
  wire [7:0] _T_860; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9054.4]
  wire [7:0] _T_861; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9055.4]
  wire  _T_862; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9056.4]
  wire  _T_863; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9057.4]
  wire  _T_864; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9058.4]
  wire  _T_865; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9059.4]
  wire [7:0] _T_867; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9060.4]
  wire [7:0] _T_868; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9061.4]
  wire  _T_869; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9062.4]
  wire  _T_870; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9063.4]
  wire  _T_871; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9064.4]
  wire  _T_872; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9065.4]
  wire [7:0] _T_874; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9066.4]
  wire [7:0] _T_875; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9067.4]
  wire  _T_876; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9068.4]
  wire  _T_877; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9069.4]
  wire  _T_878; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9070.4]
  wire  _T_879; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9071.4]
  wire [7:0] _T_881; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9072.4]
  wire [7:0] _T_882; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9073.4]
  wire  _T_883; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9074.4]
  wire  _T_884; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9075.4]
  wire  _T_885; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9076.4]
  wire  _T_886; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9077.4]
  wire [7:0] _T_888; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9078.4]
  wire [7:0] _T_889; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9079.4]
  wire  _T_890; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9080.4]
  wire  _T_891; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9081.4]
  wire  _T_892; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9082.4]
  wire  _T_893; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9083.4]
  wire [7:0] _T_895; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9084.4]
  wire [7:0] _T_896; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9085.4]
  wire  _T_897; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9086.4]
  wire  _T_898; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9087.4]
  wire  _T_899; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9088.4]
  wire  _T_900; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9089.4]
  wire [7:0] _T_902; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9090.4]
  wire [7:0] _T_903; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9091.4]
  wire  _T_904; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9092.4]
  wire  _T_905; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9093.4]
  wire  _T_906; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9094.4]
  wire  _T_907; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9095.4]
  wire [7:0] _T_909; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9096.4]
  wire [7:0] _T_910; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9097.4]
  wire  _T_911; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9098.4]
  wire  _T_912; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9099.4]
  wire  _T_913; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9100.4]
  wire  _T_914; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9101.4]
  wire [7:0] _T_916; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9102.4]
  wire [7:0] _T_917; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9103.4]
  wire  _T_918; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9104.4]
  wire  _T_919; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9105.4]
  wire  _T_920; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9106.4]
  wire  _T_921; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9107.4]
  wire [7:0] _T_923; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9108.4]
  wire [7:0] _T_924; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9109.4]
  wire  _T_925; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9110.4]
  wire  _T_926; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9111.4]
  wire  _T_927; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9112.4]
  wire  _T_928; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9113.4]
  wire [7:0] _T_930; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9114.4]
  wire [7:0] _T_931; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9115.4]
  wire  _T_932; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9116.4]
  wire  _T_933; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9117.4]
  wire  _T_934; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9118.4]
  wire  _T_935; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9119.4]
  wire [7:0] _T_937; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9120.4]
  wire [7:0] _T_938; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9121.4]
  wire  _T_939; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9122.4]
  wire  _T_940; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9123.4]
  wire  _T_941; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9124.4]
  wire  _T_942; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9125.4]
  wire [7:0] _T_944; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9126.4]
  wire [7:0] _T_945; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9127.4]
  wire  _T_946; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9128.4]
  wire  _T_947; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9129.4]
  wire  _T_948; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9130.4]
  wire  _T_949; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9131.4]
  wire [7:0] _T_951; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9132.4]
  wire [7:0] _T_952; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9133.4]
  wire  _T_953; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9134.4]
  wire  _T_954; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9135.4]
  wire  _T_955; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9136.4]
  wire  _T_956; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9137.4]
  wire [7:0] _T_958; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9138.4]
  wire [7:0] _T_959; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9139.4]
  wire  _T_960; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9140.4]
  wire  _T_961; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9141.4]
  wire  _T_962; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9142.4]
  wire  _T_963; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9143.4]
  wire [7:0] _T_965; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9144.4]
  wire [7:0] _T_966; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9145.4]
  wire  _T_967; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9146.4]
  wire  _T_968; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9147.4]
  wire  _T_969; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9148.4]
  wire  _T_970; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9149.4]
  wire [7:0] _T_972; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9150.4]
  wire [7:0] _T_973; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9151.4]
  wire  _T_974; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9152.4]
  wire  _T_975; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9153.4]
  wire  _T_976; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9154.4]
  wire  _T_977; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9155.4]
  wire [7:0] _T_979; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9156.4]
  wire [7:0] _T_980; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9157.4]
  wire  _T_981; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9158.4]
  wire  _T_982; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9159.4]
  wire  _T_983; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9160.4]
  wire  _T_984; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9161.4]
  wire [7:0] _T_986; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9162.4]
  wire [7:0] _T_987; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9163.4]
  wire  _T_988; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9164.4]
  wire  _T_989; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9165.4]
  wire  _T_990; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9166.4]
  wire  _T_991; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9167.4]
  wire [7:0] _T_993; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9168.4]
  wire [7:0] _T_994; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9169.4]
  wire  _T_995; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9170.4]
  wire  _T_996; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9171.4]
  wire  _T_997; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9172.4]
  wire  _T_998; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9173.4]
  wire [7:0] _T_1000; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9174.4]
  wire [7:0] _T_1001; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9175.4]
  wire  _T_1002; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9176.4]
  wire  _T_1003; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9177.4]
  wire  _T_1004; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9178.4]
  wire  _T_1005; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9179.4]
  wire [7:0] _T_1007; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9180.4]
  wire [7:0] _T_1008; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9181.4]
  wire  _T_1009; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9182.4]
  wire  _T_1010; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9183.4]
  wire  _T_1011; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9184.4]
  wire  _T_1012; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9185.4]
  wire [7:0] _T_1014; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9186.4]
  wire [7:0] _T_1015; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9187.4]
  wire  _T_1016; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9188.4]
  wire  _T_1017; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9189.4]
  wire  _T_1018; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9190.4]
  wire  _T_1019; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9191.4]
  wire [7:0] _T_1021; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9192.4]
  wire [7:0] _T_1022; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9193.4]
  wire  _T_1023; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9194.4]
  wire  _T_1024; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9195.4]
  wire  _T_1025; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9196.4]
  wire  _T_1026; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9197.4]
  wire [7:0] _T_1028; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9198.4]
  wire [7:0] _T_1029; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9199.4]
  wire  _T_1030; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9200.4]
  wire  _T_1031; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9201.4]
  wire  _T_1032; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9202.4]
  wire  _T_1033; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9203.4]
  wire [7:0] _T_1035; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9204.4]
  wire [7:0] _T_1036; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9205.4]
  wire [63:0] _T_1081; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9245.4]
  wire [127:0] _T_1089; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9253.4]
  wire [63:0] _T_1096; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9260.4]
  wire [255:0] _T_1105; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9269.4]
  wire  _T_1522; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:54:@9657.4]
  wire  _T_1524; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:87:@9658.4]
  wire  _T_1525; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:70:@9659.4]
  wire [255:0] _T_1106; // @[NV_NVDLA_CDMA_IMG_pack.scala 533:20:@9270.4]
  wire  _T_1529; // @[NV_NVDLA_CDMA_IMG_pack.scala 560:87:@9663.4]
  wire  _T_1530; // @[NV_NVDLA_CDMA_IMG_pack.scala 560:70:@9664.4]
  wire [255:0] _T_1107; // @[NV_NVDLA_CDMA_IMG_pack.scala 534:20:@9271.4]
  wire [511:0] _T_1108; // @[Cat.scala 30:58:@9272.4]
  wire [15:0] _T_1109; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9273.4]
  wire [7:0] _T_1110; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9274.4]
  wire [15:0] _T_1112; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9276.4]
  wire [7:0] _T_1113; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9277.4]
  wire [15:0] _T_1115; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9279.4]
  wire [7:0] _T_1116; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9280.4]
  wire [15:0] _T_1118; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9282.4]
  wire [7:0] _T_1119; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9283.4]
  wire [15:0] _T_1121; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9285.4]
  wire [7:0] _T_1122; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9286.4]
  wire [15:0] _T_1124; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9288.4]
  wire [7:0] _T_1125; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9289.4]
  wire [15:0] _T_1127; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9291.4]
  wire [7:0] _T_1128; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9292.4]
  wire [15:0] _T_1130; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9294.4]
  wire [7:0] _T_1131; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9295.4]
  wire [15:0] _T_1133; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9297.4]
  wire [7:0] _T_1134; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9298.4]
  wire [15:0] _T_1136; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9300.4]
  wire [7:0] _T_1137; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9301.4]
  wire [15:0] _T_1139; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9303.4]
  wire [7:0] _T_1140; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9304.4]
  wire [15:0] _T_1142; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9306.4]
  wire [7:0] _T_1143; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9307.4]
  wire [15:0] _T_1145; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9309.4]
  wire [7:0] _T_1146; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9310.4]
  wire [15:0] _T_1148; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9312.4]
  wire [7:0] _T_1149; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9313.4]
  wire [15:0] _T_1151; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9315.4]
  wire [7:0] _T_1152; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9316.4]
  wire [15:0] _T_1154; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9318.4]
  wire [7:0] _T_1155; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9319.4]
  wire [15:0] _T_1157; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9321.4]
  wire [7:0] _T_1158; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9322.4]
  wire [15:0] _T_1160; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9324.4]
  wire [7:0] _T_1161; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9325.4]
  wire [15:0] _T_1163; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9327.4]
  wire [7:0] _T_1164; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9328.4]
  wire [15:0] _T_1166; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9330.4]
  wire [7:0] _T_1167; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9331.4]
  wire [15:0] _T_1169; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9333.4]
  wire [7:0] _T_1170; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9334.4]
  wire [15:0] _T_1172; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9336.4]
  wire [7:0] _T_1173; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9337.4]
  wire [15:0] _T_1175; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9339.4]
  wire [7:0] _T_1176; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9340.4]
  wire [15:0] _T_1178; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9342.4]
  wire [7:0] _T_1179; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9343.4]
  wire [15:0] _T_1181; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9345.4]
  wire [7:0] _T_1182; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9346.4]
  wire [15:0] _T_1184; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9348.4]
  wire [7:0] _T_1185; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9349.4]
  wire [15:0] _T_1187; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9351.4]
  wire [7:0] _T_1188; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9352.4]
  wire [15:0] _T_1190; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9354.4]
  wire [7:0] _T_1191; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9355.4]
  wire [15:0] _T_1193; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9357.4]
  wire [7:0] _T_1194; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9358.4]
  wire [15:0] _T_1196; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9360.4]
  wire [7:0] _T_1197; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9361.4]
  wire [15:0] _T_1199; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9363.4]
  wire [7:0] _T_1200; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9364.4]
  wire [15:0] _T_1202; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9366.4]
  wire [7:0] _T_1203; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9367.4]
  wire [95:0] _T_1245; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9404.4]
  wire [191:0] _T_1249; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9408.4]
  wire [95:0] _T_1252; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9411.4]
  wire [383:0] _T_1257; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9416.4]
  wire [95:0] _T_1260; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9419.4]
  wire [191:0] _T_1264; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9423.4]
  wire [95:0] _T_1267; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9426.4]
  wire [383:0] _T_1272; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9431.4]
  wire [767:0] _T_1273; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9432.4]
  wire  _T_1275; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:59:@9433.4]
  wire  _T_1276; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:42:@9434.4]
  wire  _T_1279; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:85:@9436.4]
  wire  _T_1282; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:41:@9438.4]
  wire  _T_1284; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:87:@9440.4]
  wire  _T_1285; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:85:@9441.4]
  wire [4:0] _T_1289; // @[Cat.scala 30:58:@9445.4]
  wire  _T_1290; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:68:@9446.4]
  wire [255:0] _T_1294; // @[Bitwise.scala 72:12:@9448.4]
  wire [255:0] _T_1295; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:73:@9449.4]
  wire  _T_1296; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:68:@9450.4]
  wire [255:0] _T_1300; // @[Bitwise.scala 72:12:@9452.4]
  wire [255:0] _T_1301; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:82:@9453.4]
  wire [255:0] _T_1302; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:73:@9454.4]
  wire [255:0] _T_1303; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:93:@9455.4]
  wire  _T_1304; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:68:@9456.4]
  wire [255:0] _T_1308; // @[Bitwise.scala 72:12:@9458.4]
  wire [255:0] _T_1309; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:82:@9459.4]
  wire [255:0] _T_1310; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:73:@9460.4]
  wire [255:0] _T_1311; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:115:@9461.4]
  wire  _T_1312; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:68:@9462.4]
  wire [255:0] _T_1316; // @[Bitwise.scala 72:12:@9464.4]
  wire [255:0] _T_1317; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:82:@9465.4]
  wire [255:0] _T_1318; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:73:@9466.4]
  wire [255:0] _T_1319; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:139:@9467.4]
  wire [31:0] _T_1320; // @[NV_NVDLA_CDMA_IMG_pack.scala 548:25:@9468.4]
  wire [31:0] _T_1321; // @[NV_NVDLA_CDMA_IMG_pack.scala 549:25:@9469.4]
  wire [63:0] _T_1322; // @[Cat.scala 30:58:@9470.4]
  wire [1:0] _T_1323; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9471.4]
  wire  _T_1324; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9472.4]
  wire [1:0] _T_1326; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9474.4]
  wire  _T_1327; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9475.4]
  wire [1:0] _T_1329; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9477.4]
  wire  _T_1330; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9478.4]
  wire [1:0] _T_1332; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9480.4]
  wire  _T_1333; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9481.4]
  wire [1:0] _T_1335; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9483.4]
  wire  _T_1336; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9484.4]
  wire [1:0] _T_1338; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9486.4]
  wire  _T_1339; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9487.4]
  wire [1:0] _T_1341; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9489.4]
  wire  _T_1342; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9490.4]
  wire [1:0] _T_1344; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9492.4]
  wire  _T_1345; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9493.4]
  wire [1:0] _T_1347; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9495.4]
  wire  _T_1348; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9496.4]
  wire [1:0] _T_1350; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9498.4]
  wire  _T_1351; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9499.4]
  wire [1:0] _T_1353; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9501.4]
  wire  _T_1354; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9502.4]
  wire [1:0] _T_1356; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9504.4]
  wire  _T_1357; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9505.4]
  wire [1:0] _T_1359; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9507.4]
  wire  _T_1360; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9508.4]
  wire [1:0] _T_1362; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9510.4]
  wire  _T_1363; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9511.4]
  wire [1:0] _T_1365; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9513.4]
  wire  _T_1366; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9514.4]
  wire [1:0] _T_1368; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9516.4]
  wire  _T_1369; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9517.4]
  wire [1:0] _T_1371; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9519.4]
  wire  _T_1372; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9520.4]
  wire [1:0] _T_1374; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9522.4]
  wire  _T_1375; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9523.4]
  wire [1:0] _T_1377; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9525.4]
  wire  _T_1378; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9526.4]
  wire [1:0] _T_1380; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9528.4]
  wire  _T_1381; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9529.4]
  wire [1:0] _T_1383; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9531.4]
  wire  _T_1384; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9532.4]
  wire [1:0] _T_1386; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9534.4]
  wire  _T_1387; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9535.4]
  wire [1:0] _T_1389; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9537.4]
  wire  _T_1390; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9538.4]
  wire [1:0] _T_1392; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9540.4]
  wire  _T_1393; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9541.4]
  wire [1:0] _T_1395; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9543.4]
  wire  _T_1396; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9544.4]
  wire [1:0] _T_1398; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9546.4]
  wire  _T_1399; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9547.4]
  wire [1:0] _T_1401; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9549.4]
  wire  _T_1402; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9550.4]
  wire [1:0] _T_1404; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9552.4]
  wire  _T_1405; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9553.4]
  wire [1:0] _T_1407; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9555.4]
  wire  _T_1408; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9556.4]
  wire [1:0] _T_1410; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9558.4]
  wire  _T_1411; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9559.4]
  wire [1:0] _T_1413; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9561.4]
  wire  _T_1414; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9562.4]
  wire [1:0] _T_1416; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9564.4]
  wire  _T_1417; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9565.4]
  wire [11:0] _T_1459; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9602.4]
  wire [23:0] _T_1463; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9606.4]
  wire [11:0] _T_1466; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9609.4]
  wire [47:0] _T_1471; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9614.4]
  wire [11:0] _T_1474; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9617.4]
  wire [23:0] _T_1478; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9621.4]
  wire [11:0] _T_1481; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9624.4]
  wire [47:0] _T_1486; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9629.4]
  wire [95:0] _T_1487; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9630.4]
  wire [31:0] _T_1492; // @[Bitwise.scala 72:12:@9633.4]
  wire [31:0] _T_1493; // @[NV_NVDLA_CDMA_IMG_pack.scala 554:92:@9634.4]
  wire [31:0] _T_1498; // @[Bitwise.scala 72:12:@9637.4]
  wire [31:0] _T_1499; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:102:@9638.4]
  wire [31:0] _T_1500; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:88:@9639.4]
  wire [31:0] _T_1501; // @[NV_NVDLA_CDMA_IMG_pack.scala 554:116:@9640.4]
  wire [31:0] _T_1506; // @[Bitwise.scala 72:12:@9643.4]
  wire [31:0] _T_1507; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:102:@9644.4]
  wire [31:0] _T_1508; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:88:@9645.4]
  wire [31:0] _T_1509; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:150:@9646.4]
  wire [31:0] _T_1514; // @[Bitwise.scala 72:12:@9649.4]
  wire [31:0] _T_1515; // @[NV_NVDLA_CDMA_IMG_pack.scala 557:102:@9650.4]
  wire [31:0] _T_1516; // @[NV_NVDLA_CDMA_IMG_pack.scala 557:88:@9651.4]
  wire [31:0] _T_1517; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:189:@9652.4]
  wire  _T_1520; // @[NV_NVDLA_CDMA_IMG_pack.scala 558:58:@9655.4]
  wire [255:0] _GEN_62; // @[NV_NVDLA_CDMA_IMG_pack.scala 563:27:@9666.4]
  wire [31:0] _GEN_63; // @[NV_NVDLA_CDMA_IMG_pack.scala 563:27:@9666.4]
  wire [31:0] _GEN_69; // @[NV_NVDLA_CDMA_IMG_pack.scala 575:24:@9678.4]
  reg [255:0] _T_1542; // @[NV_NVDLA_CDMA_IMG_pack.scala 587:32:@9685.4]
  reg [255:0] _RAND_75;
  wire [127:0] _T_1717; // @[Cat.scala 30:58:@9853.4]
  wire [255:0] _T_1718; // @[Cat.scala 30:58:@9854.4]
  wire [511:0] _T_1719; // @[Cat.scala 30:58:@9855.4]
  wire [127:0] _T_1723; // @[Cat.scala 30:58:@9859.4]
  wire [255:0] _T_1724; // @[Cat.scala 30:58:@9860.4]
  wire [511:0] _T_1725; // @[Cat.scala 30:58:@9861.4]
  wire [95:0] _T_1728; // @[Cat.scala 30:58:@9864.4]
  wire [191:0] _T_1729; // @[Cat.scala 30:58:@9865.4]
  wire [383:0] _T_1730; // @[Cat.scala 30:58:@9866.4]
  wire [767:0] _T_1731; // @[Cat.scala 30:58:@9867.4]
  wire [1535:0] _T_1732; // @[Cat.scala 30:58:@9868.4]
  wire  _T_1734; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:47:@9869.4]
  wire  _T_1735; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:20:@9870.4]
  wire [511:0] _T_1736; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:19:@9871.4]
  wire [15:0] _T_1739; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9873.4]
  wire [15:0] _T_1740; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9874.4]
  wire [15:0] _T_1743; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9876.4]
  wire [15:0] _T_1744; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9877.4]
  wire [15:0] _T_1747; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9879.4]
  wire [15:0] _T_1748; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9880.4]
  wire [15:0] _T_1751; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9882.4]
  wire [15:0] _T_1752; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9883.4]
  wire [15:0] _T_1755; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9885.4]
  wire [15:0] _T_1756; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9886.4]
  wire [15:0] _T_1759; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9888.4]
  wire [15:0] _T_1760; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9889.4]
  wire [15:0] _T_1763; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9891.4]
  wire [15:0] _T_1764; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9892.4]
  wire [15:0] _T_1767; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9894.4]
  wire [15:0] _T_1768; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9895.4]
  wire [15:0] _T_1771; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9897.4]
  wire [15:0] _T_1772; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9898.4]
  wire [15:0] _T_1775; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9900.4]
  wire [15:0] _T_1776; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9901.4]
  wire [15:0] _T_1779; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9903.4]
  wire [15:0] _T_1780; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9904.4]
  wire [15:0] _T_1783; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9906.4]
  wire [15:0] _T_1784; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9907.4]
  wire [15:0] _T_1787; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9909.4]
  wire [15:0] _T_1788; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9910.4]
  wire [15:0] _T_1791; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9912.4]
  wire [15:0] _T_1792; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9913.4]
  wire [15:0] _T_1795; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9915.4]
  wire [15:0] _T_1796; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9916.4]
  wire [15:0] _T_1799; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9918.4]
  wire [15:0] _T_1800; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9919.4]
  wire [15:0] _T_1803; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9921.4]
  wire [15:0] _T_1804; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9922.4]
  wire [15:0] _T_1807; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9924.4]
  wire [15:0] _T_1808; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9925.4]
  wire [15:0] _T_1811; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9927.4]
  wire [15:0] _T_1812; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9928.4]
  wire [15:0] _T_1815; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9930.4]
  wire [15:0] _T_1816; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9931.4]
  wire [15:0] _T_1819; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9933.4]
  wire [15:0] _T_1820; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9934.4]
  wire [15:0] _T_1823; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9936.4]
  wire [15:0] _T_1824; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9937.4]
  wire [15:0] _T_1827; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9939.4]
  wire [15:0] _T_1828; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9940.4]
  wire [15:0] _T_1831; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9942.4]
  wire [15:0] _T_1832; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9943.4]
  wire [15:0] _T_1835; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9945.4]
  wire [15:0] _T_1836; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9946.4]
  wire [15:0] _T_1839; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9948.4]
  wire [15:0] _T_1840; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9949.4]
  wire [15:0] _T_1843; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9951.4]
  wire [15:0] _T_1844; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9952.4]
  wire [15:0] _T_1847; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9954.4]
  wire [15:0] _T_1848; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9955.4]
  wire [15:0] _T_1851; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9957.4]
  wire [15:0] _T_1852; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9958.4]
  wire [15:0] _T_1855; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9960.4]
  wire [15:0] _T_1856; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9961.4]
  wire [15:0] _T_1859; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9963.4]
  wire [15:0] _T_1860; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9964.4]
  wire [15:0] _T_1863; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9966.4]
  wire [15:0] _T_1864; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9967.4]
  wire [127:0] _T_1909; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10007.4]
  wire [255:0] _T_1917; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10015.4]
  wire [127:0] _T_1924; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10022.4]
  wire [511:0] _T_1933; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10031.4]
  wire  _T_1934; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10032.4]
  wire [15:0] _T_1936; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10033.4]
  wire [15:0] _T_1937; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10034.4]
  wire  _T_1938; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10035.4]
  wire [15:0] _T_1940; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10036.4]
  wire [15:0] _T_1941; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10037.4]
  wire  _T_1942; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10038.4]
  wire [15:0] _T_1944; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10039.4]
  wire [15:0] _T_1945; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10040.4]
  wire  _T_1946; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10041.4]
  wire [15:0] _T_1948; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10042.4]
  wire [15:0] _T_1949; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10043.4]
  wire  _T_1950; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10044.4]
  wire [15:0] _T_1952; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10045.4]
  wire [15:0] _T_1953; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10046.4]
  wire  _T_1954; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10047.4]
  wire [15:0] _T_1956; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10048.4]
  wire [15:0] _T_1957; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10049.4]
  wire  _T_1958; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10050.4]
  wire [15:0] _T_1960; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10051.4]
  wire [15:0] _T_1961; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10052.4]
  wire  _T_1962; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10053.4]
  wire [15:0] _T_1964; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10054.4]
  wire [15:0] _T_1965; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10055.4]
  wire  _T_1966; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10056.4]
  wire [15:0] _T_1968; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10057.4]
  wire [15:0] _T_1969; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10058.4]
  wire  _T_1970; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10059.4]
  wire [15:0] _T_1972; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10060.4]
  wire [15:0] _T_1973; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10061.4]
  wire  _T_1974; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10062.4]
  wire [15:0] _T_1976; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10063.4]
  wire [15:0] _T_1977; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10064.4]
  wire  _T_1978; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10065.4]
  wire [15:0] _T_1980; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10066.4]
  wire [15:0] _T_1981; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10067.4]
  wire  _T_1982; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10068.4]
  wire [15:0] _T_1984; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10069.4]
  wire [15:0] _T_1985; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10070.4]
  wire  _T_1986; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10071.4]
  wire [15:0] _T_1988; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10072.4]
  wire [15:0] _T_1989; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10073.4]
  wire  _T_1990; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10074.4]
  wire [15:0] _T_1992; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10075.4]
  wire [15:0] _T_1993; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10076.4]
  wire  _T_1994; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10077.4]
  wire [15:0] _T_1996; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10078.4]
  wire [15:0] _T_1997; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10079.4]
  wire  _T_1998; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10080.4]
  wire [15:0] _T_2000; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10081.4]
  wire [15:0] _T_2001; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10082.4]
  wire  _T_2002; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10083.4]
  wire [15:0] _T_2004; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10084.4]
  wire [15:0] _T_2005; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10085.4]
  wire  _T_2006; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10086.4]
  wire [15:0] _T_2008; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10087.4]
  wire [15:0] _T_2009; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10088.4]
  wire  _T_2010; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10089.4]
  wire [15:0] _T_2012; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10090.4]
  wire [15:0] _T_2013; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10091.4]
  wire  _T_2014; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10092.4]
  wire [15:0] _T_2016; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10093.4]
  wire [15:0] _T_2017; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10094.4]
  wire  _T_2018; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10095.4]
  wire [15:0] _T_2020; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10096.4]
  wire [15:0] _T_2021; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10097.4]
  wire  _T_2022; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10098.4]
  wire [15:0] _T_2024; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10099.4]
  wire [15:0] _T_2025; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10100.4]
  wire  _T_2026; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10101.4]
  wire [15:0] _T_2028; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10102.4]
  wire [15:0] _T_2029; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10103.4]
  wire  _T_2030; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10104.4]
  wire [15:0] _T_2032; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10105.4]
  wire [15:0] _T_2033; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10106.4]
  wire  _T_2034; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10107.4]
  wire [15:0] _T_2036; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10108.4]
  wire [15:0] _T_2037; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10109.4]
  wire  _T_2038; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10110.4]
  wire [15:0] _T_2040; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10111.4]
  wire [15:0] _T_2041; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10112.4]
  wire  _T_2042; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10113.4]
  wire [15:0] _T_2044; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10114.4]
  wire [15:0] _T_2045; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10115.4]
  wire  _T_2046; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10116.4]
  wire [15:0] _T_2048; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10117.4]
  wire [15:0] _T_2049; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10118.4]
  wire  _T_2050; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10119.4]
  wire [15:0] _T_2052; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10120.4]
  wire [15:0] _T_2053; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10121.4]
  wire  _T_2054; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10122.4]
  wire [15:0] _T_2056; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10123.4]
  wire [15:0] _T_2057; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10124.4]
  wire  _T_2058; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10125.4]
  wire [15:0] _T_2060; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10126.4]
  wire [15:0] _T_2061; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10127.4]
  wire  _T_2062; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10128.4]
  wire [15:0] _T_2064; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10129.4]
  wire [15:0] _T_2065; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10130.4]
  wire  _T_2066; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10131.4]
  wire [15:0] _T_2068; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10132.4]
  wire [15:0] _T_2069; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10133.4]
  wire  _T_2070; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10134.4]
  wire [15:0] _T_2072; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10135.4]
  wire [15:0] _T_2073; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10136.4]
  wire  _T_2074; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10137.4]
  wire [15:0] _T_2076; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10138.4]
  wire [15:0] _T_2077; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10139.4]
  wire  _T_2078; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10140.4]
  wire [15:0] _T_2080; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10141.4]
  wire [15:0] _T_2081; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10142.4]
  wire  _T_2082; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10143.4]
  wire [15:0] _T_2084; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10144.4]
  wire [15:0] _T_2085; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10145.4]
  wire  _T_2086; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10146.4]
  wire [15:0] _T_2088; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10147.4]
  wire [15:0] _T_2089; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10148.4]
  wire  _T_2090; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10149.4]
  wire [15:0] _T_2092; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10150.4]
  wire [15:0] _T_2093; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10151.4]
  wire  _T_2094; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10152.4]
  wire [15:0] _T_2096; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10153.4]
  wire [15:0] _T_2097; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10154.4]
  wire  _T_2098; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10155.4]
  wire [15:0] _T_2100; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10156.4]
  wire [15:0] _T_2101; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10157.4]
  wire  _T_2102; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10158.4]
  wire [15:0] _T_2104; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10159.4]
  wire [15:0] _T_2105; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10160.4]
  wire  _T_2106; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10161.4]
  wire [15:0] _T_2108; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10162.4]
  wire [15:0] _T_2109; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10163.4]
  wire  _T_2110; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10164.4]
  wire [15:0] _T_2112; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10165.4]
  wire [15:0] _T_2113; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10166.4]
  wire  _T_2114; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10167.4]
  wire [15:0] _T_2116; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10168.4]
  wire [15:0] _T_2117; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10169.4]
  wire  _T_2118; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10170.4]
  wire [15:0] _T_2120; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10171.4]
  wire [15:0] _T_2121; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10172.4]
  wire  _T_2122; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10173.4]
  wire [15:0] _T_2124; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10174.4]
  wire [15:0] _T_2125; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10175.4]
  wire  _T_2126; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10176.4]
  wire [15:0] _T_2128; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10177.4]
  wire [15:0] _T_2129; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10178.4]
  wire  _T_2130; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10179.4]
  wire [15:0] _T_2132; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10180.4]
  wire [15:0] _T_2133; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10181.4]
  wire  _T_2134; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10182.4]
  wire [15:0] _T_2136; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10183.4]
  wire [15:0] _T_2137; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10184.4]
  wire  _T_2138; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10185.4]
  wire [15:0] _T_2140; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10186.4]
  wire [15:0] _T_2141; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10187.4]
  wire  _T_2142; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10188.4]
  wire [15:0] _T_2144; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10189.4]
  wire [15:0] _T_2145; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10190.4]
  wire  _T_2146; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10191.4]
  wire [15:0] _T_2148; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10192.4]
  wire [15:0] _T_2149; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10193.4]
  wire  _T_2150; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10194.4]
  wire [15:0] _T_2152; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10195.4]
  wire [15:0] _T_2153; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10196.4]
  wire  _T_2154; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10197.4]
  wire [15:0] _T_2156; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10198.4]
  wire [15:0] _T_2157; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10199.4]
  wire  _T_2158; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10200.4]
  wire [15:0] _T_2160; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10201.4]
  wire [15:0] _T_2161; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10202.4]
  wire  _T_2162; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10203.4]
  wire [15:0] _T_2164; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10204.4]
  wire [15:0] _T_2165; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10205.4]
  wire  _T_2166; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10206.4]
  wire [15:0] _T_2168; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10207.4]
  wire [15:0] _T_2169; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10208.4]
  wire  _T_2170; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10209.4]
  wire [15:0] _T_2172; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10210.4]
  wire [15:0] _T_2173; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10211.4]
  wire  _T_2174; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10212.4]
  wire [15:0] _T_2176; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10213.4]
  wire [15:0] _T_2177; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10214.4]
  wire  _T_2178; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10215.4]
  wire [15:0] _T_2180; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10216.4]
  wire [15:0] _T_2181; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10217.4]
  wire  _T_2182; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10218.4]
  wire [15:0] _T_2184; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10219.4]
  wire [15:0] _T_2185; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10220.4]
  wire  _T_2186; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10221.4]
  wire [15:0] _T_2188; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10222.4]
  wire [15:0] _T_2189; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10223.4]
  wire  _T_2190; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10224.4]
  wire [15:0] _T_2192; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10225.4]
  wire [15:0] _T_2193; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10226.4]
  wire  _T_2194; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10227.4]
  wire [15:0] _T_2196; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10228.4]
  wire [15:0] _T_2197; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10229.4]
  wire  _T_2198; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10230.4]
  wire [15:0] _T_2200; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10231.4]
  wire [15:0] _T_2201; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10232.4]
  wire  _T_2202; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10233.4]
  wire [15:0] _T_2204; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10234.4]
  wire [15:0] _T_2205; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10235.4]
  wire  _T_2206; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10236.4]
  wire [15:0] _T_2208; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10237.4]
  wire [15:0] _T_2209; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10238.4]
  wire  _T_2210; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10239.4]
  wire [15:0] _T_2212; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10240.4]
  wire [15:0] _T_2213; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10241.4]
  wire  _T_2214; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10242.4]
  wire [15:0] _T_2216; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10243.4]
  wire [15:0] _T_2217; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10244.4]
  wire  _T_2218; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10245.4]
  wire [15:0] _T_2220; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10246.4]
  wire [15:0] _T_2221; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10247.4]
  wire  _T_2222; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10248.4]
  wire [15:0] _T_2224; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10249.4]
  wire [15:0] _T_2225; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10250.4]
  wire  _T_2226; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10251.4]
  wire [15:0] _T_2228; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10252.4]
  wire [15:0] _T_2229; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10253.4]
  wire  _T_2230; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10254.4]
  wire [15:0] _T_2232; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10255.4]
  wire [15:0] _T_2233; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10256.4]
  wire  _T_2234; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10257.4]
  wire [15:0] _T_2236; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10258.4]
  wire [15:0] _T_2237; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10259.4]
  wire  _T_2238; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10260.4]
  wire [15:0] _T_2240; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10261.4]
  wire [15:0] _T_2241; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10262.4]
  wire  _T_2242; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10263.4]
  wire [15:0] _T_2244; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10264.4]
  wire [15:0] _T_2245; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10265.4]
  wire  _T_2246; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10266.4]
  wire [15:0] _T_2248; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10267.4]
  wire [15:0] _T_2249; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10268.4]
  wire  _T_2250; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10269.4]
  wire [15:0] _T_2252; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10270.4]
  wire [15:0] _T_2253; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10271.4]
  wire  _T_2254; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10272.4]
  wire [15:0] _T_2256; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10273.4]
  wire [15:0] _T_2257; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10274.4]
  wire  _T_2258; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10275.4]
  wire [15:0] _T_2260; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10276.4]
  wire [15:0] _T_2261; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10277.4]
  wire  _T_2262; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10278.4]
  wire [15:0] _T_2264; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10279.4]
  wire [15:0] _T_2265; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10280.4]
  wire  _T_2266; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10281.4]
  wire [15:0] _T_2268; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10282.4]
  wire [15:0] _T_2269; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10283.4]
  wire  _T_2270; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10284.4]
  wire [15:0] _T_2272; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10285.4]
  wire [15:0] _T_2273; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10286.4]
  wire  _T_2274; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10287.4]
  wire [15:0] _T_2276; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10288.4]
  wire [15:0] _T_2277; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10289.4]
  wire  _T_2278; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10290.4]
  wire [15:0] _T_2280; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10291.4]
  wire [15:0] _T_2281; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10292.4]
  wire  _T_2282; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10293.4]
  wire [15:0] _T_2284; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10294.4]
  wire [15:0] _T_2285; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10295.4]
  wire  _T_2286; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10296.4]
  wire [15:0] _T_2288; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10297.4]
  wire [15:0] _T_2289; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10298.4]
  wire  _T_2290; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10299.4]
  wire [15:0] _T_2292; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10300.4]
  wire [15:0] _T_2293; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10301.4]
  wire  _T_2294; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10302.4]
  wire [15:0] _T_2296; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10303.4]
  wire [15:0] _T_2297; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10304.4]
  wire  _T_2298; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10305.4]
  wire [15:0] _T_2300; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10306.4]
  wire [15:0] _T_2301; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10307.4]
  wire  _T_2302; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10308.4]
  wire [15:0] _T_2304; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10309.4]
  wire [15:0] _T_2305; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10310.4]
  wire  _T_2306; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10311.4]
  wire [15:0] _T_2308; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10312.4]
  wire [15:0] _T_2309; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10313.4]
  wire  _T_2310; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10314.4]
  wire [15:0] _T_2312; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10315.4]
  wire [15:0] _T_2313; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10316.4]
  wire  _T_2314; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10317.4]
  wire [15:0] _T_2316; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10318.4]
  wire [15:0] _T_2317; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10319.4]
  wire [95:0] _T_2424; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10421.4]
  wire [191:0] _T_2430; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10427.4]
  wire [95:0] _T_2435; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10432.4]
  wire [383:0] _T_2442; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10439.4]
  wire [95:0] _T_2447; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10444.4]
  wire [191:0] _T_2453; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10450.4]
  wire [95:0] _T_2458; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10455.4]
  wire [767:0] _T_2466; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10463.4]
  wire [95:0] _T_2471; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10468.4]
  wire [191:0] _T_2477; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10474.4]
  wire [95:0] _T_2482; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10479.4]
  wire [383:0] _T_2489; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10486.4]
  wire [95:0] _T_2494; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10491.4]
  wire [191:0] _T_2500; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10497.4]
  wire [95:0] _T_2505; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10502.4]
  wire [1535:0] _T_2514; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10511.4]
  wire  _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 606:87:@10514.4]
  wire  _T_2520; // @[NV_NVDLA_CDMA_IMG_pack.scala 606:66:@10515.4]
  wire  _T_2526; // @[NV_NVDLA_CDMA_IMG_pack.scala 607:68:@10519.4]
  wire  _T_2527; // @[NV_NVDLA_CDMA_IMG_pack.scala 607:66:@10520.4]
  wire  _T_2533; // @[NV_NVDLA_CDMA_IMG_pack.scala 608:66:@10524.4]
  wire  _T_2540; // @[NV_NVDLA_CDMA_IMG_pack.scala 609:66:@10529.4]
  wire  _T_2546; // @[NV_NVDLA_CDMA_IMG_pack.scala 610:66:@10533.4]
  wire  _T_2553; // @[NV_NVDLA_CDMA_IMG_pack.scala 611:66:@10538.4]
  wire  _T_2559; // @[NV_NVDLA_CDMA_IMG_pack.scala 612:65:@10543.4]
  wire  _T_2564; // @[NV_NVDLA_CDMA_IMG_pack.scala 613:65:@10547.4]
  wire  _T_2565; // @[NV_NVDLA_CDMA_IMG_pack.scala 613:42:@10548.4]
  wire [7:0] _T_2572; // @[Cat.scala 30:58:@10555.4]
  wire  _T_2573; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:56:@10556.4]
  wire [511:0] _T_2577; // @[Bitwise.scala 72:12:@10558.4]
  wire [511:0] _T_2578; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:60:@10559.4]
  wire  _T_2579; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:56:@10560.4]
  wire [511:0] _T_2583; // @[Bitwise.scala 72:12:@10562.4]
  wire [511:0] _T_2584; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:71:@10563.4]
  wire [511:0] _T_2585; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:60:@10564.4]
  wire [511:0] _T_2586; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:73:@10565.4]
  wire  _T_2587; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:56:@10566.4]
  wire [511:0] _T_2591; // @[Bitwise.scala 72:12:@10568.4]
  wire [511:0] _T_2592; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:71:@10569.4]
  wire [511:0] _T_2593; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:60:@10570.4]
  wire [511:0] _T_2594; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:89:@10571.4]
  wire  _T_2595; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:56:@10572.4]
  wire [511:0] _T_2599; // @[Bitwise.scala 72:12:@10574.4]
  wire [511:0] _T_2600; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:71:@10575.4]
  wire [511:0] _T_2601; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:60:@10576.4]
  wire [511:0] _T_2602; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:100:@10577.4]
  wire  _T_2606; // @[NV_NVDLA_CDMA_IMG_pack.scala 623:72:@10582.4]
  wire  _T_2607; // @[NV_NVDLA_CDMA_IMG_pack.scala 623:43:@10583.4]
  wire [511:0] _GEN_73; // @[NV_NVDLA_CDMA_IMG_pack.scala 634:27:@10593.4]
  reg [14:0] _T_2610; // @[NV_NVDLA_CDMA_IMG_pack.scala 644:29:@10596.4]
  reg [31:0] _RAND_76;
  wire [14:0] _T_2611; // @[NV_NVDLA_CDMA_IMG_pack.scala 647:28:@10597.4]
  wire [14:0] _T_2612; // @[NV_NVDLA_CDMA_IMG_pack.scala 646:28:@10598.4]
  wire [3:0] _T_2613; // @[NV_NVDLA_CDMA_IMG_pack.scala 649:28:@10599.4]
  wire [3:0] _T_2614; // @[NV_NVDLA_CDMA_IMG_pack.scala 648:27:@10600.4]
  wire [15:0] _T_2616; // @[Cat.scala 30:58:@10601.4]
  wire [15:0] _T_2617; // @[NV_NVDLA_CDMA_IMG_pack.scala 650:99:@10602.4]
  wire [15:0] _T_2618; // @[NV_NVDLA_CDMA_IMG_pack.scala 650:29:@10603.4]
  wire [6:0] _T_2619; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:38:@10604.4]
  wire [6:0] _GEN_91; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:76:@10605.4]
  wire  _T_2620; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:76:@10605.4]
  wire [14:0] _T_2627; // @[Cat.scala 30:58:@10608.4]
  wire [15:0] _GEN_92; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10609.4]
  wire [16:0] _T_2628; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10609.4]
  wire [16:0] _T_2629; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10610.4]
  wire [14:0] _T_2630; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:124:@10611.4]
  wire [14:0] _T_2631; // @[NV_NVDLA_CDMA_IMG_pack.scala 654:81:@10612.4]
  wire [14:0] _T_2632; // @[NV_NVDLA_CDMA_IMG_pack.scala 654:27:@10613.4]
  wire  _T_2633; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:59:@10614.4]
  wire  _T_2634; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:85:@10615.4]
  wire  _T_2635; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:42:@10616.4]
  wire [14:0] _GEN_74; // @[NV_NVDLA_CDMA_IMG_pack.scala 658:24:@10617.4]
  reg [14:0] _T_2638; // @[NV_NVDLA_CDMA_IMG_pack.scala 663:33:@10620.4]
  reg [31:0] _RAND_77;
  wire  _T_2639; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:49:@10621.4]
  wire [15:0] _T_2641; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:111:@10622.4]
  wire [14:0] _T_2642; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:111:@10623.4]
  wire [14:0] _T_2643; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:31:@10624.4]
  wire  _T_2644; // @[NV_NVDLA_CDMA_IMG_pack.scala 666:63:@10625.4]
  wire  _T_2645; // @[NV_NVDLA_CDMA_IMG_pack.scala 666:46:@10626.4]
  wire [14:0] _GEN_75; // @[NV_NVDLA_CDMA_IMG_pack.scala 668:28:@10627.4]
  reg [14:0] _T_2648; // @[NV_NVDLA_CDMA_IMG_pack.scala 672:33:@10630.4]
  reg [31:0] _RAND_78;
  reg [14:0] _T_2651; // @[NV_NVDLA_CDMA_IMG_pack.scala 673:37:@10631.4]
  reg [31:0] _RAND_79;
  wire  _T_2652; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:77:@10632.4]
  wire  _T_2653; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:50:@10633.4]
  wire  _T_2655; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:54:@10634.4]
  wire  _T_2656; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:52:@10635.4]
  wire [15:0] _T_2657; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:120:@10636.4]
  wire [14:0] _T_2658; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:120:@10637.4]
  wire [14:0] _T_2659; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:31:@10638.4]
  wire [14:0] _T_2660; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:31:@10639.4]
  wire  _T_2661; // @[NV_NVDLA_CDMA_IMG_pack.scala 679:46:@10640.4]
  wire [14:0] _GEN_76; // @[NV_NVDLA_CDMA_IMG_pack.scala 682:28:@10641.4]
  wire [14:0] _GEN_77; // @[NV_NVDLA_CDMA_IMG_pack.scala 685:32:@10644.4]
  reg  _T_2664; // @[NV_NVDLA_CDMA_IMG_pack.scala 689:26:@10647.4]
  reg [31:0] _RAND_80;
  wire [15:0] _T_2665; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:41:@10648.4]
  wire [13:0] _T_2666; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:84:@10649.4]
  wire [15:0] _GEN_93; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:63:@10650.4]
  wire [16:0] _T_2667; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:63:@10650.4]
  wire  _T_2668; // @[NV_NVDLA_CDMA_IMG_pack.scala 692:63:@10651.4]
  wire  _GEN_78; // @[NV_NVDLA_CDMA_IMG_pack.scala 697:32:@10652.4]
  reg [14:0] _T_2672; // @[NV_NVDLA_CDMA_IMG_pack.scala 710:26:@10656.4]
  reg [31:0] _RAND_81;
  wire [7:0] _T_2673; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:38:@10657.4]
  wire [7:0] _GEN_94; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:76:@10658.4]
  wire  _T_2674; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:76:@10658.4]
  wire [16:0] _GEN_95; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10662.4]
  wire [17:0] _T_2682; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10662.4]
  wire [17:0] _T_2683; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10663.4]
  wire [14:0] _T_2684; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:124:@10664.4]
  wire [14:0] _T_2685; // @[NV_NVDLA_CDMA_IMG_pack.scala 714:79:@10665.4]
  wire [14:0] _T_2686; // @[NV_NVDLA_CDMA_IMG_pack.scala 714:25:@10666.4]
  wire [14:0] _GEN_79; // @[NV_NVDLA_CDMA_IMG_pack.scala 717:20:@10667.4]
  reg  _T_2689; // @[NV_NVDLA_CDMA_IMG_pack.scala 724:31:@10670.4]
  reg [31:0] _RAND_82;
  reg [14:0] _T_2692; // @[NV_NVDLA_CDMA_IMG_pack.scala 725:34:@10671.4]
  reg [31:0] _RAND_83;
  reg [3:0] _T_2695; // @[NV_NVDLA_CDMA_IMG_pack.scala 726:33:@10672.4]
  reg [31:0] _RAND_84;
  wire [14:0] _GEN_80; // @[NV_NVDLA_CDMA_IMG_pack.scala 731:23:@10676.4]
  wire [3:0] _GEN_81; // @[NV_NVDLA_CDMA_IMG_pack.scala 731:23:@10676.4]
  reg  _T_2702; // @[NV_NVDLA_CDMA_IMG_pack.scala 757:31:@10691.4]
  reg [31:0] _RAND_85;
  wire  _T_2704; // @[NV_NVDLA_CDMA_IMG_pack.scala 760:40:@10692.4]
  wire  _T_2706; // @[NV_NVDLA_CDMA_IMG_pack.scala 760:25:@10693.4]
  wire  _T_2707; // @[NV_NVDLA_CDMA_IMG_pack.scala 759:25:@10694.4]
  assign _T_117 = io_sg2pack_img_pd_valid ? io_sg2pack_img_pd_bits : 11'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 93:17:@8476.4]
  assign _T_118 = _T_117[3:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 95:26:@8477.4]
  assign _T_119 = _T_117[8:4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 96:26:@8478.4]
  assign _T_120 = _T_117[9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 97:26:@8479.4]
  assign _T_121 = _T_117[10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 98:27:@8480.4]
  assign _T_122 = ~ _T_115; // @[NV_NVDLA_CDMA_IMG_pack.scala 100:24:@8481.4]
  assign _T_123 = _T_122 & io_is_running; // @[NV_NVDLA_CDMA_IMG_pack.scala 100:39:@8482.4]
  assign _GEN_82 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:45:@8489.6]
  assign _T_133 = _GEN_82 + io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:45:@8489.6]
  assign _T_135 = _T_133 + 14'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 112:71:@8490.6]
  assign _GEN_84 = {{9'd0}, io_reg2dp_pad_right}; // @[NV_NVDLA_CDMA_IMG_pack.scala 113:78:@8494.6]
  assign _T_139 = _T_135 + _GEN_84; // @[NV_NVDLA_CDMA_IMG_pack.scala 113:78:@8494.6]
  assign _GEN_0 = io_layer_st ? {{9'd0}, io_reg2dp_pad_left} : _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  assign _GEN_1 = io_layer_st ? _T_135 : {{1'd0}, _T_129}; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  assign _GEN_2 = io_layer_st ? _T_139 : {{2'd0}, _T_132}; // @[NV_NVDLA_CDMA_IMG_pack.scala 110:18:@8487.4]
  assign _T_164 = _T_126[4:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 126:49:@8506.6]
  assign _T_170 = {_T_164,5'h0}; // @[Cat.scala 30:58:@8508.6]
  assign _T_171 = _T_170 >> io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 126:97:@8509.6]
  assign _T_179 = _T_170 >> io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 127:97:@8514.6]
  assign _T_180 = _T_129[4:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 128:49:@8516.6]
  assign _T_186 = {_T_180,5'h0}; // @[Cat.scala 30:58:@8518.6]
  assign _T_187 = _T_186 >> io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 128:97:@8519.6]
  assign _T_195 = _T_186 >> io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 129:97:@8524.6]
  assign _T_196 = _T_132[4:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 130:51:@8526.6]
  assign _T_202 = {_T_196,5'h0}; // @[Cat.scala 30:58:@8528.6]
  assign _T_203 = _T_202 >> io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 130:99:@8529.6]
  assign _T_211 = _T_202 >> io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 131:99:@8534.6]
  assign _T_213 = 8'h1 << io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 132:29:@8536.6]
  assign _T_215 = 8'h1 << io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_IMG_pack.scala 133:29:@8538.6]
  assign _GEN_3 = _T_123 ? _T_171 : {{5'd0}, _T_142}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_4 = _T_123 ? _T_179 : {{5'd0}, _T_145}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_5 = _T_123 ? _T_187 : {{5'd0}, _T_148}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_6 = _T_123 ? _T_195 : {{5'd0}, _T_151}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_7 = _T_123 ? _T_203 : {{5'd0}, _T_154}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_8 = _T_123 ? _T_211 : {{5'd0}, _T_157}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_9 = _T_123 ? _T_213 : {{2'd0}, _T_160}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _GEN_10 = _T_123 ? _T_215 : {{2'd0}, _T_163}; // @[NV_NVDLA_CDMA_IMG_pack.scala 125:23:@8505.4]
  assign _T_222 = _T_218 != 13'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 142:37:@8543.4]
  assign _T_223 = ~ _T_222; // @[NV_NVDLA_CDMA_IMG_pack.scala 142:21:@8544.4]
  assign _T_224 = _T_218 == io_sg2pack_height_total; // @[NV_NVDLA_CDMA_IMG_pack.scala 143:37:@8545.4]
  assign _T_226 = _T_218 + 13'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 144:39:@8546.4]
  assign _T_227 = _T_218 + 13'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 144:39:@8547.4]
  assign _T_229 = _T_123 ? 13'h0 : _T_227; // @[NV_NVDLA_CDMA_IMG_pack.scala 145:26:@8548.4]
  assign _T_283 = io_sg2pack_img_pd_valid | _T_281; // @[NV_NVDLA_CDMA_IMG_pack.scala 196:36:@8593.4]
  assign _T_238 = _T_234 + 4'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 162:35:@8554.4]
  assign _T_239 = _T_234 + 4'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 162:35:@8555.4]
  assign _T_240 = _T_239 >= _T_118; // @[NV_NVDLA_CDMA_IMG_pack.scala 163:37:@8556.4]
  assign _T_260 = ~ _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:45:@8574.4]
  assign _T_261 = _T_119[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:74:@8575.4]
  assign _T_262 = ~ _T_261; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:61:@8576.4]
  assign _T_263 = _T_260 | _T_262; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:59:@8577.4]
  assign _T_264 = _T_246 & _T_263; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:42:@8578.4]
  assign _T_267 = _T_264 ? 2'h1 : 2'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 182:26:@8579.4]
  assign _T_268 = _T_257 == _T_267; // @[NV_NVDLA_CDMA_IMG_pack.scala 184:37:@8580.4]
  assign _T_301 = _T_283 & _T_268; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:28:@8610.4]
  assign _T_249 = ~ io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_pack.scala 172:22:@8564.4]
  assign _T_250 = _T_249 | _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 172:39:@8565.4]
  assign _T_302 = _T_301 & _T_250; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:45:@8611.4]
  assign _T_303 = _T_302 & _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:62:@8612.4]
  assign _T_305 = _T_303 & _T_120; // @[NV_NVDLA_CDMA_IMG_pack.scala 205:93:@8614.4]
  assign _T_316 = _T_123 | _T_305; // @[NV_NVDLA_CDMA_IMG_pack.scala 210:38:@8628.4]
  assign _GEN_11 = _T_316 ? _T_229 : _T_218; // @[NV_NVDLA_CDMA_IMG_pack.scala 147:19:@8549.4]
  assign _T_241 = _T_123 | _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 166:41:@8558.6]
  assign _T_243 = _T_241 ? 4'h0 : _T_239; // @[NV_NVDLA_CDMA_IMG_pack.scala 166:23:@8559.6]
  assign _T_315 = _T_123 | _T_302; // @[NV_NVDLA_CDMA_IMG_pack.scala 209:38:@8626.4]
  assign _GEN_12 = _T_315 ? _T_243 : _T_234; // @[NV_NVDLA_CDMA_IMG_pack.scala 165:17:@8557.4]
  assign _T_251 = _T_123 | _T_250; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:43:@8567.6]
  assign _T_253 = ~ _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:70:@8568.6]
  assign _T_254 = _T_251 ? 1'h0 : _T_253; // @[NV_NVDLA_CDMA_IMG_pack.scala 175:25:@8569.6]
  assign _T_313 = _T_301 & io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_pack.scala 208:55:@8623.4]
  assign _T_314 = _T_123 | _T_313; // @[NV_NVDLA_CDMA_IMG_pack.scala 208:38:@8624.4]
  assign _GEN_13 = _T_314 ? _T_254 : _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 174:19:@8566.4]
  assign _T_269 = _T_123 | _T_268; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:43:@8582.6]
  assign _T_272 = _T_257 + 2'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:93:@8583.6]
  assign _T_273 = _T_257 + 2'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:93:@8584.6]
  assign _T_274 = _T_269 ? 2'h0 : _T_273; // @[NV_NVDLA_CDMA_IMG_pack.scala 187:25:@8585.6]
  assign _T_312 = _T_123 | _T_283; // @[NV_NVDLA_CDMA_IMG_pack.scala 207:38:@8621.4]
  assign _GEN_14 = _T_312 ? _T_274 : _T_257; // @[NV_NVDLA_CDMA_IMG_pack.scala 186:19:@8581.4]
  assign _T_284 = ~ io_is_running; // @[NV_NVDLA_CDMA_IMG_pack.scala 197:26:@8595.4]
  assign _T_288 = io_sg2pack_img_pd_valid ? 1'h1 : _T_281; // @[NV_NVDLA_CDMA_IMG_pack.scala 199:25:@8596.4]
  assign _T_289 = _T_303 ? 1'h0 : _T_288; // @[NV_NVDLA_CDMA_IMG_pack.scala 198:25:@8597.4]
  assign _T_290 = _T_284 ? 1'h0 : _T_289; // @[NV_NVDLA_CDMA_IMG_pack.scala 197:25:@8598.4]
  assign _T_311 = _T_305 & _T_224; // @[NV_NVDLA_CDMA_IMG_pack.scala 206:108:@8620.4]
  assign _T_319 = _T_301 & _T_253; // @[NV_NVDLA_CDMA_IMG_pack.scala 212:52:@8632.4]
  assign _T_320 = _T_319 & _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 212:69:@8633.4]
  assign _T_322 = _T_301 & _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 213:52:@8635.4]
  assign _T_323 = _T_322 & _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 213:68:@8636.4]
  assign _T_329 = _T_320 & _T_120; // @[NV_NVDLA_CDMA_IMG_pack.scala 215:99:@8642.4]
  assign _T_334 = _T_323 & _T_120; // @[NV_NVDLA_CDMA_IMG_pack.scala 216:98:@8647.4]
  assign _T_382 = _T_358 + 7'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 254:47:@8675.4]
  assign _T_383 = _T_358 + 7'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 254:47:@8676.4]
  assign _T_384 = _T_361 + 7'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 255:47:@8677.4]
  assign _T_385 = _T_361 + 7'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 255:47:@8678.4]
  assign _T_387 = _T_123 ? 7'h0 : _T_383; // @[NV_NVDLA_CDMA_IMG_pack.scala 256:30:@8679.4]
  assign _T_389 = _T_123 ? 7'h0 : _T_385; // @[NV_NVDLA_CDMA_IMG_pack.scala 257:30:@8680.4]
  assign _T_392 = _T_358[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:65:@8682.4]
  assign _T_393 = _T_358[6:1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:87:@8683.4]
  assign _T_395 = {1'h0,_T_392,_T_393}; // @[Cat.scala 30:58:@8685.4]
  assign _T_397 = _T_361[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 259:43:@8686.4]
  assign _T_398 = _T_361[6:1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 259:65:@8687.4]
  assign _T_400 = {1'h1,_T_397,_T_398}; // @[Cat.scala 30:58:@8689.4]
  assign _T_401 = _T_253 ? _T_395 : _T_400; // @[NV_NVDLA_CDMA_IMG_pack.scala 258:18:@8690.4]
  assign _T_403 = _T_283 & _T_253; // @[NV_NVDLA_CDMA_IMG_pack.scala 279:45:@8708.4]
  assign _T_404 = _T_123 | _T_403; // @[NV_NVDLA_CDMA_IMG_pack.scala 279:35:@8709.4]
  assign _GEN_15 = _T_404 ? _T_387 : _T_358; // @[NV_NVDLA_CDMA_IMG_pack.scala 262:20:@8692.4]
  assign _T_405 = _T_283 & _T_246; // @[NV_NVDLA_CDMA_IMG_pack.scala 280:45:@8711.4]
  assign _T_406 = _T_123 | _T_405; // @[NV_NVDLA_CDMA_IMG_pack.scala 280:35:@8712.4]
  assign _GEN_16 = _T_406 ? _T_389 : _T_361; // @[NV_NVDLA_CDMA_IMG_pack.scala 265:20:@8695.4]
  assign _GEN_19 = _T_283 ? _T_370 : _T_373; // @[NV_NVDLA_CDMA_IMG_pack.scala 274:16:@8704.4]
  assign _GEN_85 = {{8'd0}, _T_160}; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8718.4]
  assign _T_413 = _T_409 + _GEN_85; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8718.4]
  assign _T_414 = _T_409 + _GEN_85; // @[NV_NVDLA_CDMA_IMG_pack.scala 289:50:@8719.4]
  assign _GEN_86 = {{8'd0}, _T_163}; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8720.4]
  assign _T_415 = _T_412 + _GEN_86; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8720.4]
  assign _T_416 = _T_412 + _GEN_86; // @[NV_NVDLA_CDMA_IMG_pack.scala 290:50:@8721.4]
  assign _T_417 = _T_414 > _T_132; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:57:@8722.4]
  assign _T_418 = _T_414 > _T_129; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:98:@8723.4]
  assign _T_419 = _T_414 > _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 291:139:@8724.4]
  assign _T_421 = {_T_417,_T_418,_T_419}; // @[Cat.scala 30:58:@8726.4]
  assign _T_422 = _T_416 > _T_132; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:57:@8727.4]
  assign _T_423 = _T_416 > _T_129; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:98:@8728.4]
  assign _T_424 = _T_416 > _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 292:139:@8729.4]
  assign _T_426 = {_T_422,_T_423,_T_424}; // @[Cat.scala 30:58:@8731.4]
  assign _T_431 = _T_123 | _T_329; // @[NV_NVDLA_CDMA_IMG_pack.scala 298:50:@8735.6]
  assign _T_433 = _T_431 ? 14'h0 : _T_414; // @[NV_NVDLA_CDMA_IMG_pack.scala 298:32:@8736.6]
  assign _GEN_20 = _T_404 ? _T_433 : _T_409; // @[NV_NVDLA_CDMA_IMG_pack.scala 297:22:@8734.4]
  assign _T_434 = _T_123 | _T_334; // @[NV_NVDLA_CDMA_IMG_pack.scala 301:50:@8740.6]
  assign _T_436 = _T_434 ? 14'h0 : _T_416; // @[NV_NVDLA_CDMA_IMG_pack.scala 301:32:@8741.6]
  assign _GEN_21 = _T_406 ? _T_436 : _T_412; // @[NV_NVDLA_CDMA_IMG_pack.scala 300:22:@8739.4]
  assign _T_453 = _T_414 - _GEN_85; // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8752.4]
  assign _T_454 = $unsigned(_T_453); // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8753.4]
  assign _T_455 = _T_454[13:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 316:50:@8754.4]
  assign _T_456 = _T_455 > _T_129; // @[NV_NVDLA_CDMA_IMG_pack.scala 317:57:@8755.4]
  assign _T_457 = _T_455 > _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 317:99:@8756.4]
  assign _T_458 = {_T_456,_T_457}; // @[Cat.scala 30:58:@8757.4]
  assign _T_459 = _T_421[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:60:@8758.4]
  assign _T_460 = ~ _T_459; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:35:@8759.4]
  assign _T_466 = _T_458[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:62:@8761.4]
  assign _T_467 = ~ _T_466; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:37:@8762.4]
  assign _T_473 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_142; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:93:@8764.4]
  assign _T_474 = ~ _T_473; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:67:@8765.4]
  assign _T_480 = _T_467 ? _T_474 : 287'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 319:36:@8767.4]
  assign _T_481 = _T_460 ? 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : _T_480; // @[NV_NVDLA_CDMA_IMG_pack.scala 318:34:@8768.4]
  assign _T_482 = _T_421[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:60:@8769.4]
  assign _T_483 = ~ _T_482; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:35:@8770.4]
  assign _T_489 = _T_458[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:62:@8772.4]
  assign _T_490 = ~ _T_489; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:37:@8773.4]
  assign _T_496 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_148; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:92:@8775.4]
  assign _T_502 = _T_490 ? _T_496 : 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff; // @[NV_NVDLA_CDMA_IMG_pack.scala 322:36:@8777.4]
  assign _T_503 = _T_483 ? 287'h0 : _T_502; // @[NV_NVDLA_CDMA_IMG_pack.scala 321:34:@8778.4]
  assign _T_504 = _T_421[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:59:@8779.4]
  assign _T_505 = ~ _T_504; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:34:@8780.4]
  assign _T_516 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_154; // @[NV_NVDLA_CDMA_IMG_pack.scala 325:58:@8783.4]
  assign _T_517 = _T_505 ? 287'h0 : _T_516; // @[NV_NVDLA_CDMA_IMG_pack.scala 324:33:@8784.4]
  assign _T_518 = _T_481 | _T_503; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:55:@8786.4]
  assign _T_438 = _T_517[31:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 306:37:@8744.4 NV_NVDLA_CDMA_IMG_pack.scala 324:27:@8785.4]
  assign _T_519 = ~ _T_438; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:84:@8787.4]
  assign _GEN_88 = {{255'd0}, _T_519}; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:82:@8788.4]
  assign _T_520 = _T_518 & _GEN_88; // @[NV_NVDLA_CDMA_IMG_pack.scala 326:82:@8788.4]
  assign _T_521 = _T_416 - _GEN_86; // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8790.4]
  assign _T_522 = $unsigned(_T_521); // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8791.4]
  assign _T_523 = _T_522[13:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 328:50:@8792.4]
  assign _T_524 = _T_523 > _T_129; // @[NV_NVDLA_CDMA_IMG_pack.scala 329:57:@8793.4]
  assign _T_525 = _T_523 > _T_126; // @[NV_NVDLA_CDMA_IMG_pack.scala 329:99:@8794.4]
  assign _T_526 = {_T_524,_T_525}; // @[Cat.scala 30:58:@8795.4]
  assign _T_527 = _T_426[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:60:@8796.4]
  assign _T_528 = ~ _T_527; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:35:@8797.4]
  assign _T_534 = _T_526[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:62:@8799.4]
  assign _T_535 = ~ _T_534; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:37:@8800.4]
  assign _T_541 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_145; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:93:@8802.4]
  assign _T_542 = ~ _T_541; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:67:@8803.4]
  assign _T_548 = _T_535 ? _T_542 : 287'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 331:36:@8805.4]
  assign _T_549 = _T_528 ? 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : _T_548; // @[NV_NVDLA_CDMA_IMG_pack.scala 330:34:@8806.4]
  assign _T_550 = _T_426[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:60:@8807.4]
  assign _T_551 = ~ _T_550; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:35:@8808.4]
  assign _T_557 = _T_526[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:62:@8810.4]
  assign _T_558 = ~ _T_557; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:37:@8811.4]
  assign _T_564 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_151; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:92:@8813.4]
  assign _T_570 = _T_558 ? _T_564 : 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff; // @[NV_NVDLA_CDMA_IMG_pack.scala 334:36:@8815.4]
  assign _T_571 = _T_551 ? 287'h0 : _T_570; // @[NV_NVDLA_CDMA_IMG_pack.scala 333:34:@8816.4]
  assign _T_572 = _T_426[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:59:@8817.4]
  assign _T_573 = ~ _T_572; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:34:@8818.4]
  assign _T_584 = 287'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff << _T_157; // @[NV_NVDLA_CDMA_IMG_pack.scala 337:58:@8821.4]
  assign _T_585 = _T_573 ? 287'h0 : _T_584; // @[NV_NVDLA_CDMA_IMG_pack.scala 336:33:@8822.4]
  assign _T_586 = _T_549 | _T_571; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:55:@8824.4]
  assign _T_442 = _T_585[31:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 308:37:@8746.4 NV_NVDLA_CDMA_IMG_pack.scala 336:27:@8823.4]
  assign _T_587 = ~ _T_442; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:84:@8825.4]
  assign _GEN_90 = {{255'd0}, _T_587}; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:82:@8826.4]
  assign _T_588 = _T_586 & _GEN_90; // @[NV_NVDLA_CDMA_IMG_pack.scala 338:82:@8826.4]
  assign _T_440 = _T_520[31:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 307:36:@8745.4 NV_NVDLA_CDMA_IMG_pack.scala 326:26:@8789.4]
  assign _T_444 = _T_588[31:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 309:36:@8747.4 NV_NVDLA_CDMA_IMG_pack.scala 338:26:@8827.4]
  assign _T_590 = _T_253 ? _T_440 : _T_444; // @[NV_NVDLA_CDMA_IMG_pack.scala 340:22:@8829.4]
  assign _T_623 = _T_268 & _T_250; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:41:@8861.6]
  assign _T_624 = _T_623 & _T_240; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:58:@8862.6]
  assign _T_625 = _T_624 & _T_120; // @[NV_NVDLA_CDMA_IMG_pack.scala 364:73:@8863.6]
  assign _T_626 = _T_121 & _T_311; // @[NV_NVDLA_CDMA_IMG_pack.scala 366:37:@8866.6]
  assign _GEN_24 = _T_283 ? _T_246 : _T_604; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_25 = _T_283 ? 3'h0 : _T_607; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_26 = _T_283 ? _T_303 : _T_610; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_27 = _T_283 ? _T_303 : _T_613; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_28 = _T_283 ? _T_625 : _T_616; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_29 = _T_283 ? _T_223 : _T_619; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_30 = _T_283 ? _T_626 : _T_622; // @[NV_NVDLA_CDMA_IMG_pack.scala 359:13:@8856.4]
  assign _GEN_32 = _T_337 ? _T_604 : _T_639; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_33 = _T_337 ? _T_607 : _T_647; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_34 = _T_337 ? _T_610 : _T_655; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_35 = _T_337 ? _T_613 : _T_663; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_36 = _T_337 ? _T_616 : _T_671; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_37 = _T_337 ? _T_619 : _T_679; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_38 = _T_337 ? _T_622 : _T_687; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8912.4]
  assign _GEN_42 = _T_631 ? _T_639 : _T_642; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_43 = _T_631 ? _T_647 : _T_650; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_44 = _T_631 ? _T_655 : _T_658; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_45 = _T_631 ? _T_663 : _T_666; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_46 = _T_631 ? _T_671 : _T_674; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_47 = _T_631 ? _T_679 : _T_682; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _GEN_48 = _T_631 ? _T_687 : _T_690; // @[NV_NVDLA_CDMA_IMG_pack.scala 413:25:@8925.4]
  assign _T_703 = io_pixel_early_end & _T_674; // @[NV_NVDLA_CDMA_IMG_pack.scala 437:43:@8937.4]
  assign _T_704 = _T_634 & io_pixel_planar; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:34:@8938.4]
  assign _T_705 = ~ _T_703; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:54:@8939.4]
  assign _T_706 = _T_704 & _T_705; // @[NV_NVDLA_CDMA_IMG_pack.scala 438:52:@8940.4]
  assign _GEN_51 = _T_706 ? _T_650 : _T_712; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _GEN_52 = _T_706 ? _T_658 : _T_715; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _GEN_53 = _T_706 ? _T_666 : _T_718; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _GEN_54 = _T_706 ? _T_674 : _T_721; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _GEN_55 = _T_706 ? _T_682 : _T_724; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _GEN_56 = _T_706 ? _T_690 : _T_727; // @[NV_NVDLA_CDMA_IMG_pack.scala 449:22:@8949.4]
  assign _T_732 = _T_634 & _T_703; // @[NV_NVDLA_CDMA_IMG_pack.scala 468:55:@8959.4]
  assign _T_733 = _T_249 | _T_732; // @[NV_NVDLA_CDMA_IMG_pack.scala 468:41:@8960.4]
  assign _T_734 = _T_733 ? _T_634 : _T_709; // @[NV_NVDLA_CDMA_IMG_pack.scala 470:25:@8961.4]
  assign _T_735 = _T_733 ? _T_650 : _T_712; // @[NV_NVDLA_CDMA_IMG_pack.scala 471:27:@8962.4]
  assign _T_736 = _T_733 ? _T_658 : _T_715; // @[NV_NVDLA_CDMA_IMG_pack.scala 472:31:@8963.4]
  assign _T_737 = _T_733 ? _T_666 : _T_718; // @[NV_NVDLA_CDMA_IMG_pack.scala 473:30:@8964.4]
  assign _T_738 = _T_733 ? _T_674 : _T_721; // @[NV_NVDLA_CDMA_IMG_pack.scala 474:34:@8965.4]
  assign _T_739 = _T_733 ? _T_682 : _T_724; // @[NV_NVDLA_CDMA_IMG_pack.scala 475:32:@8966.4]
  assign _T_740 = _T_733 ? _T_690 : _T_727; // @[NV_NVDLA_CDMA_IMG_pack.scala 476:31:@8967.4]
  assign _T_741 = ~ _T_642; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:46:@8968.4]
  assign _T_742 = _T_123 | _T_741; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:44:@8969.4]
  assign _T_745 = _T_730 + 2'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:94:@8970.4]
  assign _T_746 = _T_730 + 2'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:94:@8971.4]
  assign _T_747 = _T_742 ? 2'h0 : _T_746; // @[NV_NVDLA_CDMA_IMG_pack.scala 479:26:@8972.4]
  assign _GEN_57 = _T_634 ? _T_747 : _T_730; // @[NV_NVDLA_CDMA_IMG_pack.scala 481:17:@8973.4]
  assign _GEN_58 = _T_734 ? _T_735 : _T_761; // @[NV_NVDLA_CDMA_IMG_pack.scala 495:20:@8984.4]
  assign _GEN_59 = _T_123 ? 4'h1 : _T_764; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  assign _GEN_60 = _T_123 ? io_sg2pack_mn_enable : _T_767; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  assign _GEN_61 = _T_123 ? io_pixel_uint : _T_770; // @[NV_NVDLA_CDMA_IMG_pack.scala 498:23:@8987.4]
  assign _T_775 = {2'h0,_T_764}; // @[Cat.scala 30:58:@8993.4]
  assign _T_778 = {_T_761,_T_770,_T_767,1'h0}; // @[Cat.scala 30:58:@8996.4]
  assign _T_813 = _T_702[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9014.4]
  assign _T_814 = io_pixel_packed_10b | _T_813; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9015.4]
  assign _T_815 = _T_696[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9016.4]
  assign _T_816 = _T_814 | _T_815; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9017.4]
  assign _T_818 = io_img2sbuf_p0_rd_data[7:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9018.4]
  assign _T_819 = _T_816 ? 8'h0 : _T_818; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9019.4]
  assign _T_820 = _T_702[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9020.4]
  assign _T_821 = io_pixel_packed_10b | _T_820; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9021.4]
  assign _T_822 = _T_696[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9022.4]
  assign _T_823 = _T_821 | _T_822; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9023.4]
  assign _T_825 = io_img2sbuf_p0_rd_data[15:8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9024.4]
  assign _T_826 = _T_823 ? 8'h0 : _T_825; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9025.4]
  assign _T_827 = _T_702[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9026.4]
  assign _T_828 = io_pixel_packed_10b | _T_827; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9027.4]
  assign _T_829 = _T_696[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9028.4]
  assign _T_830 = _T_828 | _T_829; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9029.4]
  assign _T_832 = io_img2sbuf_p0_rd_data[23:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9030.4]
  assign _T_833 = _T_830 ? 8'h0 : _T_832; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9031.4]
  assign _T_834 = _T_702[3]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9032.4]
  assign _T_835 = io_pixel_packed_10b | _T_834; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9033.4]
  assign _T_836 = _T_696[3]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9034.4]
  assign _T_837 = _T_835 | _T_836; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9035.4]
  assign _T_839 = io_img2sbuf_p0_rd_data[31:24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9036.4]
  assign _T_840 = _T_837 ? 8'h0 : _T_839; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9037.4]
  assign _T_841 = _T_702[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9038.4]
  assign _T_842 = io_pixel_packed_10b | _T_841; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9039.4]
  assign _T_843 = _T_696[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9040.4]
  assign _T_844 = _T_842 | _T_843; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9041.4]
  assign _T_846 = io_img2sbuf_p0_rd_data[39:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9042.4]
  assign _T_847 = _T_844 ? 8'h0 : _T_846; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9043.4]
  assign _T_848 = _T_702[5]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9044.4]
  assign _T_849 = io_pixel_packed_10b | _T_848; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9045.4]
  assign _T_850 = _T_696[5]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9046.4]
  assign _T_851 = _T_849 | _T_850; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9047.4]
  assign _T_853 = io_img2sbuf_p0_rd_data[47:40]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9048.4]
  assign _T_854 = _T_851 ? 8'h0 : _T_853; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9049.4]
  assign _T_855 = _T_702[6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9050.4]
  assign _T_856 = io_pixel_packed_10b | _T_855; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9051.4]
  assign _T_857 = _T_696[6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9052.4]
  assign _T_858 = _T_856 | _T_857; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9053.4]
  assign _T_860 = io_img2sbuf_p0_rd_data[55:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9054.4]
  assign _T_861 = _T_858 ? 8'h0 : _T_860; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9055.4]
  assign _T_862 = _T_702[7]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9056.4]
  assign _T_863 = io_pixel_packed_10b | _T_862; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9057.4]
  assign _T_864 = _T_696[7]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9058.4]
  assign _T_865 = _T_863 | _T_864; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9059.4]
  assign _T_867 = io_img2sbuf_p0_rd_data[63:56]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9060.4]
  assign _T_868 = _T_865 ? 8'h0 : _T_867; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9061.4]
  assign _T_869 = _T_702[8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9062.4]
  assign _T_870 = io_pixel_packed_10b | _T_869; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9063.4]
  assign _T_871 = _T_696[8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9064.4]
  assign _T_872 = _T_870 | _T_871; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9065.4]
  assign _T_874 = io_img2sbuf_p0_rd_data[71:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9066.4]
  assign _T_875 = _T_872 ? 8'h0 : _T_874; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9067.4]
  assign _T_876 = _T_702[9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9068.4]
  assign _T_877 = io_pixel_packed_10b | _T_876; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9069.4]
  assign _T_878 = _T_696[9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9070.4]
  assign _T_879 = _T_877 | _T_878; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9071.4]
  assign _T_881 = io_img2sbuf_p0_rd_data[79:72]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9072.4]
  assign _T_882 = _T_879 ? 8'h0 : _T_881; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9073.4]
  assign _T_883 = _T_702[10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9074.4]
  assign _T_884 = io_pixel_packed_10b | _T_883; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9075.4]
  assign _T_885 = _T_696[10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9076.4]
  assign _T_886 = _T_884 | _T_885; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9077.4]
  assign _T_888 = io_img2sbuf_p0_rd_data[87:80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9078.4]
  assign _T_889 = _T_886 ? 8'h0 : _T_888; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9079.4]
  assign _T_890 = _T_702[11]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9080.4]
  assign _T_891 = io_pixel_packed_10b | _T_890; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9081.4]
  assign _T_892 = _T_696[11]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9082.4]
  assign _T_893 = _T_891 | _T_892; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9083.4]
  assign _T_895 = io_img2sbuf_p0_rd_data[95:88]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9084.4]
  assign _T_896 = _T_893 ? 8'h0 : _T_895; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9085.4]
  assign _T_897 = _T_702[12]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9086.4]
  assign _T_898 = io_pixel_packed_10b | _T_897; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9087.4]
  assign _T_899 = _T_696[12]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9088.4]
  assign _T_900 = _T_898 | _T_899; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9089.4]
  assign _T_902 = io_img2sbuf_p0_rd_data[103:96]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9090.4]
  assign _T_903 = _T_900 ? 8'h0 : _T_902; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9091.4]
  assign _T_904 = _T_702[13]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9092.4]
  assign _T_905 = io_pixel_packed_10b | _T_904; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9093.4]
  assign _T_906 = _T_696[13]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9094.4]
  assign _T_907 = _T_905 | _T_906; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9095.4]
  assign _T_909 = io_img2sbuf_p0_rd_data[111:104]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9096.4]
  assign _T_910 = _T_907 ? 8'h0 : _T_909; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9097.4]
  assign _T_911 = _T_702[14]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9098.4]
  assign _T_912 = io_pixel_packed_10b | _T_911; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9099.4]
  assign _T_913 = _T_696[14]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9100.4]
  assign _T_914 = _T_912 | _T_913; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9101.4]
  assign _T_916 = io_img2sbuf_p0_rd_data[119:112]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9102.4]
  assign _T_917 = _T_914 ? 8'h0 : _T_916; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9103.4]
  assign _T_918 = _T_702[15]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9104.4]
  assign _T_919 = io_pixel_packed_10b | _T_918; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9105.4]
  assign _T_920 = _T_696[15]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9106.4]
  assign _T_921 = _T_919 | _T_920; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9107.4]
  assign _T_923 = io_img2sbuf_p0_rd_data[127:120]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9108.4]
  assign _T_924 = _T_921 ? 8'h0 : _T_923; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9109.4]
  assign _T_925 = _T_702[16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9110.4]
  assign _T_926 = io_pixel_packed_10b | _T_925; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9111.4]
  assign _T_927 = _T_696[16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9112.4]
  assign _T_928 = _T_926 | _T_927; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9113.4]
  assign _T_930 = io_img2sbuf_p0_rd_data[135:128]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9114.4]
  assign _T_931 = _T_928 ? 8'h0 : _T_930; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9115.4]
  assign _T_932 = _T_702[17]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9116.4]
  assign _T_933 = io_pixel_packed_10b | _T_932; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9117.4]
  assign _T_934 = _T_696[17]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9118.4]
  assign _T_935 = _T_933 | _T_934; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9119.4]
  assign _T_937 = io_img2sbuf_p0_rd_data[143:136]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9120.4]
  assign _T_938 = _T_935 ? 8'h0 : _T_937; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9121.4]
  assign _T_939 = _T_702[18]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9122.4]
  assign _T_940 = io_pixel_packed_10b | _T_939; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9123.4]
  assign _T_941 = _T_696[18]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9124.4]
  assign _T_942 = _T_940 | _T_941; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9125.4]
  assign _T_944 = io_img2sbuf_p0_rd_data[151:144]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9126.4]
  assign _T_945 = _T_942 ? 8'h0 : _T_944; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9127.4]
  assign _T_946 = _T_702[19]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9128.4]
  assign _T_947 = io_pixel_packed_10b | _T_946; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9129.4]
  assign _T_948 = _T_696[19]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9130.4]
  assign _T_949 = _T_947 | _T_948; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9131.4]
  assign _T_951 = io_img2sbuf_p0_rd_data[159:152]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9132.4]
  assign _T_952 = _T_949 ? 8'h0 : _T_951; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9133.4]
  assign _T_953 = _T_702[20]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9134.4]
  assign _T_954 = io_pixel_packed_10b | _T_953; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9135.4]
  assign _T_955 = _T_696[20]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9136.4]
  assign _T_956 = _T_954 | _T_955; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9137.4]
  assign _T_958 = io_img2sbuf_p0_rd_data[167:160]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9138.4]
  assign _T_959 = _T_956 ? 8'h0 : _T_958; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9139.4]
  assign _T_960 = _T_702[21]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9140.4]
  assign _T_961 = io_pixel_packed_10b | _T_960; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9141.4]
  assign _T_962 = _T_696[21]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9142.4]
  assign _T_963 = _T_961 | _T_962; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9143.4]
  assign _T_965 = io_img2sbuf_p0_rd_data[175:168]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9144.4]
  assign _T_966 = _T_963 ? 8'h0 : _T_965; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9145.4]
  assign _T_967 = _T_702[22]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9146.4]
  assign _T_968 = io_pixel_packed_10b | _T_967; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9147.4]
  assign _T_969 = _T_696[22]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9148.4]
  assign _T_970 = _T_968 | _T_969; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9149.4]
  assign _T_972 = io_img2sbuf_p0_rd_data[183:176]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9150.4]
  assign _T_973 = _T_970 ? 8'h0 : _T_972; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9151.4]
  assign _T_974 = _T_702[23]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9152.4]
  assign _T_975 = io_pixel_packed_10b | _T_974; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9153.4]
  assign _T_976 = _T_696[23]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9154.4]
  assign _T_977 = _T_975 | _T_976; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9155.4]
  assign _T_979 = io_img2sbuf_p0_rd_data[191:184]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9156.4]
  assign _T_980 = _T_977 ? 8'h0 : _T_979; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9157.4]
  assign _T_981 = _T_702[24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9158.4]
  assign _T_982 = io_pixel_packed_10b | _T_981; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9159.4]
  assign _T_983 = _T_696[24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9160.4]
  assign _T_984 = _T_982 | _T_983; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9161.4]
  assign _T_986 = io_img2sbuf_p0_rd_data[199:192]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9162.4]
  assign _T_987 = _T_984 ? 8'h0 : _T_986; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9163.4]
  assign _T_988 = _T_702[25]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9164.4]
  assign _T_989 = io_pixel_packed_10b | _T_988; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9165.4]
  assign _T_990 = _T_696[25]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9166.4]
  assign _T_991 = _T_989 | _T_990; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9167.4]
  assign _T_993 = io_img2sbuf_p0_rd_data[207:200]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9168.4]
  assign _T_994 = _T_991 ? 8'h0 : _T_993; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9169.4]
  assign _T_995 = _T_702[26]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9170.4]
  assign _T_996 = io_pixel_packed_10b | _T_995; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9171.4]
  assign _T_997 = _T_696[26]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9172.4]
  assign _T_998 = _T_996 | _T_997; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9173.4]
  assign _T_1000 = io_img2sbuf_p0_rd_data[215:208]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9174.4]
  assign _T_1001 = _T_998 ? 8'h0 : _T_1000; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9175.4]
  assign _T_1002 = _T_702[27]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9176.4]
  assign _T_1003 = io_pixel_packed_10b | _T_1002; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9177.4]
  assign _T_1004 = _T_696[27]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9178.4]
  assign _T_1005 = _T_1003 | _T_1004; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9179.4]
  assign _T_1007 = io_img2sbuf_p0_rd_data[223:216]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9180.4]
  assign _T_1008 = _T_1005 ? 8'h0 : _T_1007; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9181.4]
  assign _T_1009 = _T_702[28]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9182.4]
  assign _T_1010 = io_pixel_packed_10b | _T_1009; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9183.4]
  assign _T_1011 = _T_696[28]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9184.4]
  assign _T_1012 = _T_1010 | _T_1011; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9185.4]
  assign _T_1014 = io_img2sbuf_p0_rd_data[231:224]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9186.4]
  assign _T_1015 = _T_1012 ? 8'h0 : _T_1014; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9187.4]
  assign _T_1016 = _T_702[29]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9188.4]
  assign _T_1017 = io_pixel_packed_10b | _T_1016; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9189.4]
  assign _T_1018 = _T_696[29]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9190.4]
  assign _T_1019 = _T_1017 | _T_1018; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9191.4]
  assign _T_1021 = io_img2sbuf_p0_rd_data[239:232]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9192.4]
  assign _T_1022 = _T_1019 ? 8'h0 : _T_1021; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9193.4]
  assign _T_1023 = _T_702[30]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9194.4]
  assign _T_1024 = io_pixel_packed_10b | _T_1023; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9195.4]
  assign _T_1025 = _T_696[30]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9196.4]
  assign _T_1026 = _T_1024 | _T_1025; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9197.4]
  assign _T_1028 = io_img2sbuf_p0_rd_data[247:240]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9198.4]
  assign _T_1029 = _T_1026 ? 8'h0 : _T_1028; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9199.4]
  assign _T_1030 = _T_702[31]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:43:@9200.4]
  assign _T_1031 = io_pixel_packed_10b | _T_1030; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:33:@9201.4]
  assign _T_1032 = _T_696[31]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:55:@9202.4]
  assign _T_1033 = _T_1031 | _T_1032; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:46:@9203.4]
  assign _T_1035 = io_img2sbuf_p0_rd_data[255:248]; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:82:@9204.4]
  assign _T_1036 = _T_1033 ? 8'h0 : _T_1035; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:13:@9205.4]
  assign _T_1081 = {_T_868,_T_861,_T_854,_T_847,_T_840,_T_833,_T_826,_T_819}; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9245.4]
  assign _T_1089 = {_T_924,_T_917,_T_910,_T_903,_T_896,_T_889,_T_882,_T_875,_T_1081}; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9253.4]
  assign _T_1096 = {_T_980,_T_973,_T_966,_T_959,_T_952,_T_945,_T_938,_T_931}; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9260.4]
  assign _T_1105 = {_T_1036,_T_1029,_T_1022,_T_1015,_T_1008,_T_1001,_T_994,_T_987,_T_1096,_T_1089}; // @[NV_NVDLA_CDMA_IMG_pack.scala 531:139:@9269.4]
  assign _T_1522 = _T_704 & _T_642; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:54:@9657.4]
  assign _T_1524 = _T_730 == 2'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:87:@9658.4]
  assign _T_1525 = _T_1522 & _T_1524; // @[NV_NVDLA_CDMA_IMG_pack.scala 559:70:@9659.4]
  assign _T_1106 = _T_1525 ? _T_1105 : _T_785; // @[NV_NVDLA_CDMA_IMG_pack.scala 533:20:@9270.4]
  assign _T_1529 = _T_730 == 2'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 560:87:@9663.4]
  assign _T_1530 = _T_1522 & _T_1529; // @[NV_NVDLA_CDMA_IMG_pack.scala 560:70:@9664.4]
  assign _T_1107 = _T_1530 ? _T_1105 : _T_788; // @[NV_NVDLA_CDMA_IMG_pack.scala 534:20:@9271.4]
  assign _T_1108 = {_T_1107,_T_1106}; // @[Cat.scala 30:58:@9272.4]
  assign _T_1109 = _T_1108[15:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9273.4]
  assign _T_1110 = _T_782[7:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9274.4]
  assign _T_1112 = _T_1108[31:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9276.4]
  assign _T_1113 = _T_782[15:8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9277.4]
  assign _T_1115 = _T_1108[47:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9279.4]
  assign _T_1116 = _T_782[23:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9280.4]
  assign _T_1118 = _T_1108[63:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9282.4]
  assign _T_1119 = _T_782[31:24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9283.4]
  assign _T_1121 = _T_1108[79:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9285.4]
  assign _T_1122 = _T_782[39:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9286.4]
  assign _T_1124 = _T_1108[95:80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9288.4]
  assign _T_1125 = _T_782[47:40]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9289.4]
  assign _T_1127 = _T_1108[111:96]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9291.4]
  assign _T_1128 = _T_782[55:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9292.4]
  assign _T_1130 = _T_1108[127:112]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9294.4]
  assign _T_1131 = _T_782[63:56]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9295.4]
  assign _T_1133 = _T_1108[143:128]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9297.4]
  assign _T_1134 = _T_782[71:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9298.4]
  assign _T_1136 = _T_1108[159:144]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9300.4]
  assign _T_1137 = _T_782[79:72]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9301.4]
  assign _T_1139 = _T_1108[175:160]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9303.4]
  assign _T_1140 = _T_782[87:80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9304.4]
  assign _T_1142 = _T_1108[191:176]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9306.4]
  assign _T_1143 = _T_782[95:88]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9307.4]
  assign _T_1145 = _T_1108[207:192]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9309.4]
  assign _T_1146 = _T_782[103:96]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9310.4]
  assign _T_1148 = _T_1108[223:208]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9312.4]
  assign _T_1149 = _T_782[111:104]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9313.4]
  assign _T_1151 = _T_1108[239:224]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9315.4]
  assign _T_1152 = _T_782[119:112]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9316.4]
  assign _T_1154 = _T_1108[255:240]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9318.4]
  assign _T_1155 = _T_782[127:120]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9319.4]
  assign _T_1157 = _T_1108[271:256]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9321.4]
  assign _T_1158 = _T_782[135:128]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9322.4]
  assign _T_1160 = _T_1108[287:272]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9324.4]
  assign _T_1161 = _T_782[143:136]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9325.4]
  assign _T_1163 = _T_1108[303:288]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9327.4]
  assign _T_1164 = _T_782[151:144]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9328.4]
  assign _T_1166 = _T_1108[319:304]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9330.4]
  assign _T_1167 = _T_782[159:152]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9331.4]
  assign _T_1169 = _T_1108[335:320]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9333.4]
  assign _T_1170 = _T_782[167:160]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9334.4]
  assign _T_1172 = _T_1108[351:336]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9336.4]
  assign _T_1173 = _T_782[175:168]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9337.4]
  assign _T_1175 = _T_1108[367:352]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9339.4]
  assign _T_1176 = _T_782[183:176]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9340.4]
  assign _T_1178 = _T_1108[383:368]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9342.4]
  assign _T_1179 = _T_782[191:184]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9343.4]
  assign _T_1181 = _T_1108[399:384]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9345.4]
  assign _T_1182 = _T_782[199:192]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9346.4]
  assign _T_1184 = _T_1108[415:400]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9348.4]
  assign _T_1185 = _T_782[207:200]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9349.4]
  assign _T_1187 = _T_1108[431:416]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9351.4]
  assign _T_1188 = _T_782[215:208]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9352.4]
  assign _T_1190 = _T_1108[447:432]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9354.4]
  assign _T_1191 = _T_782[223:216]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9355.4]
  assign _T_1193 = _T_1108[463:448]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9357.4]
  assign _T_1194 = _T_782[231:224]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9358.4]
  assign _T_1196 = _T_1108[479:464]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9360.4]
  assign _T_1197 = _T_782[239:232]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9361.4]
  assign _T_1199 = _T_1108[495:480]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9363.4]
  assign _T_1200 = _T_782[247:240]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9364.4]
  assign _T_1202 = _T_1108[511:496]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:17:@9366.4]
  assign _T_1203 = _T_782[255:248]; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:45:@9367.4]
  assign _T_1245 = {_T_1118,_T_1119,_T_1115,_T_1116,_T_1112,_T_1113,_T_1109,_T_1110}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9404.4]
  assign _T_1249 = {_T_1130,_T_1131,_T_1127,_T_1128,_T_1124,_T_1125,_T_1121,_T_1122,_T_1245}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9408.4]
  assign _T_1252 = {_T_1142,_T_1143,_T_1139,_T_1140,_T_1136,_T_1137,_T_1133,_T_1134}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9411.4]
  assign _T_1257 = {_T_1154,_T_1155,_T_1151,_T_1152,_T_1148,_T_1149,_T_1145,_T_1146,_T_1252,_T_1249}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9416.4]
  assign _T_1260 = {_T_1166,_T_1167,_T_1163,_T_1164,_T_1160,_T_1161,_T_1157,_T_1158}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9419.4]
  assign _T_1264 = {_T_1178,_T_1179,_T_1175,_T_1176,_T_1172,_T_1173,_T_1169,_T_1170,_T_1260}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9423.4]
  assign _T_1267 = {_T_1190,_T_1191,_T_1187,_T_1188,_T_1184,_T_1185,_T_1181,_T_1182}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9426.4]
  assign _T_1272 = {_T_1202,_T_1203,_T_1199,_T_1200,_T_1196,_T_1197,_T_1193,_T_1194,_T_1267,_T_1264}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9431.4]
  assign _T_1273 = {_T_1272,_T_1257}; // @[NV_NVDLA_CDMA_IMG_pack.scala 537:63:@9432.4]
  assign _T_1275 = _T_730 == 2'h2; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:59:@9433.4]
  assign _T_1276 = io_pixel_planar & _T_1275; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:42:@9434.4]
  assign _T_1279 = io_pixel_planar & _T_1529; // @[NV_NVDLA_CDMA_IMG_pack.scala 539:85:@9436.4]
  assign _T_1282 = io_pixel_planar & _T_1524; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:41:@9438.4]
  assign _T_1284 = ~ io_pixel_packed_10b; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:87:@9440.4]
  assign _T_1285 = _T_249 & _T_1284; // @[NV_NVDLA_CDMA_IMG_pack.scala 540:85:@9441.4]
  assign _T_1289 = {_T_1276,_T_1279,_T_1282,_T_1285,io_pixel_packed_10b}; // @[Cat.scala 30:58:@9445.4]
  assign _T_1290 = _T_1289[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:68:@9446.4]
  assign _T_1294 = _T_1290 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@9448.4]
  assign _T_1295 = _T_1294 & _T_1105; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:73:@9449.4]
  assign _T_1296 = _T_1289[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:68:@9450.4]
  assign _T_1300 = _T_1296 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@9452.4]
  assign _T_1301 = _T_1273[255:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:82:@9453.4]
  assign _T_1302 = _T_1300 & _T_1301; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:73:@9454.4]
  assign _T_1303 = _T_1295 | _T_1302; // @[NV_NVDLA_CDMA_IMG_pack.scala 541:93:@9455.4]
  assign _T_1304 = _T_1289[3]; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:68:@9456.4]
  assign _T_1308 = _T_1304 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@9458.4]
  assign _T_1309 = _T_1273[511:256]; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:82:@9459.4]
  assign _T_1310 = _T_1308 & _T_1309; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:73:@9460.4]
  assign _T_1311 = _T_1303 | _T_1310; // @[NV_NVDLA_CDMA_IMG_pack.scala 542:115:@9461.4]
  assign _T_1312 = _T_1289[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:68:@9462.4]
  assign _T_1316 = _T_1312 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@9464.4]
  assign _T_1317 = _T_1273[767:512]; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:82:@9465.4]
  assign _T_1318 = _T_1316 & _T_1317; // @[NV_NVDLA_CDMA_IMG_pack.scala 544:73:@9466.4]
  assign _T_1319 = _T_1311 | _T_1318; // @[NV_NVDLA_CDMA_IMG_pack.scala 543:139:@9467.4]
  assign _T_1320 = _T_1525 ? _T_696 : _T_794; // @[NV_NVDLA_CDMA_IMG_pack.scala 548:25:@9468.4]
  assign _T_1321 = _T_1530 ? _T_696 : _T_797; // @[NV_NVDLA_CDMA_IMG_pack.scala 549:25:@9469.4]
  assign _T_1322 = {_T_1321,_T_1320}; // @[Cat.scala 30:58:@9470.4]
  assign _T_1323 = _T_1322[1:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9471.4]
  assign _T_1324 = _T_791[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9472.4]
  assign _T_1326 = _T_1322[3:2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9474.4]
  assign _T_1327 = _T_791[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9475.4]
  assign _T_1329 = _T_1322[5:4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9477.4]
  assign _T_1330 = _T_791[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9478.4]
  assign _T_1332 = _T_1322[7:6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9480.4]
  assign _T_1333 = _T_791[3]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9481.4]
  assign _T_1335 = _T_1322[9:8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9483.4]
  assign _T_1336 = _T_791[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9484.4]
  assign _T_1338 = _T_1322[11:10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9486.4]
  assign _T_1339 = _T_791[5]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9487.4]
  assign _T_1341 = _T_1322[13:12]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9489.4]
  assign _T_1342 = _T_791[6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9490.4]
  assign _T_1344 = _T_1322[15:14]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9492.4]
  assign _T_1345 = _T_791[7]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9493.4]
  assign _T_1347 = _T_1322[17:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9495.4]
  assign _T_1348 = _T_791[8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9496.4]
  assign _T_1350 = _T_1322[19:18]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9498.4]
  assign _T_1351 = _T_791[9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9499.4]
  assign _T_1353 = _T_1322[21:20]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9501.4]
  assign _T_1354 = _T_791[10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9502.4]
  assign _T_1356 = _T_1322[23:22]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9504.4]
  assign _T_1357 = _T_791[11]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9505.4]
  assign _T_1359 = _T_1322[25:24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9507.4]
  assign _T_1360 = _T_791[12]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9508.4]
  assign _T_1362 = _T_1322[27:26]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9510.4]
  assign _T_1363 = _T_791[13]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9511.4]
  assign _T_1365 = _T_1322[29:28]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9513.4]
  assign _T_1366 = _T_791[14]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9514.4]
  assign _T_1368 = _T_1322[31:30]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9516.4]
  assign _T_1369 = _T_791[15]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9517.4]
  assign _T_1371 = _T_1322[33:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9519.4]
  assign _T_1372 = _T_791[16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9520.4]
  assign _T_1374 = _T_1322[35:34]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9522.4]
  assign _T_1375 = _T_791[17]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9523.4]
  assign _T_1377 = _T_1322[37:36]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9525.4]
  assign _T_1378 = _T_791[18]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9526.4]
  assign _T_1380 = _T_1322[39:38]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9528.4]
  assign _T_1381 = _T_791[19]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9529.4]
  assign _T_1383 = _T_1322[41:40]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9531.4]
  assign _T_1384 = _T_791[20]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9532.4]
  assign _T_1386 = _T_1322[43:42]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9534.4]
  assign _T_1387 = _T_791[21]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9535.4]
  assign _T_1389 = _T_1322[45:44]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9537.4]
  assign _T_1390 = _T_791[22]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9538.4]
  assign _T_1392 = _T_1322[47:46]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9540.4]
  assign _T_1393 = _T_791[23]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9541.4]
  assign _T_1395 = _T_1322[49:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9543.4]
  assign _T_1396 = _T_791[24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9544.4]
  assign _T_1398 = _T_1322[51:50]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9546.4]
  assign _T_1399 = _T_791[25]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9547.4]
  assign _T_1401 = _T_1322[53:52]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9549.4]
  assign _T_1402 = _T_791[26]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9550.4]
  assign _T_1404 = _T_1322[55:54]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9552.4]
  assign _T_1405 = _T_791[27]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9553.4]
  assign _T_1407 = _T_1322[57:56]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9555.4]
  assign _T_1408 = _T_791[28]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9556.4]
  assign _T_1410 = _T_1322[59:58]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9558.4]
  assign _T_1411 = _T_791[29]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9559.4]
  assign _T_1413 = _T_1322[61:60]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9561.4]
  assign _T_1414 = _T_791[30]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9562.4]
  assign _T_1416 = _T_1322[63:62]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:22:@9564.4]
  assign _T_1417 = _T_791[31]; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:49:@9565.4]
  assign _T_1459 = {_T_1332,_T_1333,_T_1329,_T_1330,_T_1326,_T_1327,_T_1323,_T_1324}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9602.4]
  assign _T_1463 = {_T_1344,_T_1345,_T_1341,_T_1342,_T_1338,_T_1339,_T_1335,_T_1336,_T_1459}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9606.4]
  assign _T_1466 = {_T_1356,_T_1357,_T_1353,_T_1354,_T_1350,_T_1351,_T_1347,_T_1348}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9609.4]
  assign _T_1471 = {_T_1368,_T_1369,_T_1365,_T_1366,_T_1362,_T_1363,_T_1359,_T_1360,_T_1466,_T_1463}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9614.4]
  assign _T_1474 = {_T_1380,_T_1381,_T_1377,_T_1378,_T_1374,_T_1375,_T_1371,_T_1372}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9617.4]
  assign _T_1478 = {_T_1392,_T_1393,_T_1389,_T_1390,_T_1386,_T_1387,_T_1383,_T_1384,_T_1474}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9621.4]
  assign _T_1481 = {_T_1404,_T_1405,_T_1401,_T_1402,_T_1398,_T_1399,_T_1395,_T_1396}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9624.4]
  assign _T_1486 = {_T_1416,_T_1417,_T_1413,_T_1414,_T_1410,_T_1411,_T_1407,_T_1408,_T_1481,_T_1478}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9629.4]
  assign _T_1487 = {_T_1486,_T_1471}; // @[NV_NVDLA_CDMA_IMG_pack.scala 552:63:@9630.4]
  assign _T_1492 = _T_1290 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@9633.4]
  assign _T_1493 = _T_1492 & _T_696; // @[NV_NVDLA_CDMA_IMG_pack.scala 554:92:@9634.4]
  assign _T_1498 = _T_1296 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@9637.4]
  assign _T_1499 = _T_1487[31:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:102:@9638.4]
  assign _T_1500 = _T_1498 & _T_1499; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:88:@9639.4]
  assign _T_1501 = _T_1493 | _T_1500; // @[NV_NVDLA_CDMA_IMG_pack.scala 554:116:@9640.4]
  assign _T_1506 = _T_1304 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@9643.4]
  assign _T_1507 = _T_1487[63:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:102:@9644.4]
  assign _T_1508 = _T_1506 & _T_1507; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:88:@9645.4]
  assign _T_1509 = _T_1501 | _T_1508; // @[NV_NVDLA_CDMA_IMG_pack.scala 555:150:@9646.4]
  assign _T_1514 = _T_1312 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@9649.4]
  assign _T_1515 = _T_1487[95:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 557:102:@9650.4]
  assign _T_1516 = _T_1514 & _T_1515; // @[NV_NVDLA_CDMA_IMG_pack.scala 557:88:@9651.4]
  assign _T_1517 = _T_1509 | _T_1516; // @[NV_NVDLA_CDMA_IMG_pack.scala 556:189:@9652.4]
  assign _T_1520 = _T_704 & _T_741; // @[NV_NVDLA_CDMA_IMG_pack.scala 558:58:@9655.4]
  assign _GEN_62 = _T_1520 ? _T_1105 : _T_782; // @[NV_NVDLA_CDMA_IMG_pack.scala 563:27:@9666.4]
  assign _GEN_63 = _T_1520 ? _T_696 : _T_791; // @[NV_NVDLA_CDMA_IMG_pack.scala 563:27:@9666.4]
  assign _GEN_69 = _T_734 ? _T_1517 : _T_802; // @[NV_NVDLA_CDMA_IMG_pack.scala 575:24:@9678.4]
  assign _T_1717 = {io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry}; // @[Cat.scala 30:58:@9853.4]
  assign _T_1718 = {io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,_T_1717}; // @[Cat.scala 30:58:@9854.4]
  assign _T_1719 = {io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,io_reg2dp_mean_ry,_T_1717,_T_1718}; // @[Cat.scala 30:58:@9855.4]
  assign _T_1723 = {io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry}; // @[Cat.scala 30:58:@9859.4]
  assign _T_1724 = {io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1723}; // @[Cat.scala 30:58:@9860.4]
  assign _T_1725 = {io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_ax,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1723,_T_1724}; // @[Cat.scala 30:58:@9861.4]
  assign _T_1728 = {io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry}; // @[Cat.scala 30:58:@9864.4]
  assign _T_1729 = {io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1728}; // @[Cat.scala 30:58:@9865.4]
  assign _T_1730 = {io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1728,_T_1729}; // @[Cat.scala 30:58:@9866.4]
  assign _T_1731 = {io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1728,_T_1729,_T_1730}; // @[Cat.scala 30:58:@9867.4]
  assign _T_1732 = {io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,io_reg2dp_mean_bv,io_reg2dp_mean_gu,io_reg2dp_mean_ry,_T_1728,_T_1729,_T_1730,_T_1731}; // @[Cat.scala 30:58:@9868.4]
  assign _T_1734 = io_reg2dp_datain_channel != 13'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:47:@9869.4]
  assign _T_1735 = ~ _T_1734; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:20:@9870.4]
  assign _T_1736 = _T_1735 ? _T_1719 : _T_1725; // @[NV_NVDLA_CDMA_IMG_pack.scala 600:19:@9871.4]
  assign _T_1739 = _T_1736[15:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9873.4]
  assign _T_1740 = _T_813 ? 16'h0 : _T_1739; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9874.4]
  assign _T_1743 = _T_1736[31:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9876.4]
  assign _T_1744 = _T_820 ? 16'h0 : _T_1743; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9877.4]
  assign _T_1747 = _T_1736[47:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9879.4]
  assign _T_1748 = _T_827 ? 16'h0 : _T_1747; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9880.4]
  assign _T_1751 = _T_1736[63:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9882.4]
  assign _T_1752 = _T_834 ? 16'h0 : _T_1751; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9883.4]
  assign _T_1755 = _T_1736[79:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9885.4]
  assign _T_1756 = _T_841 ? 16'h0 : _T_1755; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9886.4]
  assign _T_1759 = _T_1736[95:80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9888.4]
  assign _T_1760 = _T_848 ? 16'h0 : _T_1759; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9889.4]
  assign _T_1763 = _T_1736[111:96]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9891.4]
  assign _T_1764 = _T_855 ? 16'h0 : _T_1763; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9892.4]
  assign _T_1767 = _T_1736[127:112]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9894.4]
  assign _T_1768 = _T_862 ? 16'h0 : _T_1767; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9895.4]
  assign _T_1771 = _T_1736[143:128]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9897.4]
  assign _T_1772 = _T_869 ? 16'h0 : _T_1771; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9898.4]
  assign _T_1775 = _T_1736[159:144]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9900.4]
  assign _T_1776 = _T_876 ? 16'h0 : _T_1775; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9901.4]
  assign _T_1779 = _T_1736[175:160]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9903.4]
  assign _T_1780 = _T_883 ? 16'h0 : _T_1779; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9904.4]
  assign _T_1783 = _T_1736[191:176]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9906.4]
  assign _T_1784 = _T_890 ? 16'h0 : _T_1783; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9907.4]
  assign _T_1787 = _T_1736[207:192]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9909.4]
  assign _T_1788 = _T_897 ? 16'h0 : _T_1787; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9910.4]
  assign _T_1791 = _T_1736[223:208]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9912.4]
  assign _T_1792 = _T_904 ? 16'h0 : _T_1791; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9913.4]
  assign _T_1795 = _T_1736[239:224]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9915.4]
  assign _T_1796 = _T_911 ? 16'h0 : _T_1795; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9916.4]
  assign _T_1799 = _T_1736[255:240]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9918.4]
  assign _T_1800 = _T_918 ? 16'h0 : _T_1799; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9919.4]
  assign _T_1803 = _T_1736[271:256]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9921.4]
  assign _T_1804 = _T_925 ? 16'h0 : _T_1803; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9922.4]
  assign _T_1807 = _T_1736[287:272]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9924.4]
  assign _T_1808 = _T_932 ? 16'h0 : _T_1807; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9925.4]
  assign _T_1811 = _T_1736[303:288]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9927.4]
  assign _T_1812 = _T_939 ? 16'h0 : _T_1811; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9928.4]
  assign _T_1815 = _T_1736[319:304]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9930.4]
  assign _T_1816 = _T_946 ? 16'h0 : _T_1815; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9931.4]
  assign _T_1819 = _T_1736[335:320]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9933.4]
  assign _T_1820 = _T_953 ? 16'h0 : _T_1819; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9934.4]
  assign _T_1823 = _T_1736[351:336]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9936.4]
  assign _T_1824 = _T_960 ? 16'h0 : _T_1823; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9937.4]
  assign _T_1827 = _T_1736[367:352]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9939.4]
  assign _T_1828 = _T_967 ? 16'h0 : _T_1827; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9940.4]
  assign _T_1831 = _T_1736[383:368]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9942.4]
  assign _T_1832 = _T_974 ? 16'h0 : _T_1831; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9943.4]
  assign _T_1835 = _T_1736[399:384]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9945.4]
  assign _T_1836 = _T_981 ? 16'h0 : _T_1835; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9946.4]
  assign _T_1839 = _T_1736[415:400]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9948.4]
  assign _T_1840 = _T_988 ? 16'h0 : _T_1839; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9949.4]
  assign _T_1843 = _T_1736[431:416]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9951.4]
  assign _T_1844 = _T_995 ? 16'h0 : _T_1843; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9952.4]
  assign _T_1847 = _T_1736[447:432]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9954.4]
  assign _T_1848 = _T_1002 ? 16'h0 : _T_1847; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9955.4]
  assign _T_1851 = _T_1736[463:448]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9957.4]
  assign _T_1852 = _T_1009 ? 16'h0 : _T_1851; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9958.4]
  assign _T_1855 = _T_1736[479:464]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9960.4]
  assign _T_1856 = _T_1016 ? 16'h0 : _T_1855; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9961.4]
  assign _T_1859 = _T_1736[495:480]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9963.4]
  assign _T_1860 = _T_1023 ? 16'h0 : _T_1859; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9964.4]
  assign _T_1863 = _T_1736[511:496]; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:55:@9966.4]
  assign _T_1864 = _T_1030 ? 16'h0 : _T_1863; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:13:@9967.4]
  assign _T_1909 = {_T_1768,_T_1764,_T_1760,_T_1756,_T_1752,_T_1748,_T_1744,_T_1740}; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10007.4]
  assign _T_1917 = {_T_1800,_T_1796,_T_1792,_T_1788,_T_1784,_T_1780,_T_1776,_T_1772,_T_1909}; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10015.4]
  assign _T_1924 = {_T_1832,_T_1828,_T_1824,_T_1820,_T_1816,_T_1812,_T_1808,_T_1804}; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10022.4]
  assign _T_1933 = {_T_1864,_T_1860,_T_1856,_T_1852,_T_1848,_T_1844,_T_1840,_T_1836,_T_1924,_T_1917}; // @[NV_NVDLA_CDMA_IMG_pack.scala 602:74:@10031.4]
  assign _T_1934 = _T_1487[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10032.4]
  assign _T_1936 = _T_1732[15:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10033.4]
  assign _T_1937 = _T_1934 ? 16'h0 : _T_1936; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10034.4]
  assign _T_1938 = _T_1487[1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10035.4]
  assign _T_1940 = _T_1732[31:16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10036.4]
  assign _T_1941 = _T_1938 ? 16'h0 : _T_1940; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10037.4]
  assign _T_1942 = _T_1487[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10038.4]
  assign _T_1944 = _T_1732[47:32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10039.4]
  assign _T_1945 = _T_1942 ? 16'h0 : _T_1944; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10040.4]
  assign _T_1946 = _T_1487[3]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10041.4]
  assign _T_1948 = _T_1732[63:48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10042.4]
  assign _T_1949 = _T_1946 ? 16'h0 : _T_1948; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10043.4]
  assign _T_1950 = _T_1487[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10044.4]
  assign _T_1952 = _T_1732[79:64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10045.4]
  assign _T_1953 = _T_1950 ? 16'h0 : _T_1952; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10046.4]
  assign _T_1954 = _T_1487[5]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10047.4]
  assign _T_1956 = _T_1732[95:80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10048.4]
  assign _T_1957 = _T_1954 ? 16'h0 : _T_1956; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10049.4]
  assign _T_1958 = _T_1487[6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10050.4]
  assign _T_1960 = _T_1732[111:96]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10051.4]
  assign _T_1961 = _T_1958 ? 16'h0 : _T_1960; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10052.4]
  assign _T_1962 = _T_1487[7]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10053.4]
  assign _T_1964 = _T_1732[127:112]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10054.4]
  assign _T_1965 = _T_1962 ? 16'h0 : _T_1964; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10055.4]
  assign _T_1966 = _T_1487[8]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10056.4]
  assign _T_1968 = _T_1732[143:128]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10057.4]
  assign _T_1969 = _T_1966 ? 16'h0 : _T_1968; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10058.4]
  assign _T_1970 = _T_1487[9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10059.4]
  assign _T_1972 = _T_1732[159:144]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10060.4]
  assign _T_1973 = _T_1970 ? 16'h0 : _T_1972; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10061.4]
  assign _T_1974 = _T_1487[10]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10062.4]
  assign _T_1976 = _T_1732[175:160]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10063.4]
  assign _T_1977 = _T_1974 ? 16'h0 : _T_1976; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10064.4]
  assign _T_1978 = _T_1487[11]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10065.4]
  assign _T_1980 = _T_1732[191:176]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10066.4]
  assign _T_1981 = _T_1978 ? 16'h0 : _T_1980; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10067.4]
  assign _T_1982 = _T_1487[12]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10068.4]
  assign _T_1984 = _T_1732[207:192]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10069.4]
  assign _T_1985 = _T_1982 ? 16'h0 : _T_1984; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10070.4]
  assign _T_1986 = _T_1487[13]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10071.4]
  assign _T_1988 = _T_1732[223:208]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10072.4]
  assign _T_1989 = _T_1986 ? 16'h0 : _T_1988; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10073.4]
  assign _T_1990 = _T_1487[14]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10074.4]
  assign _T_1992 = _T_1732[239:224]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10075.4]
  assign _T_1993 = _T_1990 ? 16'h0 : _T_1992; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10076.4]
  assign _T_1994 = _T_1487[15]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10077.4]
  assign _T_1996 = _T_1732[255:240]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10078.4]
  assign _T_1997 = _T_1994 ? 16'h0 : _T_1996; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10079.4]
  assign _T_1998 = _T_1487[16]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10080.4]
  assign _T_2000 = _T_1732[271:256]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10081.4]
  assign _T_2001 = _T_1998 ? 16'h0 : _T_2000; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10082.4]
  assign _T_2002 = _T_1487[17]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10083.4]
  assign _T_2004 = _T_1732[287:272]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10084.4]
  assign _T_2005 = _T_2002 ? 16'h0 : _T_2004; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10085.4]
  assign _T_2006 = _T_1487[18]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10086.4]
  assign _T_2008 = _T_1732[303:288]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10087.4]
  assign _T_2009 = _T_2006 ? 16'h0 : _T_2008; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10088.4]
  assign _T_2010 = _T_1487[19]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10089.4]
  assign _T_2012 = _T_1732[319:304]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10090.4]
  assign _T_2013 = _T_2010 ? 16'h0 : _T_2012; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10091.4]
  assign _T_2014 = _T_1487[20]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10092.4]
  assign _T_2016 = _T_1732[335:320]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10093.4]
  assign _T_2017 = _T_2014 ? 16'h0 : _T_2016; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10094.4]
  assign _T_2018 = _T_1487[21]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10095.4]
  assign _T_2020 = _T_1732[351:336]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10096.4]
  assign _T_2021 = _T_2018 ? 16'h0 : _T_2020; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10097.4]
  assign _T_2022 = _T_1487[22]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10098.4]
  assign _T_2024 = _T_1732[367:352]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10099.4]
  assign _T_2025 = _T_2022 ? 16'h0 : _T_2024; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10100.4]
  assign _T_2026 = _T_1487[23]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10101.4]
  assign _T_2028 = _T_1732[383:368]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10102.4]
  assign _T_2029 = _T_2026 ? 16'h0 : _T_2028; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10103.4]
  assign _T_2030 = _T_1487[24]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10104.4]
  assign _T_2032 = _T_1732[399:384]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10105.4]
  assign _T_2033 = _T_2030 ? 16'h0 : _T_2032; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10106.4]
  assign _T_2034 = _T_1487[25]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10107.4]
  assign _T_2036 = _T_1732[415:400]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10108.4]
  assign _T_2037 = _T_2034 ? 16'h0 : _T_2036; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10109.4]
  assign _T_2038 = _T_1487[26]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10110.4]
  assign _T_2040 = _T_1732[431:416]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10111.4]
  assign _T_2041 = _T_2038 ? 16'h0 : _T_2040; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10112.4]
  assign _T_2042 = _T_1487[27]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10113.4]
  assign _T_2044 = _T_1732[447:432]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10114.4]
  assign _T_2045 = _T_2042 ? 16'h0 : _T_2044; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10115.4]
  assign _T_2046 = _T_1487[28]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10116.4]
  assign _T_2048 = _T_1732[463:448]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10117.4]
  assign _T_2049 = _T_2046 ? 16'h0 : _T_2048; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10118.4]
  assign _T_2050 = _T_1487[29]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10119.4]
  assign _T_2052 = _T_1732[479:464]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10120.4]
  assign _T_2053 = _T_2050 ? 16'h0 : _T_2052; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10121.4]
  assign _T_2054 = _T_1487[30]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10122.4]
  assign _T_2056 = _T_1732[495:480]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10123.4]
  assign _T_2057 = _T_2054 ? 16'h0 : _T_2056; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10124.4]
  assign _T_2058 = _T_1487[31]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10125.4]
  assign _T_2060 = _T_1732[511:496]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10126.4]
  assign _T_2061 = _T_2058 ? 16'h0 : _T_2060; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10127.4]
  assign _T_2062 = _T_1487[32]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10128.4]
  assign _T_2064 = _T_1732[527:512]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10129.4]
  assign _T_2065 = _T_2062 ? 16'h0 : _T_2064; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10130.4]
  assign _T_2066 = _T_1487[33]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10131.4]
  assign _T_2068 = _T_1732[543:528]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10132.4]
  assign _T_2069 = _T_2066 ? 16'h0 : _T_2068; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10133.4]
  assign _T_2070 = _T_1487[34]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10134.4]
  assign _T_2072 = _T_1732[559:544]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10135.4]
  assign _T_2073 = _T_2070 ? 16'h0 : _T_2072; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10136.4]
  assign _T_2074 = _T_1487[35]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10137.4]
  assign _T_2076 = _T_1732[575:560]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10138.4]
  assign _T_2077 = _T_2074 ? 16'h0 : _T_2076; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10139.4]
  assign _T_2078 = _T_1487[36]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10140.4]
  assign _T_2080 = _T_1732[591:576]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10141.4]
  assign _T_2081 = _T_2078 ? 16'h0 : _T_2080; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10142.4]
  assign _T_2082 = _T_1487[37]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10143.4]
  assign _T_2084 = _T_1732[607:592]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10144.4]
  assign _T_2085 = _T_2082 ? 16'h0 : _T_2084; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10145.4]
  assign _T_2086 = _T_1487[38]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10146.4]
  assign _T_2088 = _T_1732[623:608]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10147.4]
  assign _T_2089 = _T_2086 ? 16'h0 : _T_2088; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10148.4]
  assign _T_2090 = _T_1487[39]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10149.4]
  assign _T_2092 = _T_1732[639:624]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10150.4]
  assign _T_2093 = _T_2090 ? 16'h0 : _T_2092; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10151.4]
  assign _T_2094 = _T_1487[40]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10152.4]
  assign _T_2096 = _T_1732[655:640]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10153.4]
  assign _T_2097 = _T_2094 ? 16'h0 : _T_2096; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10154.4]
  assign _T_2098 = _T_1487[41]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10155.4]
  assign _T_2100 = _T_1732[671:656]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10156.4]
  assign _T_2101 = _T_2098 ? 16'h0 : _T_2100; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10157.4]
  assign _T_2102 = _T_1487[42]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10158.4]
  assign _T_2104 = _T_1732[687:672]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10159.4]
  assign _T_2105 = _T_2102 ? 16'h0 : _T_2104; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10160.4]
  assign _T_2106 = _T_1487[43]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10161.4]
  assign _T_2108 = _T_1732[703:688]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10162.4]
  assign _T_2109 = _T_2106 ? 16'h0 : _T_2108; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10163.4]
  assign _T_2110 = _T_1487[44]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10164.4]
  assign _T_2112 = _T_1732[719:704]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10165.4]
  assign _T_2113 = _T_2110 ? 16'h0 : _T_2112; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10166.4]
  assign _T_2114 = _T_1487[45]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10167.4]
  assign _T_2116 = _T_1732[735:720]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10168.4]
  assign _T_2117 = _T_2114 ? 16'h0 : _T_2116; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10169.4]
  assign _T_2118 = _T_1487[46]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10170.4]
  assign _T_2120 = _T_1732[751:736]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10171.4]
  assign _T_2121 = _T_2118 ? 16'h0 : _T_2120; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10172.4]
  assign _T_2122 = _T_1487[47]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10173.4]
  assign _T_2124 = _T_1732[767:752]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10174.4]
  assign _T_2125 = _T_2122 ? 16'h0 : _T_2124; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10175.4]
  assign _T_2126 = _T_1487[48]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10176.4]
  assign _T_2128 = _T_1732[783:768]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10177.4]
  assign _T_2129 = _T_2126 ? 16'h0 : _T_2128; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10178.4]
  assign _T_2130 = _T_1487[49]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10179.4]
  assign _T_2132 = _T_1732[799:784]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10180.4]
  assign _T_2133 = _T_2130 ? 16'h0 : _T_2132; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10181.4]
  assign _T_2134 = _T_1487[50]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10182.4]
  assign _T_2136 = _T_1732[815:800]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10183.4]
  assign _T_2137 = _T_2134 ? 16'h0 : _T_2136; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10184.4]
  assign _T_2138 = _T_1487[51]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10185.4]
  assign _T_2140 = _T_1732[831:816]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10186.4]
  assign _T_2141 = _T_2138 ? 16'h0 : _T_2140; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10187.4]
  assign _T_2142 = _T_1487[52]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10188.4]
  assign _T_2144 = _T_1732[847:832]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10189.4]
  assign _T_2145 = _T_2142 ? 16'h0 : _T_2144; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10190.4]
  assign _T_2146 = _T_1487[53]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10191.4]
  assign _T_2148 = _T_1732[863:848]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10192.4]
  assign _T_2149 = _T_2146 ? 16'h0 : _T_2148; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10193.4]
  assign _T_2150 = _T_1487[54]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10194.4]
  assign _T_2152 = _T_1732[879:864]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10195.4]
  assign _T_2153 = _T_2150 ? 16'h0 : _T_2152; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10196.4]
  assign _T_2154 = _T_1487[55]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10197.4]
  assign _T_2156 = _T_1732[895:880]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10198.4]
  assign _T_2157 = _T_2154 ? 16'h0 : _T_2156; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10199.4]
  assign _T_2158 = _T_1487[56]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10200.4]
  assign _T_2160 = _T_1732[911:896]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10201.4]
  assign _T_2161 = _T_2158 ? 16'h0 : _T_2160; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10202.4]
  assign _T_2162 = _T_1487[57]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10203.4]
  assign _T_2164 = _T_1732[927:912]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10204.4]
  assign _T_2165 = _T_2162 ? 16'h0 : _T_2164; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10205.4]
  assign _T_2166 = _T_1487[58]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10206.4]
  assign _T_2168 = _T_1732[943:928]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10207.4]
  assign _T_2169 = _T_2166 ? 16'h0 : _T_2168; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10208.4]
  assign _T_2170 = _T_1487[59]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10209.4]
  assign _T_2172 = _T_1732[959:944]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10210.4]
  assign _T_2173 = _T_2170 ? 16'h0 : _T_2172; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10211.4]
  assign _T_2174 = _T_1487[60]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10212.4]
  assign _T_2176 = _T_1732[975:960]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10213.4]
  assign _T_2177 = _T_2174 ? 16'h0 : _T_2176; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10214.4]
  assign _T_2178 = _T_1487[61]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10215.4]
  assign _T_2180 = _T_1732[991:976]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10216.4]
  assign _T_2181 = _T_2178 ? 16'h0 : _T_2180; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10217.4]
  assign _T_2182 = _T_1487[62]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10218.4]
  assign _T_2184 = _T_1732[1007:992]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10219.4]
  assign _T_2185 = _T_2182 ? 16'h0 : _T_2184; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10220.4]
  assign _T_2186 = _T_1487[63]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10221.4]
  assign _T_2188 = _T_1732[1023:1008]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10222.4]
  assign _T_2189 = _T_2186 ? 16'h0 : _T_2188; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10223.4]
  assign _T_2190 = _T_1487[64]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10224.4]
  assign _T_2192 = _T_1732[1039:1024]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10225.4]
  assign _T_2193 = _T_2190 ? 16'h0 : _T_2192; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10226.4]
  assign _T_2194 = _T_1487[65]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10227.4]
  assign _T_2196 = _T_1732[1055:1040]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10228.4]
  assign _T_2197 = _T_2194 ? 16'h0 : _T_2196; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10229.4]
  assign _T_2198 = _T_1487[66]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10230.4]
  assign _T_2200 = _T_1732[1071:1056]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10231.4]
  assign _T_2201 = _T_2198 ? 16'h0 : _T_2200; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10232.4]
  assign _T_2202 = _T_1487[67]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10233.4]
  assign _T_2204 = _T_1732[1087:1072]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10234.4]
  assign _T_2205 = _T_2202 ? 16'h0 : _T_2204; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10235.4]
  assign _T_2206 = _T_1487[68]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10236.4]
  assign _T_2208 = _T_1732[1103:1088]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10237.4]
  assign _T_2209 = _T_2206 ? 16'h0 : _T_2208; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10238.4]
  assign _T_2210 = _T_1487[69]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10239.4]
  assign _T_2212 = _T_1732[1119:1104]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10240.4]
  assign _T_2213 = _T_2210 ? 16'h0 : _T_2212; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10241.4]
  assign _T_2214 = _T_1487[70]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10242.4]
  assign _T_2216 = _T_1732[1135:1120]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10243.4]
  assign _T_2217 = _T_2214 ? 16'h0 : _T_2216; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10244.4]
  assign _T_2218 = _T_1487[71]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10245.4]
  assign _T_2220 = _T_1732[1151:1136]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10246.4]
  assign _T_2221 = _T_2218 ? 16'h0 : _T_2220; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10247.4]
  assign _T_2222 = _T_1487[72]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10248.4]
  assign _T_2224 = _T_1732[1167:1152]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10249.4]
  assign _T_2225 = _T_2222 ? 16'h0 : _T_2224; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10250.4]
  assign _T_2226 = _T_1487[73]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10251.4]
  assign _T_2228 = _T_1732[1183:1168]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10252.4]
  assign _T_2229 = _T_2226 ? 16'h0 : _T_2228; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10253.4]
  assign _T_2230 = _T_1487[74]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10254.4]
  assign _T_2232 = _T_1732[1199:1184]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10255.4]
  assign _T_2233 = _T_2230 ? 16'h0 : _T_2232; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10256.4]
  assign _T_2234 = _T_1487[75]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10257.4]
  assign _T_2236 = _T_1732[1215:1200]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10258.4]
  assign _T_2237 = _T_2234 ? 16'h0 : _T_2236; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10259.4]
  assign _T_2238 = _T_1487[76]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10260.4]
  assign _T_2240 = _T_1732[1231:1216]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10261.4]
  assign _T_2241 = _T_2238 ? 16'h0 : _T_2240; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10262.4]
  assign _T_2242 = _T_1487[77]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10263.4]
  assign _T_2244 = _T_1732[1247:1232]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10264.4]
  assign _T_2245 = _T_2242 ? 16'h0 : _T_2244; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10265.4]
  assign _T_2246 = _T_1487[78]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10266.4]
  assign _T_2248 = _T_1732[1263:1248]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10267.4]
  assign _T_2249 = _T_2246 ? 16'h0 : _T_2248; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10268.4]
  assign _T_2250 = _T_1487[79]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10269.4]
  assign _T_2252 = _T_1732[1279:1264]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10270.4]
  assign _T_2253 = _T_2250 ? 16'h0 : _T_2252; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10271.4]
  assign _T_2254 = _T_1487[80]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10272.4]
  assign _T_2256 = _T_1732[1295:1280]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10273.4]
  assign _T_2257 = _T_2254 ? 16'h0 : _T_2256; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10274.4]
  assign _T_2258 = _T_1487[81]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10275.4]
  assign _T_2260 = _T_1732[1311:1296]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10276.4]
  assign _T_2261 = _T_2258 ? 16'h0 : _T_2260; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10277.4]
  assign _T_2262 = _T_1487[82]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10278.4]
  assign _T_2264 = _T_1732[1327:1312]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10279.4]
  assign _T_2265 = _T_2262 ? 16'h0 : _T_2264; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10280.4]
  assign _T_2266 = _T_1487[83]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10281.4]
  assign _T_2268 = _T_1732[1343:1328]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10282.4]
  assign _T_2269 = _T_2266 ? 16'h0 : _T_2268; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10283.4]
  assign _T_2270 = _T_1487[84]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10284.4]
  assign _T_2272 = _T_1732[1359:1344]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10285.4]
  assign _T_2273 = _T_2270 ? 16'h0 : _T_2272; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10286.4]
  assign _T_2274 = _T_1487[85]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10287.4]
  assign _T_2276 = _T_1732[1375:1360]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10288.4]
  assign _T_2277 = _T_2274 ? 16'h0 : _T_2276; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10289.4]
  assign _T_2278 = _T_1487[86]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10290.4]
  assign _T_2280 = _T_1732[1391:1376]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10291.4]
  assign _T_2281 = _T_2278 ? 16'h0 : _T_2280; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10292.4]
  assign _T_2282 = _T_1487[87]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10293.4]
  assign _T_2284 = _T_1732[1407:1392]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10294.4]
  assign _T_2285 = _T_2282 ? 16'h0 : _T_2284; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10295.4]
  assign _T_2286 = _T_1487[88]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10296.4]
  assign _T_2288 = _T_1732[1423:1408]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10297.4]
  assign _T_2289 = _T_2286 ? 16'h0 : _T_2288; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10298.4]
  assign _T_2290 = _T_1487[89]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10299.4]
  assign _T_2292 = _T_1732[1439:1424]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10300.4]
  assign _T_2293 = _T_2290 ? 16'h0 : _T_2292; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10301.4]
  assign _T_2294 = _T_1487[90]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10302.4]
  assign _T_2296 = _T_1732[1455:1440]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10303.4]
  assign _T_2297 = _T_2294 ? 16'h0 : _T_2296; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10304.4]
  assign _T_2298 = _T_1487[91]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10305.4]
  assign _T_2300 = _T_1732[1471:1456]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10306.4]
  assign _T_2301 = _T_2298 ? 16'h0 : _T_2300; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10307.4]
  assign _T_2302 = _T_1487[92]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10308.4]
  assign _T_2304 = _T_1732[1487:1472]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10309.4]
  assign _T_2305 = _T_2302 ? 16'h0 : _T_2304; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10310.4]
  assign _T_2306 = _T_1487[93]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10311.4]
  assign _T_2308 = _T_1732[1503:1488]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10312.4]
  assign _T_2309 = _T_2306 ? 16'h0 : _T_2308; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10313.4]
  assign _T_2310 = _T_1487[94]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10314.4]
  assign _T_2312 = _T_1732[1519:1504]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10315.4]
  assign _T_2313 = _T_2310 ? 16'h0 : _T_2312; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10316.4]
  assign _T_2314 = _T_1487[95]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:25:@10317.4]
  assign _T_2316 = _T_1732[1535:1520]; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:55:@10318.4]
  assign _T_2317 = _T_2314 ? 16'h0 : _T_2316; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:13:@10319.4]
  assign _T_2424 = {_T_1957,_T_1953,_T_1949,_T_1945,_T_1941,_T_1937}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10421.4]
  assign _T_2430 = {_T_1981,_T_1977,_T_1973,_T_1969,_T_1965,_T_1961,_T_2424}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10427.4]
  assign _T_2435 = {_T_2005,_T_2001,_T_1997,_T_1993,_T_1989,_T_1985}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10432.4]
  assign _T_2442 = {_T_2029,_T_2025,_T_2021,_T_2017,_T_2013,_T_2009,_T_2435,_T_2430}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10439.4]
  assign _T_2447 = {_T_2053,_T_2049,_T_2045,_T_2041,_T_2037,_T_2033}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10444.4]
  assign _T_2453 = {_T_2077,_T_2073,_T_2069,_T_2065,_T_2061,_T_2057,_T_2447}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10450.4]
  assign _T_2458 = {_T_2101,_T_2097,_T_2093,_T_2089,_T_2085,_T_2081}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10455.4]
  assign _T_2466 = {_T_2125,_T_2121,_T_2117,_T_2113,_T_2109,_T_2105,_T_2458,_T_2453,_T_2442}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10463.4]
  assign _T_2471 = {_T_2149,_T_2145,_T_2141,_T_2137,_T_2133,_T_2129}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10468.4]
  assign _T_2477 = {_T_2173,_T_2169,_T_2165,_T_2161,_T_2157,_T_2153,_T_2471}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10474.4]
  assign _T_2482 = {_T_2197,_T_2193,_T_2189,_T_2185,_T_2181,_T_2177}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10479.4]
  assign _T_2489 = {_T_2221,_T_2217,_T_2213,_T_2209,_T_2205,_T_2201,_T_2482,_T_2477}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10486.4]
  assign _T_2494 = {_T_2245,_T_2241,_T_2237,_T_2233,_T_2229,_T_2225}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10491.4]
  assign _T_2500 = {_T_2269,_T_2265,_T_2261,_T_2257,_T_2253,_T_2249,_T_2494}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10497.4]
  assign _T_2505 = {_T_2293,_T_2289,_T_2285,_T_2281,_T_2277,_T_2273}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10502.4]
  assign _T_2514 = {_T_2317,_T_2313,_T_2309,_T_2305,_T_2301,_T_2297,_T_2505,_T_2500,_T_2489,_T_2466}; // @[NV_NVDLA_CDMA_IMG_pack.scala 604:74:@10511.4]
  assign _T_2519 = io_pixel_precision != 2'h0; // @[NV_NVDLA_CDMA_IMG_pack.scala 606:87:@10514.4]
  assign _T_2520 = _T_1276 & _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 606:66:@10515.4]
  assign _T_2526 = ~ _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 607:68:@10519.4]
  assign _T_2527 = _T_1276 & _T_2526; // @[NV_NVDLA_CDMA_IMG_pack.scala 607:66:@10520.4]
  assign _T_2533 = _T_1279 & _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 608:66:@10524.4]
  assign _T_2540 = _T_1279 & _T_2526; // @[NV_NVDLA_CDMA_IMG_pack.scala 609:66:@10529.4]
  assign _T_2546 = _T_1282 & _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 610:66:@10533.4]
  assign _T_2553 = _T_1282 & _T_2526; // @[NV_NVDLA_CDMA_IMG_pack.scala 611:66:@10538.4]
  assign _T_2559 = _T_1285 & _T_2519; // @[NV_NVDLA_CDMA_IMG_pack.scala 612:65:@10543.4]
  assign _T_2564 = io_pixel_packed_10b | _T_2526; // @[NV_NVDLA_CDMA_IMG_pack.scala 613:65:@10547.4]
  assign _T_2565 = _T_249 & _T_2564; // @[NV_NVDLA_CDMA_IMG_pack.scala 613:42:@10548.4]
  assign _T_2572 = {_T_2520,_T_2527,_T_2533,_T_2540,_T_2546,_T_2553,_T_2559,_T_2565}; // @[Cat.scala 30:58:@10555.4]
  assign _T_2573 = _T_2572[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:56:@10556.4]
  assign _T_2577 = _T_2573 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@10558.4]
  assign _T_2578 = _T_2577 & _T_1933; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:60:@10559.4]
  assign _T_2579 = _T_2572[2]; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:56:@10560.4]
  assign _T_2583 = _T_2579 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@10562.4]
  assign _T_2584 = _T_2514[511:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:71:@10563.4]
  assign _T_2585 = _T_2583 & _T_2584; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:60:@10564.4]
  assign _T_2586 = _T_2578 | _T_2585; // @[NV_NVDLA_CDMA_IMG_pack.scala 615:73:@10565.4]
  assign _T_2587 = _T_2572[4]; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:56:@10566.4]
  assign _T_2591 = _T_2587 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@10568.4]
  assign _T_2592 = _T_2514[1023:512]; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:71:@10569.4]
  assign _T_2593 = _T_2591 & _T_2592; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:60:@10570.4]
  assign _T_2594 = _T_2586 | _T_2593; // @[NV_NVDLA_CDMA_IMG_pack.scala 616:89:@10571.4]
  assign _T_2595 = _T_2572[6]; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:56:@10572.4]
  assign _T_2599 = _T_2595 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@10574.4]
  assign _T_2600 = _T_2514[1535:1024]; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:71:@10575.4]
  assign _T_2601 = _T_2599 & _T_2600; // @[NV_NVDLA_CDMA_IMG_pack.scala 618:60:@10576.4]
  assign _T_2602 = _T_2594 | _T_2601; // @[NV_NVDLA_CDMA_IMG_pack.scala 617:100:@10577.4]
  assign _T_2606 = _T_2526 | io_pixel_packed_10b; // @[NV_NVDLA_CDMA_IMG_pack.scala 623:72:@10582.4]
  assign _T_2607 = _T_734 & _T_2606; // @[NV_NVDLA_CDMA_IMG_pack.scala 623:43:@10583.4]
  assign _GEN_73 = _T_2607 ? _T_2602 : {{256'd0}, _T_1542}; // @[NV_NVDLA_CDMA_IMG_pack.scala 634:27:@10593.4]
  assign _T_2611 = _T_740 ? io_sg2pack_entry_end : io_sg2pack_entry_mid; // @[NV_NVDLA_CDMA_IMG_pack.scala 647:28:@10597.4]
  assign _T_2612 = _T_739 ? io_sg2pack_entry_st : _T_2611; // @[NV_NVDLA_CDMA_IMG_pack.scala 646:28:@10598.4]
  assign _T_2613 = _T_740 ? io_sg2pack_sub_h_end : io_sg2pack_sub_h_mid; // @[NV_NVDLA_CDMA_IMG_pack.scala 649:28:@10599.4]
  assign _T_2614 = _T_739 ? io_sg2pack_sub_h_st : _T_2613; // @[NV_NVDLA_CDMA_IMG_pack.scala 648:27:@10600.4]
  assign _T_2616 = {1'h0,io_status2dma_wr_idx}; // @[Cat.scala 30:58:@10601.4]
  assign _T_2617 = _T_2610 + _T_2612; // @[NV_NVDLA_CDMA_IMG_pack.scala 650:99:@10602.4]
  assign _T_2618 = _T_123 ? _T_2616 : _T_2617; // @[NV_NVDLA_CDMA_IMG_pack.scala 650:29:@10603.4]
  assign _T_2619 = _T_2618[15:9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:38:@10604.4]
  assign _GEN_91 = {{1'd0}, io_pixel_bank}; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:76:@10605.4]
  assign _T_2620 = _T_2619 >= _GEN_91; // @[NV_NVDLA_CDMA_IMG_pack.scala 652:76:@10605.4]
  assign _T_2627 = {io_pixel_bank,9'h0}; // @[Cat.scala 30:58:@10608.4]
  assign _GEN_92 = {{1'd0}, _T_2627}; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10609.4]
  assign _T_2628 = _T_2618 - _GEN_92; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10609.4]
  assign _T_2629 = $unsigned(_T_2628); // @[NV_NVDLA_CDMA_IMG_pack.scala 653:54:@10610.4]
  assign _T_2630 = _T_2629[14:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 653:124:@10611.4]
  assign _T_2631 = _T_2618[14:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 654:81:@10612.4]
  assign _T_2632 = _T_2620 ? _T_2630 : _T_2631; // @[NV_NVDLA_CDMA_IMG_pack.scala 654:27:@10613.4]
  assign _T_2633 = _T_734 & _T_738; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:59:@10614.4]
  assign _T_2634 = _T_2633 & _T_736; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:85:@10615.4]
  assign _T_2635 = _T_123 | _T_2634; // @[NV_NVDLA_CDMA_IMG_pack.scala 656:42:@10616.4]
  assign _GEN_74 = _T_2635 ? _T_2632 : _T_2610; // @[NV_NVDLA_CDMA_IMG_pack.scala 658:24:@10617.4]
  assign _T_2639 = _T_123 | _T_736; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:49:@10621.4]
  assign _T_2641 = _T_2638 + io_sg2pack_data_entries; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:111:@10622.4]
  assign _T_2642 = _T_2638 + io_sg2pack_data_entries; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:111:@10623.4]
  assign _T_2643 = _T_2639 ? 15'h0 : _T_2642; // @[NV_NVDLA_CDMA_IMG_pack.scala 665:31:@10624.4]
  assign _T_2644 = _T_734 & _T_737; // @[NV_NVDLA_CDMA_IMG_pack.scala 666:63:@10625.4]
  assign _T_2645 = _T_123 | _T_2644; // @[NV_NVDLA_CDMA_IMG_pack.scala 666:46:@10626.4]
  assign _GEN_75 = _T_2645 ? _T_2643 : _T_2638; // @[NV_NVDLA_CDMA_IMG_pack.scala 668:28:@10627.4]
  assign _T_2652 = _T_738 & _T_736; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:77:@10632.4]
  assign _T_2653 = _T_123 | _T_2652; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:50:@10633.4]
  assign _T_2655 = ~ _T_736; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:54:@10634.4]
  assign _T_2656 = _T_737 & _T_2655; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:52:@10635.4]
  assign _T_2657 = _T_2648 + 15'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:120:@10636.4]
  assign _T_2658 = _T_2648 + 15'h1; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:120:@10637.4]
  assign _T_2659 = _T_2656 ? _T_2651 : _T_2658; // @[NV_NVDLA_CDMA_IMG_pack.scala 677:31:@10638.4]
  assign _T_2660 = _T_2653 ? 15'h0 : _T_2659; // @[NV_NVDLA_CDMA_IMG_pack.scala 676:31:@10639.4]
  assign _T_2661 = _T_123 | _T_734; // @[NV_NVDLA_CDMA_IMG_pack.scala 679:46:@10640.4]
  assign _GEN_76 = _T_2661 ? _T_2660 : _T_2648; // @[NV_NVDLA_CDMA_IMG_pack.scala 682:28:@10641.4]
  assign _GEN_77 = _T_123 ? _T_2660 : _T_2651; // @[NV_NVDLA_CDMA_IMG_pack.scala 685:32:@10644.4]
  assign _T_2665 = _T_2610 + _T_2638; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:41:@10648.4]
  assign _T_2666 = _T_2648[14:1]; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:84:@10649.4]
  assign _GEN_93 = {{2'd0}, _T_2666}; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:63:@10650.4]
  assign _T_2667 = _T_2665 + _GEN_93; // @[NV_NVDLA_CDMA_IMG_pack.scala 691:63:@10650.4]
  assign _T_2668 = _T_2648[0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 692:63:@10651.4]
  assign _GEN_78 = _T_734 ? _T_2668 : _T_2664; // @[NV_NVDLA_CDMA_IMG_pack.scala 697:32:@10652.4]
  assign _T_2673 = _T_2667[16:9]; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:38:@10657.4]
  assign _GEN_94 = {{2'd0}, io_pixel_bank}; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:76:@10658.4]
  assign _T_2674 = _T_2673 >= _GEN_94; // @[NV_NVDLA_CDMA_IMG_pack.scala 712:76:@10658.4]
  assign _GEN_95 = {{2'd0}, _T_2627}; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10662.4]
  assign _T_2682 = _T_2667 - _GEN_95; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10662.4]
  assign _T_2683 = $unsigned(_T_2682); // @[NV_NVDLA_CDMA_IMG_pack.scala 713:54:@10663.4]
  assign _T_2684 = _T_2683[14:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 713:124:@10664.4]
  assign _T_2685 = _T_2667[14:0]; // @[NV_NVDLA_CDMA_IMG_pack.scala 714:79:@10665.4]
  assign _T_2686 = _T_2674 ? _T_2684 : _T_2685; // @[NV_NVDLA_CDMA_IMG_pack.scala 714:25:@10666.4]
  assign _GEN_79 = _T_734 ? _T_2686 : _T_2672; // @[NV_NVDLA_CDMA_IMG_pack.scala 717:20:@10667.4]
  assign _GEN_80 = _T_2634 ? _T_2612 : _T_2692; // @[NV_NVDLA_CDMA_IMG_pack.scala 731:23:@10676.4]
  assign _GEN_81 = _T_2634 ? _T_2614 : _T_2695; // @[NV_NVDLA_CDMA_IMG_pack.scala 731:23:@10676.4]
  assign _T_2704 = _T_734 & _T_740; // @[NV_NVDLA_CDMA_IMG_pack.scala 760:40:@10692.4]
  assign _T_2706 = _T_2704 ? 1'h1 : _T_2702; // @[NV_NVDLA_CDMA_IMG_pack.scala 760:25:@10693.4]
  assign _T_2707 = _T_123 ? 1'h0 : _T_2706; // @[NV_NVDLA_CDMA_IMG_pack.scala 759:25:@10694.4]
  assign io_img2sbuf_p0_rd_addr_valid = _T_354; // @[NV_NVDLA_CDMA_IMG_pack.scala 372:30:@8869.4]
  assign io_img2sbuf_p0_rd_addr_bits = _T_373; // @[NV_NVDLA_CDMA_IMG_pack.scala 373:29:@8870.4]
  assign io_sg2pack_img_pd_ready = _T_283 & _T_303; // @[NV_NVDLA_CDMA_IMG_pack.scala 195:25:@8592.4]
  assign io_img2cvt_dat_wr_sel = _T_2664; // @[NV_NVDLA_CDMA_IMG_pack.scala 747:31:@10686.4]
  assign io_img2cvt_dat_wr_addr_valid = _T_758; // @[NV_NVDLA_CDMA_IMG_pack.scala 743:30:@10684.4]
  assign io_img2cvt_dat_wr_addr_bits = {{2'd0}, _T_2672}; // @[NV_NVDLA_CDMA_IMG_pack.scala 749:29:@10687.4]
  assign io_img2cvt_dat_wr_data = _T_799; // @[NV_NVDLA_CDMA_IMG_pack.scala 750:24:@10688.4]
  assign io_img2cvt_mn_wr_data = {{256'd0}, _T_1542}; // @[NV_NVDLA_CDMA_IMG_pack.scala 751:23:@10689.4]
  assign io_img2cvt_dat_wr_pad_mask = _T_802; // @[NV_NVDLA_CDMA_IMG_pack.scala 752:28:@10690.4]
  assign io_img2cvt_dat_wr_info_pd = {_T_778,_T_775}; // @[NV_NVDLA_CDMA_IMG_pack.scala 744:27:@10685.4]
  assign io_img2status_dat_updt_valid = _T_2689; // @[NV_NVDLA_CDMA_IMG_pack.scala 739:30:@10680.4]
  assign io_img2status_dat_updt_bits_entries = _T_2692; // @[NV_NVDLA_CDMA_IMG_pack.scala 741:37:@10683.4]
  assign io_img2status_dat_updt_bits_slices = {10'h0,_T_2695}; // @[NV_NVDLA_CDMA_IMG_pack.scala 740:36:@10682.4]
  assign io_pack_is_done = _T_2702; // @[NV_NVDLA_CDMA_IMG_pack.scala 764:17:@10696.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_115 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_126 = _RAND_1[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_132 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_142 = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_145 = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_148 = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_151 = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_154 = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_157 = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_160 = _RAND_10[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_163 = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_218 = _RAND_12[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_281 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_257 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_246 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_234 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_337 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_354 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_358 = _RAND_19[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_361 = _RAND_20[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_370 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_373 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_409 = _RAND_23[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_412 = _RAND_24[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_450 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_452 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_604 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_607 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_610 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_613 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_616 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_619 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_622 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_631 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_634 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_639 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_642 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_647 = _RAND_38[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_650 = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_655 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_658 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_663 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_666 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_671 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_674 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_679 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_682 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_687 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_690 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_694 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_696 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_700 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_702 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_709 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_712 = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_715 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_718 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_721 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_724 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_727 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_730 = _RAND_61[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_758 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_761 = _RAND_63[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_764 = _RAND_64[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_767 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_770 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {8{`RANDOM}};
  _T_782 = _RAND_67[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {8{`RANDOM}};
  _T_785 = _RAND_68[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {8{`RANDOM}};
  _T_788 = _RAND_69[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_791 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_794 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_797 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {8{`RANDOM}};
  _T_799 = _RAND_73[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_802 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {8{`RANDOM}};
  _T_1542 = _RAND_75[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_2610 = _RAND_76[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_2638 = _RAND_77[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_2648 = _RAND_78[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_2651 = _RAND_79[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_2664 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_2672 = _RAND_81[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_2689 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_2692 = _RAND_83[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_2695 = _RAND_84[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_2702 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_115 <= 1'h0;
    end else begin
      _T_115 <= io_is_running;
    end
    if (reset) begin
      _T_126 <= 14'h0;
    end else begin
      if (io_layer_st) begin
        _T_126 <= {{9'd0}, io_reg2dp_pad_left};
      end
    end
    if (reset) begin
      _T_129 <= 14'h0;
    end else begin
      _T_129 <= _GEN_1[13:0];
    end
    if (reset) begin
      _T_132 <= 14'h0;
    end else begin
      _T_132 <= _GEN_2[13:0];
    end
    if (reset) begin
      _T_142 <= 5'h0;
    end else begin
      _T_142 <= _GEN_3[4:0];
    end
    if (reset) begin
      _T_145 <= 5'h0;
    end else begin
      _T_145 <= _GEN_4[4:0];
    end
    if (reset) begin
      _T_148 <= 5'h0;
    end else begin
      _T_148 <= _GEN_5[4:0];
    end
    if (reset) begin
      _T_151 <= 5'h0;
    end else begin
      _T_151 <= _GEN_6[4:0];
    end
    if (reset) begin
      _T_154 <= 5'h0;
    end else begin
      _T_154 <= _GEN_7[4:0];
    end
    if (reset) begin
      _T_157 <= 5'h0;
    end else begin
      _T_157 <= _GEN_8[4:0];
    end
    if (reset) begin
      _T_160 <= 6'h0;
    end else begin
      _T_160 <= _GEN_9[5:0];
    end
    if (reset) begin
      _T_163 <= 6'h0;
    end else begin
      _T_163 <= _GEN_10[5:0];
    end
    if (reset) begin
      _T_218 <= 13'h0;
    end else begin
      if (_T_316) begin
        if (_T_123) begin
          _T_218 <= 13'h0;
        end else begin
          _T_218 <= _T_227;
        end
      end
    end
    if (reset) begin
      _T_281 <= 1'h0;
    end else begin
      if (_T_284) begin
        _T_281 <= 1'h0;
      end else begin
        if (_T_303) begin
          _T_281 <= 1'h0;
        end else begin
          if (io_sg2pack_img_pd_valid) begin
            _T_281 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_257 <= 2'h0;
    end else begin
      if (_T_312) begin
        if (_T_269) begin
          _T_257 <= 2'h0;
        end else begin
          _T_257 <= _T_273;
        end
      end
    end
    if (reset) begin
      _T_246 <= 1'h0;
    end else begin
      if (_T_314) begin
        if (_T_251) begin
          _T_246 <= 1'h0;
        end else begin
          _T_246 <= _T_253;
        end
      end
    end
    if (reset) begin
      _T_234 <= 4'h0;
    end else begin
      if (_T_315) begin
        if (_T_241) begin
          _T_234 <= 4'h0;
        end else begin
          _T_234 <= _T_239;
        end
      end
    end
    if (reset) begin
      _T_337 <= 1'h0;
    end else begin
      _T_337 <= _T_283;
    end
    if (reset) begin
      _T_354 <= 1'h0;
    end else begin
      _T_354 <= _T_283;
    end
    if (reset) begin
      _T_358 <= 7'h0;
    end else begin
      if (_T_404) begin
        if (_T_123) begin
          _T_358 <= 7'h0;
        end else begin
          _T_358 <= _T_383;
        end
      end
    end
    if (reset) begin
      _T_361 <= 7'h0;
    end else begin
      if (_T_406) begin
        if (_T_123) begin
          _T_361 <= 7'h0;
        end else begin
          _T_361 <= _T_385;
        end
      end
    end
    if (reset) begin
      _T_370 <= 8'h0;
    end else begin
      if (_T_253) begin
        _T_370 <= _T_395;
      end else begin
        _T_370 <= _T_400;
      end
    end
    if (reset) begin
      _T_373 <= 8'h0;
    end else begin
      if (_T_283) begin
        _T_373 <= _T_370;
      end
    end
    if (reset) begin
      _T_409 <= 14'h0;
    end else begin
      if (_T_404) begin
        if (_T_431) begin
          _T_409 <= 14'h0;
        end else begin
          _T_409 <= _T_414;
        end
      end
    end
    if (reset) begin
      _T_412 <= 14'h0;
    end else begin
      if (_T_406) begin
        if (_T_434) begin
          _T_412 <= 14'h0;
        end else begin
          _T_412 <= _T_416;
        end
      end
    end
    if (_T_283) begin
      if (_T_253) begin
        _T_450 <= _T_440;
      end else begin
        _T_450 <= _T_444;
      end
    end
    if (_T_283) begin
      if (_T_253) begin
        _T_452 <= _T_440;
      end else begin
        _T_452 <= _T_444;
      end
    end
    if (reset) begin
      _T_604 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_604 <= _T_246;
      end
    end
    if (reset) begin
      _T_607 <= 3'h0;
    end else begin
      if (_T_283) begin
        _T_607 <= 3'h0;
      end
    end
    if (reset) begin
      _T_610 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_610 <= _T_303;
      end
    end
    if (reset) begin
      _T_613 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_613 <= _T_303;
      end
    end
    if (reset) begin
      _T_616 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_616 <= _T_625;
      end
    end
    if (reset) begin
      _T_619 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_619 <= _T_223;
      end
    end
    if (reset) begin
      _T_622 <= 1'h0;
    end else begin
      if (_T_283) begin
        _T_622 <= _T_626;
      end
    end
    if (reset) begin
      _T_631 <= 1'h0;
    end else begin
      _T_631 <= _T_337;
    end
    if (reset) begin
      _T_634 <= 1'h0;
    end else begin
      _T_634 <= _T_631;
    end
    if (reset) begin
      _T_639 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_639 <= _T_604;
      end
    end
    if (reset) begin
      _T_642 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_642 <= _T_639;
      end
    end
    if (reset) begin
      _T_647 <= 3'h0;
    end else begin
      if (_T_337) begin
        _T_647 <= _T_607;
      end
    end
    if (reset) begin
      _T_650 <= 3'h0;
    end else begin
      if (_T_631) begin
        _T_650 <= _T_647;
      end
    end
    if (reset) begin
      _T_655 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_655 <= _T_610;
      end
    end
    if (reset) begin
      _T_658 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_658 <= _T_655;
      end
    end
    if (reset) begin
      _T_663 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_663 <= _T_613;
      end
    end
    if (reset) begin
      _T_666 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_666 <= _T_663;
      end
    end
    if (reset) begin
      _T_671 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_671 <= _T_616;
      end
    end
    if (reset) begin
      _T_674 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_674 <= _T_671;
      end
    end
    if (reset) begin
      _T_679 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_679 <= _T_619;
      end
    end
    if (reset) begin
      _T_682 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_682 <= _T_679;
      end
    end
    if (reset) begin
      _T_687 <= 1'h0;
    end else begin
      if (_T_337) begin
        _T_687 <= _T_622;
      end
    end
    if (reset) begin
      _T_690 <= 1'h0;
    end else begin
      if (_T_631) begin
        _T_690 <= _T_687;
      end
    end
    if (_T_337) begin
      _T_694 <= _T_452;
    end
    if (_T_631) begin
      _T_696 <= _T_694;
    end
    if (_T_337) begin
      _T_700 <= _T_450;
    end
    if (_T_631) begin
      _T_702 <= _T_700;
    end
    if (reset) begin
      _T_709 <= 1'h0;
    end else begin
      _T_709 <= _T_706;
    end
    if (reset) begin
      _T_712 <= 3'h0;
    end else begin
      if (_T_706) begin
        _T_712 <= _T_650;
      end
    end
    if (reset) begin
      _T_715 <= 1'h0;
    end else begin
      if (_T_706) begin
        _T_715 <= _T_658;
      end
    end
    if (reset) begin
      _T_718 <= 1'h0;
    end else begin
      if (_T_706) begin
        _T_718 <= _T_666;
      end
    end
    if (reset) begin
      _T_721 <= 1'h0;
    end else begin
      if (_T_706) begin
        _T_721 <= _T_674;
      end
    end
    if (reset) begin
      _T_724 <= 1'h0;
    end else begin
      if (_T_706) begin
        _T_724 <= _T_682;
      end
    end
    if (reset) begin
      _T_727 <= 1'h0;
    end else begin
      if (_T_706) begin
        _T_727 <= _T_690;
      end
    end
    if (reset) begin
      _T_730 <= 2'h0;
    end else begin
      if (_T_634) begin
        if (_T_742) begin
          _T_730 <= 2'h0;
        end else begin
          _T_730 <= _T_746;
        end
      end
    end
    if (reset) begin
      _T_758 <= 1'h0;
    end else begin
      if (_T_733) begin
        _T_758 <= _T_634;
      end else begin
        _T_758 <= _T_709;
      end
    end
    if (reset) begin
      _T_761 <= 3'h0;
    end else begin
      if (_T_734) begin
        if (_T_733) begin
          _T_761 <= _T_650;
        end else begin
          _T_761 <= _T_712;
        end
      end
    end
    if (reset) begin
      _T_764 <= 4'h0;
    end else begin
      if (_T_123) begin
        _T_764 <= 4'h1;
      end
    end
    if (reset) begin
      _T_767 <= 1'h0;
    end else begin
      if (_T_123) begin
        _T_767 <= io_sg2pack_mn_enable;
      end
    end
    if (reset) begin
      _T_770 <= 1'h0;
    end else begin
      if (_T_123) begin
        _T_770 <= io_pixel_uint;
      end
    end
    if (reset) begin
      _T_782 <= 256'h0;
    end else begin
      if (_T_1520) begin
        _T_782 <= _T_1105;
      end
    end
    if (reset) begin
      _T_785 <= 256'h0;
    end else begin
      if (_T_1525) begin
        _T_785 <= _T_1105;
      end
    end
    if (reset) begin
      _T_788 <= 256'h0;
    end else begin
      if (_T_1530) begin
        _T_788 <= _T_1105;
      end
    end
    if (reset) begin
      _T_791 <= 32'h0;
    end else begin
      if (_T_1520) begin
        _T_791 <= _T_696;
      end
    end
    if (reset) begin
      _T_794 <= 32'h0;
    end else begin
      if (_T_1525) begin
        _T_794 <= _T_696;
      end
    end
    if (reset) begin
      _T_797 <= 32'h0;
    end else begin
      if (_T_1530) begin
        _T_797 <= _T_696;
      end
    end
    if (_T_734) begin
      _T_799 <= _T_1319;
    end
    if (reset) begin
      _T_802 <= 32'h0;
    end else begin
      if (_T_734) begin
        _T_802 <= _T_1517;
      end
    end
    if (reset) begin
      _T_1542 <= 256'h0;
    end else begin
      _T_1542 <= _GEN_73[255:0];
    end
    if (reset) begin
      _T_2610 <= 15'h0;
    end else begin
      if (_T_2635) begin
        if (_T_2620) begin
          _T_2610 <= _T_2630;
        end else begin
          _T_2610 <= _T_2631;
        end
      end
    end
    if (reset) begin
      _T_2638 <= 15'h0;
    end else begin
      if (_T_2645) begin
        if (_T_2639) begin
          _T_2638 <= 15'h0;
        end else begin
          _T_2638 <= _T_2642;
        end
      end
    end
    if (reset) begin
      _T_2648 <= 15'h0;
    end else begin
      if (_T_2661) begin
        if (_T_2653) begin
          _T_2648 <= 15'h0;
        end else begin
          if (_T_2656) begin
            _T_2648 <= _T_2651;
          end else begin
            _T_2648 <= _T_2658;
          end
        end
      end
    end
    if (reset) begin
      _T_2651 <= 15'h0;
    end else begin
      if (_T_123) begin
        if (_T_2653) begin
          _T_2651 <= 15'h0;
        end else begin
          if (!(_T_2656)) begin
            _T_2651 <= _T_2658;
          end
        end
      end
    end
    if (reset) begin
      _T_2664 <= 1'h0;
    end else begin
      if (_T_734) begin
        _T_2664 <= _T_2668;
      end
    end
    if (reset) begin
      _T_2672 <= 15'h0;
    end else begin
      if (_T_734) begin
        if (_T_2674) begin
          _T_2672 <= _T_2684;
        end else begin
          _T_2672 <= _T_2685;
        end
      end
    end
    if (reset) begin
      _T_2689 <= 1'h0;
    end else begin
      _T_2689 <= _T_2634;
    end
    if (reset) begin
      _T_2692 <= 15'h0;
    end else begin
      if (_T_2634) begin
        if (_T_739) begin
          _T_2692 <= io_sg2pack_entry_st;
        end else begin
          if (_T_740) begin
            _T_2692 <= io_sg2pack_entry_end;
          end else begin
            _T_2692 <= io_sg2pack_entry_mid;
          end
        end
      end
    end
    if (reset) begin
      _T_2695 <= 4'h0;
    end else begin
      if (_T_2634) begin
        if (_T_739) begin
          _T_2695 <= io_sg2pack_sub_h_st;
        end else begin
          if (_T_740) begin
            _T_2695 <= io_sg2pack_sub_h_end;
          end else begin
            _T_2695 <= io_sg2pack_sub_h_mid;
          end
        end
      end
    end
    if (reset) begin
      _T_2702 <= 1'h1;
    end else begin
      if (_T_123) begin
        _T_2702 <= 1'h0;
      end else begin
        if (_T_2704) begin
          _T_2702 <= 1'h1;
        end
      end
    end
  end
endmodule
module NV_NVDLA_CDMA_img( // @[:@10698.2]
  input          reset, // @[:@10700.4]
  input          io_nvdla_core_clk, // @[:@10701.4]
  input          io_nvdla_core_ng_clk, // @[:@10701.4]
  input          io_img_dat2mcif_rd_req_pd_ready, // @[:@10701.4]
  output         io_img_dat2mcif_rd_req_pd_valid, // @[:@10701.4]
  output [78:0]  io_img_dat2mcif_rd_req_pd_bits, // @[:@10701.4]
  output         io_mcif2img_dat_rd_rsp_pd_ready, // @[:@10701.4]
  input          io_mcif2img_dat_rd_rsp_pd_valid, // @[:@10701.4]
  input  [256:0] io_mcif2img_dat_rd_rsp_pd_bits, // @[:@10701.4]
  input          io_img_dat2cvif_rd_req_pd_ready, // @[:@10701.4]
  output         io_img_dat2cvif_rd_req_pd_valid, // @[:@10701.4]
  output [78:0]  io_img_dat2cvif_rd_req_pd_bits, // @[:@10701.4]
  output         io_cvif2img_dat_rd_rsp_pd_ready, // @[:@10701.4]
  input          io_cvif2img_dat_rd_rsp_pd_valid, // @[:@10701.4]
  input  [256:0] io_cvif2img_dat_rd_rsp_pd_bits, // @[:@10701.4]
  output         io_img2cvt_dat_wr_sel, // @[:@10701.4]
  output         io_img2cvt_dat_wr_addr_valid, // @[:@10701.4]
  output [16:0]  io_img2cvt_dat_wr_addr_bits, // @[:@10701.4]
  output [255:0] io_img2cvt_dat_wr_data, // @[:@10701.4]
  output [511:0] io_img2cvt_mn_wr_data, // @[:@10701.4]
  output [31:0]  io_img2cvt_dat_wr_pad_mask, // @[:@10701.4]
  output [11:0]  io_img2cvt_dat_wr_info_pd, // @[:@10701.4]
  output [1:0]   io_img2status_state, // @[:@10701.4]
  output         io_img2status_dat_updt_valid, // @[:@10701.4]
  output [14:0]  io_img2status_dat_updt_bits_entries, // @[:@10701.4]
  output [13:0]  io_img2status_dat_updt_bits_slices, // @[:@10701.4]
  input  [14:0]  io_status2dma_free_entries, // @[:@10701.4]
  input  [14:0]  io_status2dma_wr_idx, // @[:@10701.4]
  input          io_status2dma_fsm_switch, // @[:@10701.4]
  output         io_img2sbuf_p0_wr_addr_valid, // @[:@10701.4]
  output [7:0]   io_img2sbuf_p0_wr_addr_bits, // @[:@10701.4]
  output [255:0] io_img2sbuf_p0_wr_data, // @[:@10701.4]
  output         io_img2sbuf_p0_rd_addr_valid, // @[:@10701.4]
  output [7:0]   io_img2sbuf_p0_rd_addr_bits, // @[:@10701.4]
  input  [255:0] io_img2sbuf_p0_rd_data, // @[:@10701.4]
  input          io_sc2cdma_dat_pending_req, // @[:@10701.4]
  input          io_reg2dp_op_en, // @[:@10701.4]
  input          io_reg2dp_conv_mode, // @[:@10701.4]
  input          io_reg2dp_data_reuse, // @[:@10701.4]
  input          io_reg2dp_skip_data_rls, // @[:@10701.4]
  input          io_reg2dp_datain_format, // @[:@10701.4]
  input  [5:0]   io_reg2dp_pixel_format, // @[:@10701.4]
  input          io_reg2dp_pixel_sign_override, // @[:@10701.4]
  input  [12:0]  io_reg2dp_datain_width, // @[:@10701.4]
  input  [12:0]  io_reg2dp_datain_height, // @[:@10701.4]
  input  [12:0]  io_reg2dp_datain_channel, // @[:@10701.4]
  input  [4:0]   io_reg2dp_pixel_x_offset, // @[:@10701.4]
  input          io_reg2dp_datain_ram_type, // @[:@10701.4]
  input  [31:0]  io_reg2dp_datain_addr_high_0, // @[:@10701.4]
  input  [31:0]  io_reg2dp_datain_addr_low_0, // @[:@10701.4]
  input  [31:0]  io_reg2dp_datain_addr_low_1, // @[:@10701.4]
  input  [31:0]  io_reg2dp_line_stride, // @[:@10701.4]
  input  [31:0]  io_reg2dp_uv_line_stride, // @[:@10701.4]
  input  [31:0]  io_reg2dp_datain_addr_high_1, // @[:@10701.4]
  input          io_reg2dp_mean_format, // @[:@10701.4]
  input  [15:0]  io_reg2dp_mean_ry, // @[:@10701.4]
  input  [15:0]  io_reg2dp_mean_gu, // @[:@10701.4]
  input  [15:0]  io_reg2dp_mean_bv, // @[:@10701.4]
  input  [15:0]  io_reg2dp_mean_ax, // @[:@10701.4]
  input  [13:0]  io_reg2dp_entries, // @[:@10701.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@10701.4]
  input  [5:0]   io_reg2dp_pad_right, // @[:@10701.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@10701.4]
  input          io_reg2dp_dma_en, // @[:@10701.4]
  output [31:0]  io_dp2reg_img_rd_stall, // @[:@10701.4]
  output [31:0]  io_dp2reg_img_rd_latency // @[:@10701.4]
);
  wire  u_ctrl_reset; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_nvdla_core_ng_clk; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pack_is_done; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_sg_is_done; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [1:0] u_ctrl_io_img2status_state; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_is_running; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_layer_st; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [5:0] u_ctrl_io_pixel_bank; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_early_end; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [10:0] u_ctrl_io_pixel_order; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_packed_10b; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_planar; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [1:0] u_ctrl_io_pixel_precision; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_uint; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [3:0] u_ctrl_io_pixel_planar0_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [3:0] u_ctrl_io_pixel_planar0_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_pixel_planar0_byte_sft; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [3:0] u_ctrl_io_pixel_planar0_lp_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_planar0_lp_vld; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [3:0] u_ctrl_io_pixel_planar0_rp_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_planar0_rp_vld; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [2:0] u_ctrl_io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [13:0] u_ctrl_io_pixel_planar0_width_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_pixel_planar1_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_pixel_planar1_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_pixel_planar1_byte_sft; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [2:0] u_ctrl_io_pixel_planar1_lp_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_planar1_lp_vld; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [2:0] u_ctrl_io_pixel_planar1_rp_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_pixel_planar1_rp_vld; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [2:0] u_ctrl_io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [13:0] u_ctrl_io_pixel_planar1_width_burst; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_op_en; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_conv_mode; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_datain_format; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [5:0] u_ctrl_io_reg2dp_pixel_format; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_pixel_sign_override; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [12:0] u_ctrl_io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_data_reuse; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_ctrl_io_reg2dp_skip_data_rls; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_reg2dp_data_bank; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_reg2dp_pixel_x_offset; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [4:0] u_ctrl_io_reg2dp_pad_left; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire [5:0] u_ctrl_io_reg2dp_pad_right; // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
  wire  u_sg_reset; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [78:0] u_sg_io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [256:0] u_sg_io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [78:0] u_sg_io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [256:0] u_sg_io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_img2status_dat_entries; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img2status_dat_updt; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_status2dma_free_entries; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_status2dma_fsm_switch; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_is_running; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_layer_st; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [10:0] u_sg_io_pixel_order; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_pixel_planar; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_pixel_planar0_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_pixel_planar0_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [4:0] u_sg_io_pixel_planar0_byte_sft; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [4:0] u_sg_io_pixel_planar1_byte_sft; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_pixel_planar0_lp_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_pixel_planar0_lp_vld; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_pixel_planar0_rp_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_pixel_planar0_rp_vld; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [13:0] u_sg_io_pixel_planar0_width_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [4:0] u_sg_io_pixel_planar1_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [4:0] u_sg_io_pixel_planar1_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [2:0] u_sg_io_pixel_planar1_lp_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_pixel_planar1_lp_vld; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [2:0] u_sg_io_pixel_planar1_rp_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_pixel_planar1_rp_vld; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [13:0] u_sg_io_pixel_planar1_width_burst; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_sg2pack_img_pd_ready; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_sg2pack_img_pd_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [10:0] u_sg_io_sg2pack_img_pd_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_sg2pack_data_entries; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_sg2pack_entry_end; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_sg2pack_entry_mid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [14:0] u_sg_io_sg2pack_entry_st; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [12:0] u_sg_io_sg2pack_height_total; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_sg2pack_mn_enable; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_sg2pack_sub_h_end; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_sg2pack_sub_h_mid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [3:0] u_sg_io_sg2pack_sub_h_st; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_sg_is_done; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_img2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [16:0] u_sg_io_img2sbuf_p0_wr_addr_bits; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [255:0] u_sg_io_img2sbuf_p0_wr_data; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_reg2dp_op_en; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [12:0] u_sg_io_reg2dp_datain_height; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_reg2dp_datain_ram_type; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_datain_addr_high_0; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_datain_addr_low_0; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_datain_addr_high_1; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_datain_addr_low_1; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_line_stride; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_reg2dp_uv_line_stride; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_reg2dp_mean_format; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [13:0] u_sg_io_reg2dp_entries; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_sg_io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_dp2reg_img_rd_stall; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire [31:0] u_sg_io_dp2reg_img_rd_latency; // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
  wire  u_pack_reset; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_img2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [7:0] u_pack_io_img2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [255:0] u_pack_io_img2sbuf_p0_rd_data; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_is_running; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_layer_st; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [5:0] u_pack_io_pixel_bank; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_pixel_early_end; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_pixel_packed_10b; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_pixel_planar; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [2:0] u_pack_io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [2:0] u_pack_io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [1:0] u_pack_io_pixel_precision; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_pixel_uint; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_sg2pack_img_pd_ready; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_sg2pack_img_pd_valid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [10:0] u_pack_io_sg2pack_img_pd_bits; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_sg2pack_data_entries; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_sg2pack_entry_end; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_sg2pack_entry_mid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_sg2pack_entry_st; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [12:0] u_pack_io_sg2pack_height_total; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_sg2pack_mn_enable; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [3:0] u_pack_io_sg2pack_sub_h_end; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [3:0] u_pack_io_sg2pack_sub_h_mid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [3:0] u_pack_io_sg2pack_sub_h_st; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_status2dma_wr_idx; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_img2cvt_dat_wr_sel; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [16:0] u_pack_io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [255:0] u_pack_io_img2cvt_dat_wr_data; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [511:0] u_pack_io_img2cvt_mn_wr_data; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [31:0] u_pack_io_img2cvt_dat_wr_pad_mask; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [11:0] u_pack_io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_img2status_dat_updt_valid; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [14:0] u_pack_io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [13:0] u_pack_io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire  u_pack_io_pack_is_done; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [12:0] u_pack_io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [12:0] u_pack_io_reg2dp_datain_channel; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [15:0] u_pack_io_reg2dp_mean_ry; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [15:0] u_pack_io_reg2dp_mean_gu; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [15:0] u_pack_io_reg2dp_mean_bv; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [15:0] u_pack_io_reg2dp_mean_ax; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [4:0] u_pack_io_reg2dp_pad_left; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  wire [5:0] u_pack_io_reg2dp_pad_right; // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
  NV_NVDLA_CDMA_IMG_ctrl u_ctrl ( // @[NV_NVDLA_CDMA_img.scala 107:24:@10703.4]
    .reset(u_ctrl_reset),
    .io_nvdla_core_clk(u_ctrl_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(u_ctrl_io_nvdla_core_ng_clk),
    .io_pack_is_done(u_ctrl_io_pack_is_done),
    .io_sc2cdma_dat_pending_req(u_ctrl_io_sc2cdma_dat_pending_req),
    .io_sg_is_done(u_ctrl_io_sg_is_done),
    .io_img2status_state(u_ctrl_io_img2status_state),
    .io_is_running(u_ctrl_io_is_running),
    .io_layer_st(u_ctrl_io_layer_st),
    .io_pixel_bank(u_ctrl_io_pixel_bank),
    .io_pixel_early_end(u_ctrl_io_pixel_early_end),
    .io_pixel_order(u_ctrl_io_pixel_order),
    .io_pixel_packed_10b(u_ctrl_io_pixel_packed_10b),
    .io_pixel_planar(u_ctrl_io_pixel_planar),
    .io_pixel_precision(u_ctrl_io_pixel_precision),
    .io_pixel_uint(u_ctrl_io_pixel_uint),
    .io_pixel_planar0_bundle_limit(u_ctrl_io_pixel_planar0_bundle_limit),
    .io_pixel_planar0_bundle_limit_1st(u_ctrl_io_pixel_planar0_bundle_limit_1st),
    .io_pixel_planar0_byte_sft(u_ctrl_io_pixel_planar0_byte_sft),
    .io_pixel_planar0_lp_burst(u_ctrl_io_pixel_planar0_lp_burst),
    .io_pixel_planar0_lp_vld(u_ctrl_io_pixel_planar0_lp_vld),
    .io_pixel_planar0_rp_burst(u_ctrl_io_pixel_planar0_rp_burst),
    .io_pixel_planar0_rp_vld(u_ctrl_io_pixel_planar0_rp_vld),
    .io_pixel_planar0_sft(u_ctrl_io_pixel_planar0_sft),
    .io_pixel_planar0_width_burst(u_ctrl_io_pixel_planar0_width_burst),
    .io_pixel_planar1_bundle_limit(u_ctrl_io_pixel_planar1_bundle_limit),
    .io_pixel_planar1_bundle_limit_1st(u_ctrl_io_pixel_planar1_bundle_limit_1st),
    .io_pixel_planar1_byte_sft(u_ctrl_io_pixel_planar1_byte_sft),
    .io_pixel_planar1_lp_burst(u_ctrl_io_pixel_planar1_lp_burst),
    .io_pixel_planar1_lp_vld(u_ctrl_io_pixel_planar1_lp_vld),
    .io_pixel_planar1_rp_burst(u_ctrl_io_pixel_planar1_rp_burst),
    .io_pixel_planar1_rp_vld(u_ctrl_io_pixel_planar1_rp_vld),
    .io_pixel_planar1_sft(u_ctrl_io_pixel_planar1_sft),
    .io_pixel_planar1_width_burst(u_ctrl_io_pixel_planar1_width_burst),
    .io_reg2dp_op_en(u_ctrl_io_reg2dp_op_en),
    .io_reg2dp_conv_mode(u_ctrl_io_reg2dp_conv_mode),
    .io_reg2dp_datain_format(u_ctrl_io_reg2dp_datain_format),
    .io_reg2dp_pixel_format(u_ctrl_io_reg2dp_pixel_format),
    .io_reg2dp_pixel_sign_override(u_ctrl_io_reg2dp_pixel_sign_override),
    .io_reg2dp_datain_width(u_ctrl_io_reg2dp_datain_width),
    .io_reg2dp_data_reuse(u_ctrl_io_reg2dp_data_reuse),
    .io_reg2dp_skip_data_rls(u_ctrl_io_reg2dp_skip_data_rls),
    .io_reg2dp_data_bank(u_ctrl_io_reg2dp_data_bank),
    .io_reg2dp_pixel_x_offset(u_ctrl_io_reg2dp_pixel_x_offset),
    .io_reg2dp_pad_left(u_ctrl_io_reg2dp_pad_left),
    .io_reg2dp_pad_right(u_ctrl_io_reg2dp_pad_right)
  );
  NV_NVDLA_CDMA_IMG_sg u_sg ( // @[NV_NVDLA_CDMA_img.scala 134:22:@10728.4]
    .reset(u_sg_reset),
    .io_nvdla_core_clk(u_sg_io_nvdla_core_clk),
    .io_img_dat2mcif_rd_req_pd_ready(u_sg_io_img_dat2mcif_rd_req_pd_ready),
    .io_img_dat2mcif_rd_req_pd_valid(u_sg_io_img_dat2mcif_rd_req_pd_valid),
    .io_img_dat2mcif_rd_req_pd_bits(u_sg_io_img_dat2mcif_rd_req_pd_bits),
    .io_mcif2img_dat_rd_rsp_pd_ready(u_sg_io_mcif2img_dat_rd_rsp_pd_ready),
    .io_mcif2img_dat_rd_rsp_pd_valid(u_sg_io_mcif2img_dat_rd_rsp_pd_valid),
    .io_mcif2img_dat_rd_rsp_pd_bits(u_sg_io_mcif2img_dat_rd_rsp_pd_bits),
    .io_img_dat2cvif_rd_req_pd_ready(u_sg_io_img_dat2cvif_rd_req_pd_ready),
    .io_img_dat2cvif_rd_req_pd_valid(u_sg_io_img_dat2cvif_rd_req_pd_valid),
    .io_img_dat2cvif_rd_req_pd_bits(u_sg_io_img_dat2cvif_rd_req_pd_bits),
    .io_cvif2img_dat_rd_rsp_pd_ready(u_sg_io_cvif2img_dat_rd_rsp_pd_ready),
    .io_cvif2img_dat_rd_rsp_pd_valid(u_sg_io_cvif2img_dat_rd_rsp_pd_valid),
    .io_cvif2img_dat_rd_rsp_pd_bits(u_sg_io_cvif2img_dat_rd_rsp_pd_bits),
    .io_img2status_dat_entries(u_sg_io_img2status_dat_entries),
    .io_img2status_dat_updt(u_sg_io_img2status_dat_updt),
    .io_status2dma_free_entries(u_sg_io_status2dma_free_entries),
    .io_status2dma_fsm_switch(u_sg_io_status2dma_fsm_switch),
    .io_is_running(u_sg_io_is_running),
    .io_layer_st(u_sg_io_layer_st),
    .io_pixel_order(u_sg_io_pixel_order),
    .io_pixel_planar(u_sg_io_pixel_planar),
    .io_pixel_planar0_bundle_limit(u_sg_io_pixel_planar0_bundle_limit),
    .io_pixel_planar0_bundle_limit_1st(u_sg_io_pixel_planar0_bundle_limit_1st),
    .io_pixel_planar0_byte_sft(u_sg_io_pixel_planar0_byte_sft),
    .io_pixel_planar1_byte_sft(u_sg_io_pixel_planar1_byte_sft),
    .io_pixel_planar0_lp_burst(u_sg_io_pixel_planar0_lp_burst),
    .io_pixel_planar0_lp_vld(u_sg_io_pixel_planar0_lp_vld),
    .io_pixel_planar0_rp_burst(u_sg_io_pixel_planar0_rp_burst),
    .io_pixel_planar0_rp_vld(u_sg_io_pixel_planar0_rp_vld),
    .io_pixel_planar0_width_burst(u_sg_io_pixel_planar0_width_burst),
    .io_pixel_planar1_bundle_limit(u_sg_io_pixel_planar1_bundle_limit),
    .io_pixel_planar1_bundle_limit_1st(u_sg_io_pixel_planar1_bundle_limit_1st),
    .io_pixel_planar1_lp_burst(u_sg_io_pixel_planar1_lp_burst),
    .io_pixel_planar1_lp_vld(u_sg_io_pixel_planar1_lp_vld),
    .io_pixel_planar1_rp_burst(u_sg_io_pixel_planar1_rp_burst),
    .io_pixel_planar1_rp_vld(u_sg_io_pixel_planar1_rp_vld),
    .io_pixel_planar1_width_burst(u_sg_io_pixel_planar1_width_burst),
    .io_sg2pack_img_pd_ready(u_sg_io_sg2pack_img_pd_ready),
    .io_sg2pack_img_pd_valid(u_sg_io_sg2pack_img_pd_valid),
    .io_sg2pack_img_pd_bits(u_sg_io_sg2pack_img_pd_bits),
    .io_sg2pack_data_entries(u_sg_io_sg2pack_data_entries),
    .io_sg2pack_entry_end(u_sg_io_sg2pack_entry_end),
    .io_sg2pack_entry_mid(u_sg_io_sg2pack_entry_mid),
    .io_sg2pack_entry_st(u_sg_io_sg2pack_entry_st),
    .io_sg2pack_height_total(u_sg_io_sg2pack_height_total),
    .io_sg2pack_mn_enable(u_sg_io_sg2pack_mn_enable),
    .io_sg2pack_sub_h_end(u_sg_io_sg2pack_sub_h_end),
    .io_sg2pack_sub_h_mid(u_sg_io_sg2pack_sub_h_mid),
    .io_sg2pack_sub_h_st(u_sg_io_sg2pack_sub_h_st),
    .io_sg_is_done(u_sg_io_sg_is_done),
    .io_img2sbuf_p0_wr_addr_valid(u_sg_io_img2sbuf_p0_wr_addr_valid),
    .io_img2sbuf_p0_wr_addr_bits(u_sg_io_img2sbuf_p0_wr_addr_bits),
    .io_img2sbuf_p0_wr_data(u_sg_io_img2sbuf_p0_wr_data),
    .io_reg2dp_op_en(u_sg_io_reg2dp_op_en),
    .io_reg2dp_datain_height(u_sg_io_reg2dp_datain_height),
    .io_reg2dp_datain_ram_type(u_sg_io_reg2dp_datain_ram_type),
    .io_reg2dp_datain_addr_high_0(u_sg_io_reg2dp_datain_addr_high_0),
    .io_reg2dp_datain_addr_low_0(u_sg_io_reg2dp_datain_addr_low_0),
    .io_reg2dp_datain_addr_high_1(u_sg_io_reg2dp_datain_addr_high_1),
    .io_reg2dp_datain_addr_low_1(u_sg_io_reg2dp_datain_addr_low_1),
    .io_reg2dp_line_stride(u_sg_io_reg2dp_line_stride),
    .io_reg2dp_uv_line_stride(u_sg_io_reg2dp_uv_line_stride),
    .io_reg2dp_mean_format(u_sg_io_reg2dp_mean_format),
    .io_reg2dp_entries(u_sg_io_reg2dp_entries),
    .io_reg2dp_dma_en(u_sg_io_reg2dp_dma_en),
    .io_dp2reg_img_rd_stall(u_sg_io_dp2reg_img_rd_stall),
    .io_dp2reg_img_rd_latency(u_sg_io_dp2reg_img_rd_latency)
  );
  NV_NVDLA_CDMA_IMG_pack u_pack ( // @[NV_NVDLA_CDMA_img.scala 191:24:@10788.4]
    .reset(u_pack_reset),
    .io_nvdla_core_clk(u_pack_io_nvdla_core_clk),
    .io_img2sbuf_p0_rd_addr_valid(u_pack_io_img2sbuf_p0_rd_addr_valid),
    .io_img2sbuf_p0_rd_addr_bits(u_pack_io_img2sbuf_p0_rd_addr_bits),
    .io_img2sbuf_p0_rd_data(u_pack_io_img2sbuf_p0_rd_data),
    .io_is_running(u_pack_io_is_running),
    .io_layer_st(u_pack_io_layer_st),
    .io_pixel_bank(u_pack_io_pixel_bank),
    .io_pixel_early_end(u_pack_io_pixel_early_end),
    .io_pixel_packed_10b(u_pack_io_pixel_packed_10b),
    .io_pixel_planar(u_pack_io_pixel_planar),
    .io_pixel_planar0_sft(u_pack_io_pixel_planar0_sft),
    .io_pixel_planar1_sft(u_pack_io_pixel_planar1_sft),
    .io_pixel_precision(u_pack_io_pixel_precision),
    .io_pixel_uint(u_pack_io_pixel_uint),
    .io_sg2pack_img_pd_ready(u_pack_io_sg2pack_img_pd_ready),
    .io_sg2pack_img_pd_valid(u_pack_io_sg2pack_img_pd_valid),
    .io_sg2pack_img_pd_bits(u_pack_io_sg2pack_img_pd_bits),
    .io_sg2pack_data_entries(u_pack_io_sg2pack_data_entries),
    .io_sg2pack_entry_end(u_pack_io_sg2pack_entry_end),
    .io_sg2pack_entry_mid(u_pack_io_sg2pack_entry_mid),
    .io_sg2pack_entry_st(u_pack_io_sg2pack_entry_st),
    .io_sg2pack_height_total(u_pack_io_sg2pack_height_total),
    .io_sg2pack_mn_enable(u_pack_io_sg2pack_mn_enable),
    .io_sg2pack_sub_h_end(u_pack_io_sg2pack_sub_h_end),
    .io_sg2pack_sub_h_mid(u_pack_io_sg2pack_sub_h_mid),
    .io_sg2pack_sub_h_st(u_pack_io_sg2pack_sub_h_st),
    .io_status2dma_wr_idx(u_pack_io_status2dma_wr_idx),
    .io_img2cvt_dat_wr_sel(u_pack_io_img2cvt_dat_wr_sel),
    .io_img2cvt_dat_wr_addr_valid(u_pack_io_img2cvt_dat_wr_addr_valid),
    .io_img2cvt_dat_wr_addr_bits(u_pack_io_img2cvt_dat_wr_addr_bits),
    .io_img2cvt_dat_wr_data(u_pack_io_img2cvt_dat_wr_data),
    .io_img2cvt_mn_wr_data(u_pack_io_img2cvt_mn_wr_data),
    .io_img2cvt_dat_wr_pad_mask(u_pack_io_img2cvt_dat_wr_pad_mask),
    .io_img2cvt_dat_wr_info_pd(u_pack_io_img2cvt_dat_wr_info_pd),
    .io_img2status_dat_updt_valid(u_pack_io_img2status_dat_updt_valid),
    .io_img2status_dat_updt_bits_entries(u_pack_io_img2status_dat_updt_bits_entries),
    .io_img2status_dat_updt_bits_slices(u_pack_io_img2status_dat_updt_bits_slices),
    .io_pack_is_done(u_pack_io_pack_is_done),
    .io_reg2dp_datain_width(u_pack_io_reg2dp_datain_width),
    .io_reg2dp_datain_channel(u_pack_io_reg2dp_datain_channel),
    .io_reg2dp_mean_ry(u_pack_io_reg2dp_mean_ry),
    .io_reg2dp_mean_gu(u_pack_io_reg2dp_mean_gu),
    .io_reg2dp_mean_bv(u_pack_io_reg2dp_mean_bv),
    .io_reg2dp_mean_ax(u_pack_io_reg2dp_mean_ax),
    .io_reg2dp_pad_left(u_pack_io_reg2dp_pad_left),
    .io_reg2dp_pad_right(u_pack_io_reg2dp_pad_right)
  );
  assign io_img_dat2mcif_rd_req_pd_valid = u_sg_io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_img.scala 141:31:@10739.4]
  assign io_img_dat2mcif_rd_req_pd_bits = u_sg_io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_img.scala 141:31:@10738.4]
  assign io_mcif2img_dat_rd_rsp_pd_ready = u_sg_io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_img.scala 142:36:@10743.4]
  assign io_img_dat2cvif_rd_req_pd_valid = u_sg_io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_img.scala 138:39:@10733.4]
  assign io_img_dat2cvif_rd_req_pd_bits = u_sg_io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_img.scala 138:39:@10732.4]
  assign io_cvif2img_dat_rd_rsp_pd_ready = u_sg_io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_img.scala 139:44:@10737.4]
  assign io_img2cvt_dat_wr_sel = u_pack_io_img2cvt_dat_wr_sel; // @[NV_NVDLA_CDMA_img.scala 223:35:@10820.4]
  assign io_img2cvt_dat_wr_addr_valid = u_pack_io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_CDMA_img.scala 225:23:@10823.4]
  assign io_img2cvt_dat_wr_addr_bits = u_pack_io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_CDMA_img.scala 225:23:@10822.4]
  assign io_img2cvt_dat_wr_data = u_pack_io_img2cvt_dat_wr_data; // @[NV_NVDLA_CDMA_img.scala 225:23:@10821.4]
  assign io_img2cvt_mn_wr_data = u_pack_io_img2cvt_mn_wr_data; // @[NV_NVDLA_CDMA_img.scala 226:27:@10824.4]
  assign io_img2cvt_dat_wr_pad_mask = u_pack_io_img2cvt_dat_wr_pad_mask; // @[NV_NVDLA_CDMA_img.scala 227:32:@10825.4]
  assign io_img2cvt_dat_wr_info_pd = u_pack_io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_CDMA_img.scala 228:31:@10826.4]
  assign io_img2status_state = u_ctrl_io_img2status_state; // @[NV_NVDLA_CDMA_img.scala 114:25:@10710.4]
  assign io_img2status_dat_updt_valid = u_pack_io_img2status_dat_updt_valid; // @[NV_NVDLA_CDMA_img.scala 230:28:@10829.4]
  assign io_img2status_dat_updt_bits_entries = u_pack_io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_img.scala 230:28:@10828.4]
  assign io_img2status_dat_updt_bits_slices = u_pack_io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_CDMA_img.scala 230:28:@10827.4]
  assign io_img2sbuf_p0_wr_addr_valid = u_sg_io_img2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_CDMA_img.scala 172:23:@10773.4]
  assign io_img2sbuf_p0_wr_addr_bits = u_sg_io_img2sbuf_p0_wr_addr_bits[7:0]; // @[NV_NVDLA_CDMA_img.scala 172:23:@10772.4]
  assign io_img2sbuf_p0_wr_data = u_sg_io_img2sbuf_p0_wr_data; // @[NV_NVDLA_CDMA_img.scala 172:23:@10771.4]
  assign io_img2sbuf_p0_rd_addr_valid = u_pack_io_img2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_CDMA_img.scala 194:23:@10794.4]
  assign io_img2sbuf_p0_rd_addr_bits = u_pack_io_img2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_CDMA_img.scala 194:23:@10793.4]
  assign io_dp2reg_img_rd_stall = u_sg_io_dp2reg_img_rd_stall; // @[NV_NVDLA_CDMA_img.scala 187:28:@10786.4]
  assign io_dp2reg_img_rd_latency = u_sg_io_dp2reg_img_rd_latency; // @[NV_NVDLA_CDMA_img.scala 188:30:@10787.4]
  assign u_ctrl_reset = reset; // @[:@10705.4]
  assign u_ctrl_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 108:30:@10706.4]
  assign u_ctrl_io_nvdla_core_ng_clk = io_nvdla_core_ng_clk; // @[NV_NVDLA_CDMA_img.scala 109:33:@10707.4]
  assign u_ctrl_io_pack_is_done = u_pack_io_pack_is_done; // @[NV_NVDLA_CDMA_img.scala 231:28:@10830.4]
  assign u_ctrl_io_sc2cdma_dat_pending_req = io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CDMA_img.scala 111:39:@10708.4]
  assign u_ctrl_io_sg_is_done = u_sg_io_sg_is_done; // @[NV_NVDLA_CDMA_img.scala 147:26:@10746.4]
  assign u_ctrl_io_reg2dp_op_en = io_reg2dp_op_en; // @[NV_NVDLA_CDMA_img.scala 118:28:@10713.4]
  assign u_ctrl_io_reg2dp_conv_mode = io_reg2dp_conv_mode; // @[NV_NVDLA_CDMA_img.scala 119:32:@10714.4]
  assign u_ctrl_io_reg2dp_datain_format = io_reg2dp_datain_format; // @[NV_NVDLA_CDMA_img.scala 122:36:@10717.4]
  assign u_ctrl_io_reg2dp_pixel_format = io_reg2dp_pixel_format; // @[NV_NVDLA_CDMA_img.scala 123:35:@10718.4]
  assign u_ctrl_io_reg2dp_pixel_sign_override = io_reg2dp_pixel_sign_override; // @[NV_NVDLA_CDMA_img.scala 125:42:@10720.4]
  assign u_ctrl_io_reg2dp_datain_width = io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_img.scala 126:35:@10721.4]
  assign u_ctrl_io_reg2dp_data_reuse = io_reg2dp_data_reuse; // @[NV_NVDLA_CDMA_img.scala 127:33:@10722.4]
  assign u_ctrl_io_reg2dp_skip_data_rls = io_reg2dp_skip_data_rls; // @[NV_NVDLA_CDMA_img.scala 128:36:@10723.4]
  assign u_ctrl_io_reg2dp_data_bank = io_reg2dp_data_bank; // @[NV_NVDLA_CDMA_img.scala 129:32:@10724.4]
  assign u_ctrl_io_reg2dp_pixel_x_offset = io_reg2dp_pixel_x_offset; // @[NV_NVDLA_CDMA_img.scala 130:37:@10725.4]
  assign u_ctrl_io_reg2dp_pad_left = io_reg2dp_pad_left; // @[NV_NVDLA_CDMA_img.scala 131:31:@10726.4]
  assign u_ctrl_io_reg2dp_pad_right = io_reg2dp_pad_right; // @[NV_NVDLA_CDMA_img.scala 132:32:@10727.4]
  assign u_sg_reset = reset; // @[:@10730.4]
  assign u_sg_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 136:28:@10731.4]
  assign u_sg_io_img_dat2mcif_rd_req_pd_ready = io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_img.scala 141:31:@10740.4]
  assign u_sg_io_mcif2img_dat_rd_rsp_pd_valid = io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_img.scala 142:36:@10742.4]
  assign u_sg_io_mcif2img_dat_rd_rsp_pd_bits = io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_img.scala 142:36:@10741.4]
  assign u_sg_io_img_dat2cvif_rd_req_pd_ready = io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_img.scala 138:39:@10734.4]
  assign u_sg_io_cvif2img_dat_rd_rsp_pd_valid = io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_img.scala 139:44:@10736.4]
  assign u_sg_io_cvif2img_dat_rd_rsp_pd_bits = io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_img.scala 139:44:@10735.4]
  assign u_sg_io_img2status_dat_entries = io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_img.scala 144:36:@10744.4]
  assign u_sg_io_img2status_dat_updt = io_img2status_dat_updt_valid; // @[NV_NVDLA_CDMA_img.scala 145:33:@10745.4]
  assign u_sg_io_status2dma_free_entries = io_status2dma_free_entries; // @[NV_NVDLA_CDMA_img.scala 170:37:@10769.4]
  assign u_sg_io_status2dma_fsm_switch = io_status2dma_fsm_switch; // @[NV_NVDLA_CDMA_img.scala 171:35:@10770.4]
  assign u_sg_io_is_running = u_ctrl_io_is_running; // @[NV_NVDLA_CDMA_img.scala 148:24:@10747.4]
  assign u_sg_io_layer_st = u_ctrl_io_layer_st; // @[NV_NVDLA_CDMA_img.scala 149:22:@10748.4]
  assign u_sg_io_pixel_order = u_ctrl_io_pixel_order; // @[NV_NVDLA_CDMA_img.scala 150:25:@10749.4]
  assign u_sg_io_pixel_planar = u_ctrl_io_pixel_planar; // @[NV_NVDLA_CDMA_img.scala 151:26:@10750.4]
  assign u_sg_io_pixel_planar0_bundle_limit = u_ctrl_io_pixel_planar0_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 152:40:@10751.4]
  assign u_sg_io_pixel_planar0_bundle_limit_1st = u_ctrl_io_pixel_planar0_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 153:44:@10752.4]
  assign u_sg_io_pixel_planar0_byte_sft = u_ctrl_io_pixel_planar0_byte_sft; // @[NV_NVDLA_CDMA_img.scala 154:36:@10753.4]
  assign u_sg_io_pixel_planar1_byte_sft = u_ctrl_io_pixel_planar1_byte_sft; // @[NV_NVDLA_CDMA_img.scala 155:36:@10754.4]
  assign u_sg_io_pixel_planar0_lp_burst = u_ctrl_io_pixel_planar0_lp_burst; // @[NV_NVDLA_CDMA_img.scala 156:36:@10755.4]
  assign u_sg_io_pixel_planar0_lp_vld = u_ctrl_io_pixel_planar0_lp_vld; // @[NV_NVDLA_CDMA_img.scala 157:34:@10756.4]
  assign u_sg_io_pixel_planar0_rp_burst = u_ctrl_io_pixel_planar0_rp_burst; // @[NV_NVDLA_CDMA_img.scala 158:36:@10757.4]
  assign u_sg_io_pixel_planar0_rp_vld = u_ctrl_io_pixel_planar0_rp_vld; // @[NV_NVDLA_CDMA_img.scala 159:34:@10758.4]
  assign u_sg_io_pixel_planar0_width_burst = u_ctrl_io_pixel_planar0_width_burst; // @[NV_NVDLA_CDMA_img.scala 160:39:@10759.4]
  assign u_sg_io_pixel_planar1_bundle_limit = u_ctrl_io_pixel_planar1_bundle_limit; // @[NV_NVDLA_CDMA_img.scala 161:40:@10760.4]
  assign u_sg_io_pixel_planar1_bundle_limit_1st = u_ctrl_io_pixel_planar1_bundle_limit_1st; // @[NV_NVDLA_CDMA_img.scala 162:44:@10761.4]
  assign u_sg_io_pixel_planar1_lp_burst = u_ctrl_io_pixel_planar1_lp_burst; // @[NV_NVDLA_CDMA_img.scala 163:36:@10762.4]
  assign u_sg_io_pixel_planar1_lp_vld = u_ctrl_io_pixel_planar1_lp_vld; // @[NV_NVDLA_CDMA_img.scala 164:34:@10763.4]
  assign u_sg_io_pixel_planar1_rp_burst = u_ctrl_io_pixel_planar1_rp_burst; // @[NV_NVDLA_CDMA_img.scala 165:36:@10764.4]
  assign u_sg_io_pixel_planar1_rp_vld = u_ctrl_io_pixel_planar1_rp_vld; // @[NV_NVDLA_CDMA_img.scala 166:34:@10765.4]
  assign u_sg_io_pixel_planar1_width_burst = u_ctrl_io_pixel_planar1_width_burst; // @[NV_NVDLA_CDMA_img.scala 167:39:@10766.4]
  assign u_sg_io_sg2pack_img_pd_ready = u_pack_io_sg2pack_img_pd_ready; // @[NV_NVDLA_CDMA_img.scala 215:30:@10814.4]
  assign u_sg_io_reg2dp_op_en = io_reg2dp_op_en; // @[NV_NVDLA_CDMA_img.scala 169:26:@10768.4]
  assign u_sg_io_reg2dp_datain_height = io_reg2dp_datain_height; // @[NV_NVDLA_CDMA_img.scala 175:34:@10775.4]
  assign u_sg_io_reg2dp_datain_ram_type = io_reg2dp_datain_ram_type; // @[NV_NVDLA_CDMA_img.scala 176:36:@10776.4]
  assign u_sg_io_reg2dp_datain_addr_high_0 = io_reg2dp_datain_addr_high_0; // @[NV_NVDLA_CDMA_img.scala 177:39:@10777.4]
  assign u_sg_io_reg2dp_datain_addr_low_0 = io_reg2dp_datain_addr_low_0; // @[NV_NVDLA_CDMA_img.scala 178:38:@10778.4]
  assign u_sg_io_reg2dp_datain_addr_high_1 = io_reg2dp_datain_addr_high_1; // @[NV_NVDLA_CDMA_img.scala 179:39:@10779.4]
  assign u_sg_io_reg2dp_datain_addr_low_1 = io_reg2dp_datain_addr_low_1; // @[NV_NVDLA_CDMA_img.scala 180:38:@10780.4]
  assign u_sg_io_reg2dp_line_stride = io_reg2dp_line_stride; // @[NV_NVDLA_CDMA_img.scala 181:32:@10781.4]
  assign u_sg_io_reg2dp_uv_line_stride = io_reg2dp_uv_line_stride; // @[NV_NVDLA_CDMA_img.scala 182:35:@10782.4]
  assign u_sg_io_reg2dp_mean_format = io_reg2dp_mean_format; // @[NV_NVDLA_CDMA_img.scala 183:32:@10783.4]
  assign u_sg_io_reg2dp_entries = io_reg2dp_entries; // @[NV_NVDLA_CDMA_img.scala 184:28:@10784.4]
  assign u_sg_io_reg2dp_dma_en = io_reg2dp_dma_en; // @[NV_NVDLA_CDMA_img.scala 185:27:@10785.4]
  assign u_pack_reset = reset; // @[:@10790.4]
  assign u_pack_io_nvdla_core_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_img.scala 192:30:@10791.4]
  assign u_pack_io_img2sbuf_p0_rd_data = io_img2sbuf_p0_rd_data; // @[NV_NVDLA_CDMA_img.scala 194:23:@10792.4]
  assign u_pack_io_is_running = u_ctrl_io_is_running; // @[NV_NVDLA_CDMA_img.scala 196:26:@10795.4]
  assign u_pack_io_layer_st = u_ctrl_io_layer_st; // @[NV_NVDLA_CDMA_img.scala 197:24:@10796.4]
  assign u_pack_io_pixel_bank = u_ctrl_io_pixel_bank; // @[NV_NVDLA_CDMA_img.scala 199:26:@10797.4]
  assign u_pack_io_pixel_early_end = u_ctrl_io_pixel_early_end; // @[NV_NVDLA_CDMA_img.scala 202:31:@10800.4]
  assign u_pack_io_pixel_packed_10b = u_ctrl_io_pixel_packed_10b; // @[NV_NVDLA_CDMA_img.scala 203:32:@10801.4]
  assign u_pack_io_pixel_planar = u_ctrl_io_pixel_planar; // @[NV_NVDLA_CDMA_img.scala 204:28:@10802.4]
  assign u_pack_io_pixel_planar0_sft = u_ctrl_io_pixel_planar0_sft; // @[NV_NVDLA_CDMA_img.scala 205:33:@10803.4]
  assign u_pack_io_pixel_planar1_sft = u_ctrl_io_pixel_planar1_sft; // @[NV_NVDLA_CDMA_img.scala 206:33:@10804.4]
  assign u_pack_io_pixel_precision = u_ctrl_io_pixel_precision; // @[NV_NVDLA_CDMA_img.scala 207:31:@10805.4]
  assign u_pack_io_pixel_uint = u_ctrl_io_pixel_uint; // @[NV_NVDLA_CDMA_img.scala 208:26:@10806.4]
  assign u_pack_io_sg2pack_img_pd_valid = u_sg_io_sg2pack_img_pd_valid; // @[NV_NVDLA_CDMA_img.scala 215:30:@10813.4]
  assign u_pack_io_sg2pack_img_pd_bits = u_sg_io_sg2pack_img_pd_bits; // @[NV_NVDLA_CDMA_img.scala 215:30:@10812.4]
  assign u_pack_io_sg2pack_data_entries = u_sg_io_sg2pack_data_entries; // @[NV_NVDLA_CDMA_img.scala 210:36:@10807.4]
  assign u_pack_io_sg2pack_entry_end = u_sg_io_sg2pack_entry_end; // @[NV_NVDLA_CDMA_img.scala 211:33:@10808.4]
  assign u_pack_io_sg2pack_entry_mid = u_sg_io_sg2pack_entry_mid; // @[NV_NVDLA_CDMA_img.scala 212:33:@10809.4]
  assign u_pack_io_sg2pack_entry_st = u_sg_io_sg2pack_entry_st; // @[NV_NVDLA_CDMA_img.scala 213:32:@10810.4]
  assign u_pack_io_sg2pack_height_total = u_sg_io_sg2pack_height_total; // @[NV_NVDLA_CDMA_img.scala 214:36:@10811.4]
  assign u_pack_io_sg2pack_mn_enable = u_sg_io_sg2pack_mn_enable; // @[NV_NVDLA_CDMA_img.scala 216:33:@10815.4]
  assign u_pack_io_sg2pack_sub_h_end = u_sg_io_sg2pack_sub_h_end; // @[NV_NVDLA_CDMA_img.scala 217:33:@10816.4]
  assign u_pack_io_sg2pack_sub_h_mid = u_sg_io_sg2pack_sub_h_mid; // @[NV_NVDLA_CDMA_img.scala 218:33:@10817.4]
  assign u_pack_io_sg2pack_sub_h_st = u_sg_io_sg2pack_sub_h_st; // @[NV_NVDLA_CDMA_img.scala 219:32:@10818.4]
  assign u_pack_io_status2dma_wr_idx = io_status2dma_wr_idx; // @[NV_NVDLA_CDMA_img.scala 220:33:@10819.4]
  assign u_pack_io_reg2dp_datain_width = io_reg2dp_datain_width; // @[NV_NVDLA_CDMA_img.scala 233:35:@10831.4]
  assign u_pack_io_reg2dp_datain_channel = io_reg2dp_datain_channel; // @[NV_NVDLA_CDMA_img.scala 234:37:@10832.4]
  assign u_pack_io_reg2dp_mean_ry = io_reg2dp_mean_ry; // @[NV_NVDLA_CDMA_img.scala 235:30:@10833.4]
  assign u_pack_io_reg2dp_mean_gu = io_reg2dp_mean_gu; // @[NV_NVDLA_CDMA_img.scala 236:30:@10834.4]
  assign u_pack_io_reg2dp_mean_bv = io_reg2dp_mean_bv; // @[NV_NVDLA_CDMA_img.scala 237:30:@10835.4]
  assign u_pack_io_reg2dp_mean_ax = io_reg2dp_mean_ax; // @[NV_NVDLA_CDMA_img.scala 238:30:@10836.4]
  assign u_pack_io_reg2dp_pad_left = io_reg2dp_pad_left; // @[NV_NVDLA_CDMA_img.scala 239:31:@10837.4]
  assign u_pack_io_reg2dp_pad_right = io_reg2dp_pad_right; // @[NV_NVDLA_CDMA_img.scala 240:32:@10838.4]
endmodule
module NV_NVDLA_CDMA_dma_mux( // @[:@11035.2]
  input          reset, // @[:@11037.4]
  input          io_nvdla_core_clk, // @[:@11038.4]
  output         io_dc_dat2mcif_rd_req_pd_ready, // @[:@11038.4]
  input          io_dc_dat2mcif_rd_req_pd_valid, // @[:@11038.4]
  input  [78:0]  io_dc_dat2mcif_rd_req_pd_bits, // @[:@11038.4]
  input          io_mcif2dc_dat_rd_rsp_pd_ready, // @[:@11038.4]
  output         io_mcif2dc_dat_rd_rsp_pd_valid, // @[:@11038.4]
  output [256:0] io_mcif2dc_dat_rd_rsp_pd_bits, // @[:@11038.4]
  output         io_img_dat2mcif_rd_req_pd_ready, // @[:@11038.4]
  input          io_img_dat2mcif_rd_req_pd_valid, // @[:@11038.4]
  input  [78:0]  io_img_dat2mcif_rd_req_pd_bits, // @[:@11038.4]
  input          io_mcif2img_dat_rd_rsp_pd_ready, // @[:@11038.4]
  output         io_mcif2img_dat_rd_rsp_pd_valid, // @[:@11038.4]
  output [256:0] io_mcif2img_dat_rd_rsp_pd_bits, // @[:@11038.4]
  input          io_cdma_dat2mcif_rd_req_pd_ready, // @[:@11038.4]
  output         io_cdma_dat2mcif_rd_req_pd_valid, // @[:@11038.4]
  output [78:0]  io_cdma_dat2mcif_rd_req_pd_bits, // @[:@11038.4]
  output         io_mcif2cdma_dat_rd_rsp_pd_ready, // @[:@11038.4]
  input          io_mcif2cdma_dat_rd_rsp_pd_valid, // @[:@11038.4]
  input  [256:0] io_mcif2cdma_dat_rd_rsp_pd_bits, // @[:@11038.4]
  output         io_dc_dat2cvif_rd_req_pd_ready, // @[:@11038.4]
  input          io_dc_dat2cvif_rd_req_pd_valid, // @[:@11038.4]
  input  [78:0]  io_dc_dat2cvif_rd_req_pd_bits, // @[:@11038.4]
  input          io_cvif2dc_dat_rd_rsp_pd_ready, // @[:@11038.4]
  output         io_cvif2dc_dat_rd_rsp_pd_valid, // @[:@11038.4]
  output [256:0] io_cvif2dc_dat_rd_rsp_pd_bits, // @[:@11038.4]
  output         io_img_dat2cvif_rd_req_pd_ready, // @[:@11038.4]
  input          io_img_dat2cvif_rd_req_pd_valid, // @[:@11038.4]
  input  [78:0]  io_img_dat2cvif_rd_req_pd_bits, // @[:@11038.4]
  input          io_cvif2img_dat_rd_rsp_pd_ready, // @[:@11038.4]
  output         io_cvif2img_dat_rd_rsp_pd_valid, // @[:@11038.4]
  output [256:0] io_cvif2img_dat_rd_rsp_pd_bits, // @[:@11038.4]
  input          io_cdma_dat2cvif_rd_req_pd_ready, // @[:@11038.4]
  output         io_cdma_dat2cvif_rd_req_pd_valid, // @[:@11038.4]
  output [78:0]  io_cdma_dat2cvif_rd_req_pd_bits, // @[:@11038.4]
  output         io_cvif2cdma_dat_rd_rsp_pd_ready, // @[:@11038.4]
  input          io_cvif2cdma_dat_rd_rsp_pd_valid, // @[:@11038.4]
  input  [256:0] io_cvif2cdma_dat_rd_rsp_pd_bits // @[:@11038.4]
);
  wire  NV_NVDLA_IS_pipe_reset; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_io_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire [78:0] NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_io_ri; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire [78:0] NV_NVDLA_IS_pipe_io_di; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_io_vi; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
  wire  NV_NVDLA_IS_pipe_1_reset; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_1_io_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire [256:0] NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_1_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_1_io_ri; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire [256:0] NV_NVDLA_IS_pipe_1_io_di; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_1_io_vi; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_1_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
  wire  NV_NVDLA_IS_pipe_2_reset; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_2_io_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire [78:0] NV_NVDLA_IS_pipe_2_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_2_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_2_io_ri; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire [78:0] NV_NVDLA_IS_pipe_2_io_di; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_2_io_vi; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_2_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
  wire  NV_NVDLA_IS_pipe_3_reset; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  NV_NVDLA_IS_pipe_3_io_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire [78:0] NV_NVDLA_IS_pipe_3_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  NV_NVDLA_IS_pipe_3_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  NV_NVDLA_IS_pipe_3_io_ri; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire [78:0] NV_NVDLA_IS_pipe_3_io_di; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  NV_NVDLA_IS_pipe_3_io_vi; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  NV_NVDLA_IS_pipe_3_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
  wire  _T_115; // @[NV_NVDLA_CDMA_dma_mux.scala 69:56:@11040.4]
  wire [78:0] _T_119; // @[Bitwise.scala 72:12:@11042.4]
  wire [78:0] _T_120; // @[NV_NVDLA_CDMA_dma_mux.scala 70:70:@11043.4]
  wire [78:0] _T_124; // @[Bitwise.scala 72:12:@11045.4]
  wire [78:0] _T_125; // @[NV_NVDLA_CDMA_dma_mux.scala 71:71:@11046.4]
  wire  _T_132; // @[NV_NVDLA_CDMA_dma_mux.scala 89:68:@11063.4]
  reg  _T_134; // @[Reg.scala 19:20:@11064.4]
  reg [31:0] _RAND_0;
  wire  _GEN_0; // @[Reg.scala 20:19:@11065.4]
  reg  _T_138; // @[Reg.scala 19:20:@11069.4]
  reg [31:0] _RAND_1;
  wire  _GEN_1; // @[Reg.scala 20:19:@11070.4]
  wire [256:0] _T_146; // @[Bitwise.scala 72:12:@11087.4]
  wire [256:0] _T_151; // @[Bitwise.scala 72:12:@11091.4]
  wire  _T_153; // @[NV_NVDLA_CDMA_dma_mux.scala 114:35:@11094.4]
  wire  _T_154; // @[NV_NVDLA_CDMA_dma_mux.scala 114:81:@11095.4]
  wire  _T_156; // @[NV_NVDLA_CDMA_dma_mux.scala 125:60:@11098.4]
  wire [78:0] _T_160; // @[Bitwise.scala 72:12:@11100.4]
  wire [78:0] _T_161; // @[NV_NVDLA_CDMA_dma_mux.scala 126:70:@11101.4]
  wire [78:0] _T_165; // @[Bitwise.scala 72:12:@11103.4]
  wire [78:0] _T_166; // @[NV_NVDLA_CDMA_dma_mux.scala 127:71:@11104.4]
  wire  _T_173; // @[NV_NVDLA_CDMA_dma_mux.scala 145:68:@11121.4]
  reg  _T_175; // @[Reg.scala 19:20:@11122.4]
  reg [31:0] _RAND_2;
  wire  _GEN_2; // @[Reg.scala 20:19:@11123.4]
  reg  _T_179; // @[Reg.scala 19:20:@11127.4]
  reg [31:0] _RAND_3;
  wire  _GEN_3; // @[Reg.scala 20:19:@11128.4]
  wire [256:0] _T_187; // @[Bitwise.scala 72:12:@11145.4]
  wire [256:0] _GEN_4; // @[NV_NVDLA_CDMA_dma_mux.scala 167:86:@11146.4]
  wire [256:0] _T_192; // @[Bitwise.scala 72:12:@11149.4]
  wire  _T_194; // @[NV_NVDLA_CDMA_dma_mux.scala 169:35:@11152.4]
  wire  _T_195; // @[NV_NVDLA_CDMA_dma_mux.scala 169:85:@11153.4]
  NV_NVDLA_IS_pipe NV_NVDLA_IS_pipe ( // @[NV_NVDLA_CDMA_dma_mux.scala 74:25:@11049.4]
    .reset(NV_NVDLA_IS_pipe_reset),
    .io_clk(NV_NVDLA_IS_pipe_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_io_ri),
    .io_di(NV_NVDLA_IS_pipe_io_di),
    .io_vi(NV_NVDLA_IS_pipe_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_io_ro)
  );
  NV_NVDLA_IS_pipe_2 NV_NVDLA_IS_pipe_1 ( // @[NV_NVDLA_CDMA_dma_mux.scala 100:25:@11074.4]
    .reset(NV_NVDLA_IS_pipe_1_reset),
    .io_clk(NV_NVDLA_IS_pipe_1_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_1_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_1_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_1_io_ri),
    .io_di(NV_NVDLA_IS_pipe_1_io_di),
    .io_vi(NV_NVDLA_IS_pipe_1_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_1_io_ro)
  );
  NV_NVDLA_IS_pipe NV_NVDLA_IS_pipe_2 ( // @[NV_NVDLA_CDMA_dma_mux.scala 130:25:@11107.4]
    .reset(NV_NVDLA_IS_pipe_2_reset),
    .io_clk(NV_NVDLA_IS_pipe_2_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_2_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_2_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_2_io_ri),
    .io_di(NV_NVDLA_IS_pipe_2_io_di),
    .io_vi(NV_NVDLA_IS_pipe_2_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_2_io_ro)
  );
  NV_NVDLA_IS_pipe NV_NVDLA_IS_pipe_3 ( // @[NV_NVDLA_CDMA_dma_mux.scala 155:25:@11132.4]
    .reset(NV_NVDLA_IS_pipe_3_reset),
    .io_clk(NV_NVDLA_IS_pipe_3_io_clk),
    .io_dout(NV_NVDLA_IS_pipe_3_io_dout),
    .io_vo(NV_NVDLA_IS_pipe_3_io_vo),
    .io_ri(NV_NVDLA_IS_pipe_3_io_ri),
    .io_di(NV_NVDLA_IS_pipe_3_io_di),
    .io_vi(NV_NVDLA_IS_pipe_3_io_vi),
    .io_ro(NV_NVDLA_IS_pipe_3_io_ro)
  );
  assign _T_115 = io_dc_dat2mcif_rd_req_pd_valid | io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 69:56:@11040.4]
  assign _T_119 = io_dc_dat2mcif_rd_req_pd_valid ? 79'h7fffffffffffffffffff : 79'h0; // @[Bitwise.scala 72:12:@11042.4]
  assign _T_120 = _T_119 & io_dc_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dma_mux.scala 70:70:@11043.4]
  assign _T_124 = io_img_dat2mcif_rd_req_pd_valid ? 79'h7fffffffffffffffffff : 79'h0; // @[Bitwise.scala 72:12:@11045.4]
  assign _T_125 = _T_124 & io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dma_mux.scala 71:71:@11046.4]
  assign _T_132 = _T_115 & NV_NVDLA_IS_pipe_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 89:68:@11063.4]
  assign _GEN_0 = _T_132 ? io_dc_dat2mcif_rd_req_pd_valid : _T_134; // @[Reg.scala 20:19:@11065.4]
  assign _GEN_1 = _T_132 ? io_img_dat2mcif_rd_req_pd_valid : _T_138; // @[Reg.scala 20:19:@11070.4]
  assign _T_146 = _T_134 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@11087.4]
  assign _T_151 = _T_138 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@11091.4]
  assign _T_153 = _T_134 & io_mcif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 114:35:@11094.4]
  assign _T_154 = _T_138 & io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 114:81:@11095.4]
  assign _T_156 = io_dc_dat2cvif_rd_req_pd_valid | io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 125:60:@11098.4]
  assign _T_160 = io_dc_dat2cvif_rd_req_pd_valid ? 79'h7fffffffffffffffffff : 79'h0; // @[Bitwise.scala 72:12:@11100.4]
  assign _T_161 = _T_160 & io_dc_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dma_mux.scala 126:70:@11101.4]
  assign _T_165 = io_img_dat2cvif_rd_req_pd_valid ? 79'h7fffffffffffffffffff : 79'h0; // @[Bitwise.scala 72:12:@11103.4]
  assign _T_166 = _T_165 & io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_CDMA_dma_mux.scala 127:71:@11104.4]
  assign _T_173 = _T_156 & NV_NVDLA_IS_pipe_2_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 145:68:@11121.4]
  assign _GEN_2 = _T_173 ? io_dc_dat2cvif_rd_req_pd_valid : _T_175; // @[Reg.scala 20:19:@11123.4]
  assign _GEN_3 = _T_173 ? io_img_dat2cvif_rd_req_pd_valid : _T_179; // @[Reg.scala 20:19:@11128.4]
  assign _T_187 = _T_175 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@11145.4]
  assign _GEN_4 = {{178'd0}, NV_NVDLA_IS_pipe_3_io_dout}; // @[NV_NVDLA_CDMA_dma_mux.scala 167:86:@11146.4]
  assign _T_192 = _T_179 ? 257'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 257'h0; // @[Bitwise.scala 72:12:@11149.4]
  assign _T_194 = _T_175 & io_cvif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 169:35:@11152.4]
  assign _T_195 = _T_179 & io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 169:85:@11153.4]
  assign io_dc_dat2mcif_rd_req_pd_ready = NV_NVDLA_IS_pipe_io_ro & io_dc_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 83:36:@11057.4]
  assign io_mcif2dc_dat_rd_rsp_pd_valid = NV_NVDLA_IS_pipe_1_io_vo & _T_134; // @[NV_NVDLA_CDMA_dma_mux.scala 110:37:@11083.4]
  assign io_mcif2dc_dat_rd_rsp_pd_bits = _T_146 & NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 112:35:@11089.4]
  assign io_img_dat2mcif_rd_req_pd_ready = NV_NVDLA_IS_pipe_io_ro & io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 84:37:@11059.4]
  assign io_mcif2img_dat_rd_rsp_pd_valid = NV_NVDLA_IS_pipe_1_io_vo & _T_138; // @[NV_NVDLA_CDMA_dma_mux.scala 111:37:@11085.4]
  assign io_mcif2img_dat_rd_rsp_pd_bits = _T_151 & NV_NVDLA_IS_pipe_1_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 113:36:@11093.4]
  assign io_cdma_dat2mcif_rd_req_pd_valid = NV_NVDLA_IS_pipe_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 85:38:@11060.4]
  assign io_cdma_dat2mcif_rd_req_pd_bits = NV_NVDLA_IS_pipe_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 86:37:@11061.4]
  assign io_mcif2cdma_dat_rd_rsp_pd_ready = NV_NVDLA_IS_pipe_1_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 109:38:@11081.4]
  assign io_dc_dat2cvif_rd_req_pd_ready = NV_NVDLA_IS_pipe_2_io_ro & io_dc_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 139:40:@11115.4]
  assign io_cvif2dc_dat_rd_rsp_pd_valid = NV_NVDLA_IS_pipe_3_io_vo & _T_175; // @[NV_NVDLA_CDMA_dma_mux.scala 165:40:@11141.4]
  assign io_cvif2dc_dat_rd_rsp_pd_bits = _T_187 & _GEN_4; // @[NV_NVDLA_CDMA_dma_mux.scala 167:39:@11147.4]
  assign io_img_dat2cvif_rd_req_pd_ready = NV_NVDLA_IS_pipe_2_io_ro & io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 140:41:@11117.4]
  assign io_cvif2img_dat_rd_rsp_pd_valid = NV_NVDLA_IS_pipe_3_io_vo & _T_179; // @[NV_NVDLA_CDMA_dma_mux.scala 166:41:@11143.4]
  assign io_cvif2img_dat_rd_rsp_pd_bits = _T_192 & _GEN_4; // @[NV_NVDLA_CDMA_dma_mux.scala 168:40:@11151.4]
  assign io_cdma_dat2cvif_rd_req_pd_valid = NV_NVDLA_IS_pipe_2_io_vo; // @[NV_NVDLA_CDMA_dma_mux.scala 141:42:@11118.4]
  assign io_cdma_dat2cvif_rd_req_pd_bits = NV_NVDLA_IS_pipe_2_io_dout; // @[NV_NVDLA_CDMA_dma_mux.scala 142:41:@11119.4]
  assign io_cvif2cdma_dat_rd_rsp_pd_ready = NV_NVDLA_IS_pipe_3_io_ro; // @[NV_NVDLA_CDMA_dma_mux.scala 164:42:@11139.4]
  assign NV_NVDLA_IS_pipe_reset = reset; // @[:@11051.4]
  assign NV_NVDLA_IS_pipe_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 75:20:@11052.4]
  assign NV_NVDLA_IS_pipe_io_ri = io_cdma_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 80:19:@11055.4]
  assign NV_NVDLA_IS_pipe_io_di = _T_120 | _T_125; // @[NV_NVDLA_CDMA_dma_mux.scala 78:19:@11054.4]
  assign NV_NVDLA_IS_pipe_io_vi = io_dc_dat2mcif_rd_req_pd_valid | io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 76:19:@11053.4]
  assign NV_NVDLA_IS_pipe_1_reset = reset; // @[:@11076.4]
  assign NV_NVDLA_IS_pipe_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 101:20:@11077.4]
  assign NV_NVDLA_IS_pipe_1_io_ri = _T_153 | _T_154; // @[NV_NVDLA_CDMA_dma_mux.scala 106:19:@11080.4]
  assign NV_NVDLA_IS_pipe_1_io_di = io_mcif2cdma_dat_rd_rsp_pd_bits; // @[NV_NVDLA_CDMA_dma_mux.scala 104:19:@11079.4]
  assign NV_NVDLA_IS_pipe_1_io_vi = io_mcif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 102:19:@11078.4]
  assign NV_NVDLA_IS_pipe_2_reset = reset; // @[:@11109.4]
  assign NV_NVDLA_IS_pipe_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 131:20:@11110.4]
  assign NV_NVDLA_IS_pipe_2_io_ri = io_cdma_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_CDMA_dma_mux.scala 136:19:@11113.4]
  assign NV_NVDLA_IS_pipe_2_io_di = _T_161 | _T_166; // @[NV_NVDLA_CDMA_dma_mux.scala 134:19:@11112.4]
  assign NV_NVDLA_IS_pipe_2_io_vi = io_dc_dat2cvif_rd_req_pd_valid | io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 132:19:@11111.4]
  assign NV_NVDLA_IS_pipe_3_reset = reset; // @[:@11134.4]
  assign NV_NVDLA_IS_pipe_3_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_dma_mux.scala 156:20:@11135.4]
  assign NV_NVDLA_IS_pipe_3_io_ri = _T_194 | _T_195; // @[NV_NVDLA_CDMA_dma_mux.scala 161:19:@11138.4]
  assign NV_NVDLA_IS_pipe_3_io_di = io_cvif2cdma_dat_rd_rsp_pd_bits[78:0]; // @[NV_NVDLA_CDMA_dma_mux.scala 159:19:@11137.4]
  assign NV_NVDLA_IS_pipe_3_io_vi = io_cvif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_CDMA_dma_mux.scala 157:19:@11136.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_134 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_138 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_175 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_179 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_134 <= 1'h0;
    end else begin
      if (_T_132) begin
        _T_134 <= io_dc_dat2mcif_rd_req_pd_valid;
      end
    end
    if (reset) begin
      _T_138 <= 1'h0;
    end else begin
      if (_T_132) begin
        _T_138 <= io_img_dat2mcif_rd_req_pd_valid;
      end
    end
    if (reset) begin
      _T_175 <= 1'h0;
    end else begin
      if (_T_173) begin
        _T_175 <= io_dc_dat2cvif_rd_req_pd_valid;
      end
    end
    if (reset) begin
      _T_179 <= 1'h0;
    end else begin
      if (_T_173) begin
        _T_179 <= io_img_dat2cvif_rd_req_pd_valid;
      end
    end
  end
endmodule
module NV_NVDLA_BC_pipe( // @[:@11164.2]
  input         reset, // @[:@11166.4]
  input         io_clk, // @[:@11167.4]
  input         io_vi, // @[:@11167.4]
  output        io_ro, // @[:@11167.4]
  input  [17:0] io_di, // @[:@11167.4]
  output        io_vo, // @[:@11167.4]
  input         io_ri, // @[:@11167.4]
  output [17:0] io_dout // @[:@11167.4]
);
  reg  _T_21; // @[BC_pipe.scala 49:29:@11169.4]
  reg [31:0] _RAND_0;
  reg [17:0] _T_23; // @[BC_pipe.scala 50:24:@11170.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[BC_pipe.scala 53:22:@11172.4]
  wire  _T_29; // @[BC_pipe.scala 54:28:@11174.4]
  wire  _T_31; // @[BC_pipe.scala 55:28:@11177.4]
  assign _T_27 = io_ro ? io_vi : 1'h1; // @[BC_pipe.scala 53:22:@11172.4]
  assign _T_29 = _T_21 == 1'h0; // @[BC_pipe.scala 54:28:@11174.4]
  assign _T_31 = io_ro & io_vi; // @[BC_pipe.scala 55:28:@11177.4]
  assign io_ro = io_ri | _T_29; // @[BC_pipe.scala 54:11:@11176.4]
  assign io_vo = _T_21; // @[BC_pipe.scala 59:11:@11181.4]
  assign io_dout = _T_23; // @[BC_pipe.scala 60:13:@11182.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_23 = _RAND_1[17:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      if (io_ro) begin
        _T_21 <= io_vi;
      end else begin
        _T_21 <= 1'h1;
      end
    end
    if (_T_31) begin
      _T_23 <= io_di;
    end
  end
endmodule
module NV_NVDLA_BC_pipe_1( // @[:@11184.2]
  input         reset, // @[:@11186.4]
  input         io_clk, // @[:@11187.4]
  input         io_vi, // @[:@11187.4]
  output        io_ro, // @[:@11187.4]
  input  [33:0] io_di, // @[:@11187.4]
  output        io_vo, // @[:@11187.4]
  input         io_ri, // @[:@11187.4]
  output [33:0] io_dout // @[:@11187.4]
);
  reg  _T_21; // @[BC_pipe.scala 49:29:@11189.4]
  reg [31:0] _RAND_0;
  reg [33:0] _T_23; // @[BC_pipe.scala 50:24:@11190.4]
  reg [63:0] _RAND_1;
  wire  _T_27; // @[BC_pipe.scala 53:22:@11192.4]
  wire  _T_29; // @[BC_pipe.scala 54:28:@11194.4]
  wire  _T_31; // @[BC_pipe.scala 55:28:@11197.4]
  assign _T_27 = io_ro ? io_vi : 1'h1; // @[BC_pipe.scala 53:22:@11192.4]
  assign _T_29 = _T_21 == 1'h0; // @[BC_pipe.scala 54:28:@11194.4]
  assign _T_31 = io_ro & io_vi; // @[BC_pipe.scala 55:28:@11197.4]
  assign io_ro = io_ri | _T_29; // @[BC_pipe.scala 54:11:@11196.4]
  assign io_vo = _T_21; // @[BC_pipe.scala 59:11:@11201.4]
  assign io_dout = _T_23; // @[BC_pipe.scala 60:13:@11202.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_23 = _RAND_1[33:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      if (io_ro) begin
        _T_21 <= io_vi;
      end else begin
        _T_21 <= 1'h1;
      end
    end
    if (_T_31) begin
      _T_23 <= io_di;
    end
  end
endmodule
module NV_soDLA_HLS_shiftrightsu( // @[:@11204.2]
  input  [33:0] io_data_in, // @[:@11207.4]
  input  [5:0]  io_shift_num, // @[:@11207.4]
  output [16:0] io_data_out // @[:@11207.4]
);
  wire  data_sign; // @[NV_NVDLA_HLS_shiftrightsu.scala 25:28:@11218.4]
  wire [33:0] _T_24; // @[Bitwise.scala 72:12:@11221.4]
  wire [101:0] _T_31; // @[Cat.scala 30:58:@11224.4]
  wire [101:0] _T_32; // @[NV_NVDLA_HLS_shiftrightsu.scala 27:87:@11225.4]
  wire [33:0] data_shift; // @[NV_NVDLA_HLS_shiftrightsu.scala 29:104:@11234.4]
  wire  guide; // @[NV_NVDLA_HLS_shiftrightsu.scala 31:99:@11242.4]
  wire [32:0] _T_72; // @[NV_NVDLA_HLS_shiftrightsu.scala 33:99:@11250.4]
  wire  _T_73; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:24:@11252.4]
  wire [33:0] stick; // @[NV_NVDLA_HLS_shiftrightsu.scala 17:21:@11211.4 NV_NVDLA_HLS_shiftrightsu.scala 33:11:@11251.4]
  wire  _T_75; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:43:@11253.4]
  wire  _T_76; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:35:@11254.4]
  wire  point5; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:21:@11255.4]
  wire [16:0] _T_78; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:29:@11257.4]
  wire [16:0] _GEN_0; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11258.4]
  wire [17:0] _T_79; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11258.4]
  wire [16:0] data_round; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11259.4]
  wire [16:0] _T_81; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:49:@11261.4]
  wire [16:0] _T_82; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:75:@11262.4]
  wire  _T_84; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:75:@11263.4]
  wire  _T_85; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:37:@11264.4]
  wire  _T_86; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:35:@11265.4]
  wire  _T_90; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:75:@11268.4]
  wire  _T_91; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:35:@11269.4]
  wire  _T_92; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:82:@11270.4]
  wire [15:0] _T_94; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:52:@11272.4]
  wire [16:0] _T_95; // @[Cat.scala 30:58:@11273.4]
  wire [16:0] _T_96; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:86:@11274.4]
  wire  _T_98; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:86:@11275.4]
  wire  _T_99; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:35:@11276.4]
  wire  tru_need_sat; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:81:@11277.4]
  wire [16:0] data_max; // @[NV_NVDLA_HLS_shiftrightsu.scala 43:20:@11284.4]
  wire  _T_118; // @[NV_NVDLA_HLS_shiftrightsu.scala 45:37:@11286.4]
  wire [16:0] _T_124; // @[NV_NVDLA_HLS_shiftrightsu.scala 45:81:@11288.4]
  assign data_sign = io_data_in[33]; // @[NV_NVDLA_HLS_shiftrightsu.scala 25:28:@11218.4]
  assign _T_24 = data_sign ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@11221.4]
  assign _T_31 = {_T_24,io_data_in,34'h0}; // @[Cat.scala 30:58:@11224.4]
  assign _T_32 = _T_31 >> io_shift_num; // @[NV_NVDLA_HLS_shiftrightsu.scala 27:87:@11225.4]
  assign data_shift = _T_32[67:34]; // @[NV_NVDLA_HLS_shiftrightsu.scala 29:104:@11234.4]
  assign guide = _T_32[33]; // @[NV_NVDLA_HLS_shiftrightsu.scala 31:99:@11242.4]
  assign _T_72 = _T_32[32:0]; // @[NV_NVDLA_HLS_shiftrightsu.scala 33:99:@11250.4]
  assign _T_73 = ~ data_sign; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:24:@11252.4]
  assign stick = {{1'd0}, _T_72}; // @[NV_NVDLA_HLS_shiftrightsu.scala 17:21:@11211.4 NV_NVDLA_HLS_shiftrightsu.scala 33:11:@11251.4]
  assign _T_75 = stick != 34'h0; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:43:@11253.4]
  assign _T_76 = _T_73 | _T_75; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:35:@11254.4]
  assign point5 = guide & _T_76; // @[NV_NVDLA_HLS_shiftrightsu.scala 35:21:@11255.4]
  assign _T_78 = data_shift[16:0]; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:29:@11257.4]
  assign _GEN_0 = {{16'd0}, point5}; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11258.4]
  assign _T_79 = _T_78 + _GEN_0; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11258.4]
  assign data_round = _T_78 + _GEN_0; // @[NV_NVDLA_HLS_shiftrightsu.scala 37:46:@11259.4]
  assign _T_81 = data_shift[32:16]; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:49:@11261.4]
  assign _T_82 = ~ _T_81; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:75:@11262.4]
  assign _T_84 = _T_82 == 17'h0; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:75:@11263.4]
  assign _T_85 = ~ _T_84; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:37:@11264.4]
  assign _T_86 = data_sign & _T_85; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:35:@11265.4]
  assign _T_90 = _T_81 != 17'h0; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:75:@11268.4]
  assign _T_91 = _T_73 & _T_90; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:35:@11269.4]
  assign _T_92 = _T_86 | _T_91; // @[NV_NVDLA_HLS_shiftrightsu.scala 39:82:@11270.4]
  assign _T_94 = data_shift[15:0]; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:52:@11272.4]
  assign _T_95 = {_T_94,point5}; // @[Cat.scala 30:58:@11273.4]
  assign _T_96 = ~ _T_95; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:86:@11274.4]
  assign _T_98 = _T_96 == 17'h0; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:86:@11275.4]
  assign _T_99 = _T_73 & _T_98; // @[NV_NVDLA_HLS_shiftrightsu.scala 41:35:@11276.4]
  assign tru_need_sat = _T_92 | _T_99; // @[NV_NVDLA_HLS_shiftrightsu.scala 40:81:@11277.4]
  assign data_max = data_sign ? 17'h10000 : 17'hffff; // @[NV_NVDLA_HLS_shiftrightsu.scala 43:20:@11284.4]
  assign _T_118 = io_shift_num >= 6'h22; // @[NV_NVDLA_HLS_shiftrightsu.scala 45:37:@11286.4]
  assign _T_124 = tru_need_sat ? data_max : data_round; // @[NV_NVDLA_HLS_shiftrightsu.scala 45:81:@11288.4]
  assign io_data_out = _T_118 ? 17'h0 : _T_124; // @[NV_NVDLA_HLS_shiftrightsu.scala 45:17:@11290.4]
endmodule
module NV_soDLA_HLS_saturate( // @[:@11292.2]
  input  [16:0] io_data_in, // @[:@11295.4]
  output [15:0] io_data_out // @[:@11295.4]
);
  wire  data_sign; // @[NV_NVDLA_HLS_saturate.scala 18:28:@11300.4]
  wire  _T_13; // @[NV_NVDLA_HLS_saturate.scala 20:46:@11302.4]
  wire  _T_14; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11303.4]
  wire  _T_16; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11304.4]
  wire  _T_17; // @[NV_NVDLA_HLS_saturate.scala 20:34:@11305.4]
  wire  _T_18; // @[NV_NVDLA_HLS_saturate.scala 20:32:@11306.4]
  wire  _T_19; // @[NV_NVDLA_HLS_saturate.scala 20:82:@11307.4]
  wire  _T_23; // @[NV_NVDLA_HLS_saturate.scala 20:93:@11310.4]
  wire  tru_need_sat; // @[NV_NVDLA_HLS_saturate.scala 20:79:@11311.4]
  wire [15:0] data_max; // @[NV_NVDLA_HLS_saturate.scala 22:20:@11318.4]
  wire [16:0] _T_41; // @[NV_NVDLA_HLS_saturate.scala 24:23:@11320.4]
  assign data_sign = io_data_in[16]; // @[NV_NVDLA_HLS_saturate.scala 18:28:@11300.4]
  assign _T_13 = io_data_in[15]; // @[NV_NVDLA_HLS_saturate.scala 20:46:@11302.4]
  assign _T_14 = ~ _T_13; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11303.4]
  assign _T_16 = _T_14 == 1'h0; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11304.4]
  assign _T_17 = ~ _T_16; // @[NV_NVDLA_HLS_saturate.scala 20:34:@11305.4]
  assign _T_18 = data_sign & _T_17; // @[NV_NVDLA_HLS_saturate.scala 20:32:@11306.4]
  assign _T_19 = ~ data_sign; // @[NV_NVDLA_HLS_saturate.scala 20:82:@11307.4]
  assign _T_23 = _T_19 & _T_13; // @[NV_NVDLA_HLS_saturate.scala 20:93:@11310.4]
  assign tru_need_sat = _T_18 | _T_23; // @[NV_NVDLA_HLS_saturate.scala 20:79:@11311.4]
  assign data_max = data_sign ? 16'h8000 : 16'h7fff; // @[NV_NVDLA_HLS_saturate.scala 22:20:@11318.4]
  assign _T_41 = tru_need_sat ? {{1'd0}, data_max} : io_data_in; // @[NV_NVDLA_HLS_saturate.scala 24:23:@11320.4]
  assign io_data_out = _T_41[15:0]; // @[NV_NVDLA_HLS_saturate.scala 24:17:@11321.4]
endmodule
module NV_soDLA_HLS_saturate_1( // @[:@11323.2]
  input  [16:0] io_data_in, // @[:@11326.4]
  output [7:0]  io_data_out // @[:@11326.4]
);
  wire  data_sign; // @[NV_NVDLA_HLS_saturate.scala 18:28:@11331.4]
  wire [8:0] _T_13; // @[NV_NVDLA_HLS_saturate.scala 20:46:@11333.4]
  wire [8:0] _T_14; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11334.4]
  wire  _T_16; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11335.4]
  wire  _T_17; // @[NV_NVDLA_HLS_saturate.scala 20:34:@11336.4]
  wire  _T_18; // @[NV_NVDLA_HLS_saturate.scala 20:32:@11337.4]
  wire  _T_19; // @[NV_NVDLA_HLS_saturate.scala 20:82:@11338.4]
  wire  _T_22; // @[NV_NVDLA_HLS_saturate.scala 20:132:@11340.4]
  wire  _T_23; // @[NV_NVDLA_HLS_saturate.scala 20:93:@11341.4]
  wire  tru_need_sat; // @[NV_NVDLA_HLS_saturate.scala 20:79:@11342.4]
  wire [7:0] data_max; // @[NV_NVDLA_HLS_saturate.scala 22:20:@11349.4]
  wire [16:0] _T_41; // @[NV_NVDLA_HLS_saturate.scala 24:23:@11351.4]
  assign data_sign = io_data_in[16]; // @[NV_NVDLA_HLS_saturate.scala 18:28:@11331.4]
  assign _T_13 = io_data_in[15:7]; // @[NV_NVDLA_HLS_saturate.scala 20:46:@11333.4]
  assign _T_14 = ~ _T_13; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11334.4]
  assign _T_16 = _T_14 == 9'h0; // @[NV_NVDLA_HLS_saturate.scala 20:72:@11335.4]
  assign _T_17 = ~ _T_16; // @[NV_NVDLA_HLS_saturate.scala 20:34:@11336.4]
  assign _T_18 = data_sign & _T_17; // @[NV_NVDLA_HLS_saturate.scala 20:32:@11337.4]
  assign _T_19 = ~ data_sign; // @[NV_NVDLA_HLS_saturate.scala 20:82:@11338.4]
  assign _T_22 = _T_13 != 9'h0; // @[NV_NVDLA_HLS_saturate.scala 20:132:@11340.4]
  assign _T_23 = _T_19 & _T_22; // @[NV_NVDLA_HLS_saturate.scala 20:93:@11341.4]
  assign tru_need_sat = _T_18 | _T_23; // @[NV_NVDLA_HLS_saturate.scala 20:79:@11342.4]
  assign data_max = data_sign ? 8'h80 : 8'h7f; // @[NV_NVDLA_HLS_saturate.scala 22:20:@11349.4]
  assign _T_41 = tru_need_sat ? {{9'd0}, data_max} : io_data_in; // @[NV_NVDLA_HLS_saturate.scala 24:23:@11351.4]
  assign io_data_out = _T_41[7:0]; // @[NV_NVDLA_HLS_saturate.scala 24:17:@11352.4]
endmodule
module NV_NVDLA_BC_pipe_2( // @[:@11354.2]
  input         reset, // @[:@11356.4]
  input         io_clk, // @[:@11357.4]
  input         io_vi, // @[:@11357.4]
  output        io_ro, // @[:@11357.4]
  input  [15:0] io_di, // @[:@11357.4]
  input         io_ri, // @[:@11357.4]
  output [15:0] io_dout // @[:@11357.4]
);
  reg  _T_21; // @[BC_pipe.scala 49:29:@11359.4]
  reg [31:0] _RAND_0;
  reg [15:0] _T_23; // @[BC_pipe.scala 50:24:@11360.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[BC_pipe.scala 53:22:@11362.4]
  wire  _T_29; // @[BC_pipe.scala 54:28:@11364.4]
  wire  _T_31; // @[BC_pipe.scala 55:28:@11367.4]
  assign _T_27 = io_ro ? io_vi : 1'h1; // @[BC_pipe.scala 53:22:@11362.4]
  assign _T_29 = _T_21 == 1'h0; // @[BC_pipe.scala 54:28:@11364.4]
  assign _T_31 = io_ro & io_vi; // @[BC_pipe.scala 55:28:@11367.4]
  assign io_ro = io_ri | _T_29; // @[BC_pipe.scala 54:11:@11366.4]
  assign io_dout = _T_23; // @[BC_pipe.scala 60:13:@11372.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_21 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_23 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      if (io_ro) begin
        _T_21 <= io_vi;
      end else begin
        _T_21 <= 1'h1;
      end
    end
    if (_T_31) begin
      _T_23 <= io_di;
    end
  end
endmodule
module NV_NVDLA_CDMA_CVT_cell( // @[:@11374.2]
  input         reset, // @[:@11376.4]
  input         io_nvdla_core_clk, // @[:@11377.4]
  input  [15:0] io_cfg_mul_in_rsc, // @[:@11377.4]
  input  [1:0]  io_cfg_out_precision, // @[:@11377.4]
  input  [5:0]  io_cfg_truncate, // @[:@11377.4]
  input         io_chn_alu_in_rsc_valid, // @[:@11377.4]
  input  [15:0] io_chn_alu_in_rsc_bits, // @[:@11377.4]
  input         io_chn_data_in_rsc_valid, // @[:@11377.4]
  input  [16:0] io_chn_data_in_rsc_bits, // @[:@11377.4]
  output [15:0] io_chn_data_out_rsc_bits // @[:@11377.4]
);
  wire  NV_NVDLA_BC_pipe_reset; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_io_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_io_vi; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_io_ro; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire [17:0] NV_NVDLA_BC_pipe_io_di; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_io_vo; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_io_ri; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire [17:0] NV_NVDLA_BC_pipe_io_dout; // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
  wire  NV_NVDLA_BC_pipe_1_reset; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire  NV_NVDLA_BC_pipe_1_io_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire  NV_NVDLA_BC_pipe_1_io_vi; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire  NV_NVDLA_BC_pipe_1_io_ro; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire [33:0] NV_NVDLA_BC_pipe_1_io_di; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire  NV_NVDLA_BC_pipe_1_io_vo; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire  NV_NVDLA_BC_pipe_1_io_ri; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire [33:0] NV_NVDLA_BC_pipe_1_io_dout; // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
  wire [33:0] NV_NVDLA_HLS_shiftrightsu_io_data_in; // @[NV_NVDLA_CDMA_CVT_cell.scala 80:33:@11417.4]
  wire [5:0] NV_NVDLA_HLS_shiftrightsu_io_shift_num; // @[NV_NVDLA_CDMA_CVT_cell.scala 80:33:@11417.4]
  wire [16:0] NV_NVDLA_HLS_shiftrightsu_io_data_out; // @[NV_NVDLA_CDMA_CVT_cell.scala 80:33:@11417.4]
  wire [16:0] NV_NVDLA_HLS_saturate_io_data_in; // @[NV_NVDLA_CDMA_CVT_cell.scala 85:34:@11422.4]
  wire [15:0] NV_NVDLA_HLS_saturate_io_data_out; // @[NV_NVDLA_CDMA_CVT_cell.scala 85:34:@11422.4]
  wire [16:0] NV_NVDLA_HLS_saturate_1_io_data_in; // @[NV_NVDLA_CDMA_CVT_cell.scala 89:33:@11426.4]
  wire [7:0] NV_NVDLA_HLS_saturate_1_io_data_out; // @[NV_NVDLA_CDMA_CVT_cell.scala 89:33:@11426.4]
  wire  NV_NVDLA_BC_pipe_2_reset; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire  NV_NVDLA_BC_pipe_2_io_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire  NV_NVDLA_BC_pipe_2_io_vi; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire  NV_NVDLA_BC_pipe_2_io_ro; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire [15:0] NV_NVDLA_BC_pipe_2_io_di; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire  NV_NVDLA_BC_pipe_2_io_ri; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire [15:0] NV_NVDLA_BC_pipe_2_io_dout; // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
  wire [16:0] _T_49; // @[NV_NVDLA_CDMA_CVT_cell.scala 53:45:@11385.4]
  wire [15:0] _T_52; // @[NV_NVDLA_CDMA_CVT_cell.scala 55:43:@11388.4]
  wire [17:0] _T_48; // @[NV_NVDLA_CDMA_CVT_cell.scala 52:28:@11384.4 NV_NVDLA_CDMA_CVT_cell.scala 53:18:@11386.4]
  wire [17:0] _T_51; // @[NV_NVDLA_CDMA_CVT_cell.scala 54:27:@11387.4 NV_NVDLA_CDMA_CVT_cell.scala 55:17:@11389.4]
  wire [18:0] _T_56; // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11398.4]
  wire [17:0] _T_57; // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11399.4]
  wire [17:0] _T_58; // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11400.4]
  wire [17:0] _T_62; // @[NV_NVDLA_CDMA_CVT_cell.scala 74:36:@11411.4]
  wire [15:0] _T_63; // @[NV_NVDLA_CDMA_CVT_cell.scala 74:64:@11412.4]
  wire [17:0] _GEN_0; // @[NV_NVDLA_CDMA_CVT_cell.scala 74:43:@11413.4]
  wire [33:0] _T_64; // @[NV_NVDLA_CDMA_CVT_cell.scala 74:43:@11413.4]
  wire  _T_67; // @[NV_NVDLA_CDMA_CVT_cell.scala 97:48:@11436.4]
  NV_NVDLA_BC_pipe NV_NVDLA_BC_pipe ( // @[NV_NVDLA_CDMA_CVT_cell.scala 59:25:@11391.4]
    .reset(NV_NVDLA_BC_pipe_reset),
    .io_clk(NV_NVDLA_BC_pipe_io_clk),
    .io_vi(NV_NVDLA_BC_pipe_io_vi),
    .io_ro(NV_NVDLA_BC_pipe_io_ro),
    .io_di(NV_NVDLA_BC_pipe_io_di),
    .io_vo(NV_NVDLA_BC_pipe_io_vo),
    .io_ri(NV_NVDLA_BC_pipe_io_ri),
    .io_dout(NV_NVDLA_BC_pipe_io_dout)
  );
  NV_NVDLA_BC_pipe_1 NV_NVDLA_BC_pipe_1 ( // @[NV_NVDLA_CDMA_CVT_cell.scala 70:25:@11405.4]
    .reset(NV_NVDLA_BC_pipe_1_reset),
    .io_clk(NV_NVDLA_BC_pipe_1_io_clk),
    .io_vi(NV_NVDLA_BC_pipe_1_io_vi),
    .io_ro(NV_NVDLA_BC_pipe_1_io_ro),
    .io_di(NV_NVDLA_BC_pipe_1_io_di),
    .io_vo(NV_NVDLA_BC_pipe_1_io_vo),
    .io_ri(NV_NVDLA_BC_pipe_1_io_ri),
    .io_dout(NV_NVDLA_BC_pipe_1_io_dout)
  );
  NV_soDLA_HLS_shiftrightsu NV_soDLA_HLS_shiftrightsu ( // @[NV_NVDLA_CDMA_CVT_cell.scala 80:33:@11417.4]
    .io_data_in(NV_NVDLA_HLS_shiftrightsu_io_data_in),
    .io_shift_num(NV_NVDLA_HLS_shiftrightsu_io_shift_num),
    .io_data_out(NV_NVDLA_HLS_shiftrightsu_io_data_out)
  );
  NV_soDLA_HLS_saturate NV_soDLA_HLS_saturate ( // @[NV_NVDLA_CDMA_CVT_cell.scala 85:34:@11422.4]
    .io_data_in(NV_NVDLA_HLS_saturate_io_data_in),
    .io_data_out(NV_NVDLA_HLS_saturate_io_data_out)
  );
  NV_soDLA_HLS_saturate_1 NV_soDLA_HLS_saturate_1 ( // @[NV_NVDLA_CDMA_CVT_cell.scala 89:33:@11426.4]
    .io_data_in(NV_NVDLA_HLS_saturate_1_io_data_in),
    .io_data_out(NV_NVDLA_HLS_saturate_1_io_data_out)
  );
  NV_NVDLA_BC_pipe_2 NV_NVDLA_BC_pipe_2 ( // @[NV_NVDLA_CDMA_CVT_cell.scala 93:25:@11430.4]
    .reset(NV_NVDLA_BC_pipe_2_reset),
    .io_clk(NV_NVDLA_BC_pipe_2_io_clk),
    .io_vi(NV_NVDLA_BC_pipe_2_io_vi),
    .io_ro(NV_NVDLA_BC_pipe_2_io_ro),
    .io_di(NV_NVDLA_BC_pipe_2_io_di),
    .io_ri(NV_NVDLA_BC_pipe_2_io_ri),
    .io_dout(NV_NVDLA_BC_pipe_2_io_dout)
  );
  assign _T_49 = $signed(io_chn_data_in_rsc_bits); // @[NV_NVDLA_CDMA_CVT_cell.scala 53:45:@11385.4]
  assign _T_52 = $signed(io_chn_alu_in_rsc_bits); // @[NV_NVDLA_CDMA_CVT_cell.scala 55:43:@11388.4]
  assign _T_48 = {{1{_T_49[16]}},_T_49}; // @[NV_NVDLA_CDMA_CVT_cell.scala 52:28:@11384.4 NV_NVDLA_CDMA_CVT_cell.scala 53:18:@11386.4]
  assign _T_51 = {{2{_T_52[15]}},_T_52}; // @[NV_NVDLA_CDMA_CVT_cell.scala 54:27:@11387.4 NV_NVDLA_CDMA_CVT_cell.scala 55:17:@11389.4]
  assign _T_56 = $signed(_T_48) - $signed(_T_51); // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11398.4]
  assign _T_57 = $signed(_T_48) - $signed(_T_51); // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11399.4]
  assign _T_58 = $signed(_T_57); // @[NV_NVDLA_CDMA_CVT_cell.scala 63:36:@11400.4]
  assign _T_62 = $signed(NV_NVDLA_BC_pipe_io_dout); // @[NV_NVDLA_CDMA_CVT_cell.scala 74:36:@11411.4]
  assign _T_63 = $signed(io_cfg_mul_in_rsc); // @[NV_NVDLA_CDMA_CVT_cell.scala 74:64:@11412.4]
  assign _GEN_0 = {{2{_T_63[15]}},_T_63}; // @[NV_NVDLA_CDMA_CVT_cell.scala 74:43:@11413.4]
  assign _T_64 = $signed(_T_62) * $signed(_GEN_0); // @[NV_NVDLA_CDMA_CVT_cell.scala 74:43:@11413.4]
  assign _T_67 = io_cfg_out_precision == 2'h1; // @[NV_NVDLA_CDMA_CVT_cell.scala 97:48:@11436.4]
  assign io_chn_data_out_rsc_bits = NV_NVDLA_BC_pipe_2_io_dout; // @[NV_NVDLA_CDMA_CVT_cell.scala 100:31:@11441.4]
  assign NV_NVDLA_BC_pipe_reset = reset; // @[:@11393.4]
  assign NV_NVDLA_BC_pipe_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 60:20:@11394.4]
  assign NV_NVDLA_BC_pipe_io_vi = io_chn_alu_in_rsc_valid & io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_CVT_cell.scala 61:19:@11396.4]
  assign NV_NVDLA_BC_pipe_io_di = $unsigned(_T_58); // @[NV_NVDLA_CDMA_CVT_cell.scala 63:19:@11402.4]
  assign NV_NVDLA_BC_pipe_io_ri = NV_NVDLA_BC_pipe_1_io_ro; // @[NV_NVDLA_CDMA_CVT_cell.scala 65:19:@11403.4]
  assign NV_NVDLA_BC_pipe_1_reset = reset; // @[:@11407.4]
  assign NV_NVDLA_BC_pipe_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 71:20:@11408.4]
  assign NV_NVDLA_BC_pipe_1_io_vi = NV_NVDLA_BC_pipe_io_vo; // @[NV_NVDLA_CDMA_CVT_cell.scala 72:19:@11409.4]
  assign NV_NVDLA_BC_pipe_1_io_di = $unsigned(_T_64); // @[NV_NVDLA_CDMA_CVT_cell.scala 74:19:@11415.4]
  assign NV_NVDLA_BC_pipe_1_io_ri = NV_NVDLA_BC_pipe_2_io_ro; // @[NV_NVDLA_CDMA_CVT_cell.scala 76:19:@11416.4]
  assign NV_NVDLA_HLS_shiftrightsu_io_data_in = NV_NVDLA_BC_pipe_1_io_dout; // @[NV_NVDLA_CDMA_CVT_cell.scala 81:32:@11420.4]
  assign NV_NVDLA_HLS_shiftrightsu_io_shift_num = io_cfg_truncate; // @[NV_NVDLA_CDMA_CVT_cell.scala 82:34:@11421.4]
  assign NV_NVDLA_HLS_saturate_io_data_in = NV_NVDLA_HLS_shiftrightsu_io_data_out; // @[NV_NVDLA_CDMA_CVT_cell.scala 86:33:@11425.4]
  assign NV_NVDLA_HLS_saturate_1_io_data_in = NV_NVDLA_HLS_shiftrightsu_io_data_out; // @[NV_NVDLA_CDMA_CVT_cell.scala 90:32:@11429.4]
  assign NV_NVDLA_BC_pipe_2_reset = reset; // @[:@11432.4]
  assign NV_NVDLA_BC_pipe_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_CVT_cell.scala 94:20:@11433.4]
  assign NV_NVDLA_BC_pipe_2_io_vi = NV_NVDLA_BC_pipe_1_io_vo; // @[NV_NVDLA_CDMA_CVT_cell.scala 95:19:@11434.4]
  assign NV_NVDLA_BC_pipe_2_io_di = _T_67 ? NV_NVDLA_HLS_saturate_io_data_out : {{8'd0}, NV_NVDLA_HLS_saturate_1_io_data_out}; // @[NV_NVDLA_CDMA_CVT_cell.scala 97:19:@11438.4]
  assign NV_NVDLA_BC_pipe_2_io_ri = 1'h1; // @[NV_NVDLA_CDMA_CVT_cell.scala 99:19:@11440.4]
endmodule
module NV_NVDLA_CDMA_cvt( // @[:@20092.2]
  input          reset, // @[:@20094.4]
  input          io_nvdla_core_clk, // @[:@20095.4]
  input          io_nvdla_core_ng_clk, // @[:@20095.4]
  input          io_nvdla_hls_clk, // @[:@20095.4]
  input          io_dc2cvt_dat_wr_sel, // @[:@20095.4]
  input          io_dc2cvt_dat_wr_addr_valid, // @[:@20095.4]
  input  [16:0]  io_dc2cvt_dat_wr_addr_bits, // @[:@20095.4]
  input  [255:0] io_dc2cvt_dat_wr_data, // @[:@20095.4]
  input  [11:0]  io_dc2cvt_dat_wr_info_pd, // @[:@20095.4]
  input          io_img2cvt_dat_wr_sel, // @[:@20095.4]
  input          io_img2cvt_dat_wr_addr_valid, // @[:@20095.4]
  input  [16:0]  io_img2cvt_dat_wr_addr_bits, // @[:@20095.4]
  input  [255:0] io_img2cvt_dat_wr_data, // @[:@20095.4]
  input  [511:0] io_img2cvt_mn_wr_data, // @[:@20095.4]
  input  [31:0]  io_img2cvt_dat_wr_pad_mask, // @[:@20095.4]
  input  [11:0]  io_img2cvt_dat_wr_info_pd, // @[:@20095.4]
  output [1:0]   io_cdma2buf_dat_wr_sel, // @[:@20095.4]
  output         io_cdma2buf_dat_wr_addr_valid, // @[:@20095.4]
  output [16:0]  io_cdma2buf_dat_wr_addr_bits, // @[:@20095.4]
  output [255:0] io_cdma2buf_dat_wr_data, // @[:@20095.4]
  input          io_reg2dp_op_en, // @[:@20095.4]
  input  [1:0]   io_reg2dp_proc_precision, // @[:@20095.4]
  input          io_reg2dp_cvt_en, // @[:@20095.4]
  input  [5:0]   io_reg2dp_cvt_truncate, // @[:@20095.4]
  input  [15:0]  io_reg2dp_cvt_offset, // @[:@20095.4]
  input  [15:0]  io_reg2dp_cvt_scale, // @[:@20095.4]
  input  [15:0]  io_reg2dp_pad_value, // @[:@20095.4]
  input          io_dp2reg_done, // @[:@20095.4]
  output         io_dp2reg_dat_flush_done // @[:@20095.4]
);
  wire  NV_NVDLA_CDMA_CVT_cell_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire  NV_NVDLA_CDMA_CVT_cell_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire  NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire  NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
  wire  NV_NVDLA_CDMA_CVT_cell_1_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire  NV_NVDLA_CDMA_CVT_cell_1_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_1_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_1_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_1_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire  NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire  NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
  wire  NV_NVDLA_CDMA_CVT_cell_2_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire  NV_NVDLA_CDMA_CVT_cell_2_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_2_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_2_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_2_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire  NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire  NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
  wire  NV_NVDLA_CDMA_CVT_cell_3_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire  NV_NVDLA_CDMA_CVT_cell_3_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_3_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_3_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_3_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire  NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire  NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
  wire  NV_NVDLA_CDMA_CVT_cell_4_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire  NV_NVDLA_CDMA_CVT_cell_4_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_4_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_4_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_4_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire  NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire  NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
  wire  NV_NVDLA_CDMA_CVT_cell_5_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire  NV_NVDLA_CDMA_CVT_cell_5_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_5_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_5_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_5_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire  NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire  NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
  wire  NV_NVDLA_CDMA_CVT_cell_6_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire  NV_NVDLA_CDMA_CVT_cell_6_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_6_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_6_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_6_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire  NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire  NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
  wire  NV_NVDLA_CDMA_CVT_cell_7_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire  NV_NVDLA_CDMA_CVT_cell_7_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_7_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_7_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_7_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire  NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire  NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
  wire  NV_NVDLA_CDMA_CVT_cell_8_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire  NV_NVDLA_CDMA_CVT_cell_8_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_8_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_8_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_8_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire  NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire  NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
  wire  NV_NVDLA_CDMA_CVT_cell_9_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire  NV_NVDLA_CDMA_CVT_cell_9_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_9_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_9_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_9_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire  NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire  NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
  wire  NV_NVDLA_CDMA_CVT_cell_10_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire  NV_NVDLA_CDMA_CVT_cell_10_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_10_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_10_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_10_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire  NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire  NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
  wire  NV_NVDLA_CDMA_CVT_cell_11_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire  NV_NVDLA_CDMA_CVT_cell_11_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_11_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_11_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_11_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire  NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire  NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
  wire  NV_NVDLA_CDMA_CVT_cell_12_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire  NV_NVDLA_CDMA_CVT_cell_12_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_12_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_12_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_12_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire  NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire  NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
  wire  NV_NVDLA_CDMA_CVT_cell_13_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire  NV_NVDLA_CDMA_CVT_cell_13_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_13_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_13_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_13_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire  NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire  NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
  wire  NV_NVDLA_CDMA_CVT_cell_14_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire  NV_NVDLA_CDMA_CVT_cell_14_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_14_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_14_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_14_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire  NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire  NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
  wire  NV_NVDLA_CDMA_CVT_cell_15_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire  NV_NVDLA_CDMA_CVT_cell_15_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_15_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_15_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_15_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire  NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire  NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
  wire  NV_NVDLA_CDMA_CVT_cell_16_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire  NV_NVDLA_CDMA_CVT_cell_16_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_16_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_16_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_16_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire  NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire  NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
  wire  NV_NVDLA_CDMA_CVT_cell_17_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire  NV_NVDLA_CDMA_CVT_cell_17_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_17_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_17_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_17_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire  NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire  NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
  wire  NV_NVDLA_CDMA_CVT_cell_18_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire  NV_NVDLA_CDMA_CVT_cell_18_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_18_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_18_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_18_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire  NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire  NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
  wire  NV_NVDLA_CDMA_CVT_cell_19_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire  NV_NVDLA_CDMA_CVT_cell_19_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_19_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_19_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_19_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire  NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire  NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
  wire  NV_NVDLA_CDMA_CVT_cell_20_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire  NV_NVDLA_CDMA_CVT_cell_20_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_20_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_20_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_20_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire  NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire  NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
  wire  NV_NVDLA_CDMA_CVT_cell_21_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire  NV_NVDLA_CDMA_CVT_cell_21_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_21_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_21_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_21_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire  NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire  NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
  wire  NV_NVDLA_CDMA_CVT_cell_22_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire  NV_NVDLA_CDMA_CVT_cell_22_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_22_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_22_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_22_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire  NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire  NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
  wire  NV_NVDLA_CDMA_CVT_cell_23_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire  NV_NVDLA_CDMA_CVT_cell_23_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_23_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_23_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_23_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire  NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire  NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
  wire  NV_NVDLA_CDMA_CVT_cell_24_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire  NV_NVDLA_CDMA_CVT_cell_24_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_24_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_24_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_24_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire  NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire  NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
  wire  NV_NVDLA_CDMA_CVT_cell_25_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire  NV_NVDLA_CDMA_CVT_cell_25_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_25_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_25_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_25_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire  NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire  NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
  wire  NV_NVDLA_CDMA_CVT_cell_26_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire  NV_NVDLA_CDMA_CVT_cell_26_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_26_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_26_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_26_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire  NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire  NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
  wire  NV_NVDLA_CDMA_CVT_cell_27_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire  NV_NVDLA_CDMA_CVT_cell_27_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_27_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_27_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_27_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire  NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire  NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
  wire  NV_NVDLA_CDMA_CVT_cell_28_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire  NV_NVDLA_CDMA_CVT_cell_28_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_28_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_28_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_28_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire  NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire  NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
  wire  NV_NVDLA_CDMA_CVT_cell_29_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire  NV_NVDLA_CDMA_CVT_cell_29_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_29_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_29_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_29_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire  NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire  NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
  wire  NV_NVDLA_CDMA_CVT_cell_30_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire  NV_NVDLA_CDMA_CVT_cell_30_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_30_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_30_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_30_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire  NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire  NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
  wire  NV_NVDLA_CDMA_CVT_cell_31_reset; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire  NV_NVDLA_CDMA_CVT_cell_31_io_nvdla_core_clk; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_31_io_cfg_mul_in_rsc; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [1:0] NV_NVDLA_CDMA_CVT_cell_31_io_cfg_out_precision; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [5:0] NV_NVDLA_CDMA_CVT_cell_31_io_cfg_truncate; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire  NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire  NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_valid; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [16:0] NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  wire [15:0] NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
  reg  _T_89; // @[NV_NVDLA_CDMA_cvt.scala 77:20:@20097.4]
  reg [31:0] _RAND_0;
  reg [1:0] _T_92; // @[NV_NVDLA_CDMA_cvt.scala 78:33:@20098.4]
  reg [31:0] _RAND_1;
  reg [15:0] _T_95; // @[NV_NVDLA_CDMA_cvt.scala 79:24:@20099.4]
  reg [31:0] _RAND_2;
  reg [5:0] _T_98; // @[NV_NVDLA_CDMA_cvt.scala 80:27:@20100.4]
  reg [31:0] _RAND_3;
  reg [15:0] _T_101; // @[NV_NVDLA_CDMA_cvt.scala 81:25:@20101.4]
  reg [31:0] _RAND_4;
  reg [5:0] _T_104; // @[NV_NVDLA_CDMA_cvt.scala 82:25:@20102.4]
  reg [31:0] _RAND_5;
  reg [15:0] _T_113; // @[NV_NVDLA_CDMA_cvt.scala 85:28:@20105.4]
  reg [31:0] _RAND_6;
  wire  _T_126; // @[NV_NVDLA_CDMA_cvt.scala 91:15:@20110.4]
  wire  _T_127; // @[NV_NVDLA_CDMA_cvt.scala 91:31:@20111.4]
  wire  _T_128; // @[NV_NVDLA_CDMA_cvt.scala 92:28:@20112.4]
  wire  _T_129; // @[NV_NVDLA_CDMA_cvt.scala 92:26:@20113.4]
  wire [5:0] _T_140; // @[Bitwise.scala 72:12:@20125.6]
  wire [1:0] _GEN_0; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [15:0] _GEN_1; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [5:0] _GEN_2; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [15:0] _GEN_3; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [5:0] _GEN_4; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [15:0] _GEN_7; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  wire [11:0] _T_153; // @[Bitwise.scala 72:12:@20150.4]
  wire [11:0] _T_154; // @[NV_NVDLA_CDMA_cvt.scala 127:61:@20151.4]
  wire [11:0] _T_158; // @[Bitwise.scala 72:12:@20153.4]
  wire [11:0] _T_159; // @[NV_NVDLA_CDMA_cvt.scala 128:62:@20154.4]
  wire [11:0] _T_160; // @[NV_NVDLA_CDMA_cvt.scala 127:88:@20155.4]
  wire [3:0] _T_161; // @[NV_NVDLA_CDMA_cvt.scala 130:33:@20156.4]
  wire  _T_162; // @[NV_NVDLA_CDMA_cvt.scala 131:33:@20157.4]
  wire  _T_163; // @[NV_NVDLA_CDMA_cvt.scala 132:33:@20158.4]
  wire  _T_165; // @[NV_NVDLA_CDMA_cvt.scala 135:46:@20160.4]
  wire  _T_167; // @[NV_NVDLA_CDMA_cvt.scala 138:27:@20161.4]
  wire  _T_168; // @[NV_NVDLA_CDMA_cvt.scala 137:27:@20162.4]
  wire [31:0] _T_170; // @[NV_NVDLA_CDMA_cvt.scala 140:26:@20163.4]
  wire [16:0] _T_174; // @[Bitwise.scala 72:12:@20165.4]
  wire [16:0] _T_175; // @[NV_NVDLA_CDMA_cvt.scala 141:57:@20166.4]
  wire [16:0] _T_179; // @[Bitwise.scala 72:12:@20168.4]
  wire [16:0] _T_180; // @[NV_NVDLA_CDMA_cvt.scala 142:58:@20169.4]
  wire [16:0] _T_181; // @[NV_NVDLA_CDMA_cvt.scala 141:86:@20170.4]
  wire [255:0] _T_185; // @[Bitwise.scala 72:12:@20172.4]
  wire [255:0] _T_186; // @[NV_NVDLA_CDMA_cvt.scala 143:79:@20173.4]
  wire [255:0] _T_190; // @[Bitwise.scala 72:12:@20175.4]
  wire [255:0] _T_191; // @[NV_NVDLA_CDMA_cvt.scala 144:80:@20176.4]
  wire [255:0] _T_192; // @[NV_NVDLA_CDMA_cvt.scala 143:103:@20177.4]
  wire  _T_195; // @[NV_NVDLA_CDMA_cvt.scala 155:45:@20179.4]
  wire  _T_196; // @[NV_NVDLA_CDMA_cvt.scala 155:33:@20180.4]
  wire  _T_197; // @[NV_NVDLA_CDMA_cvt.scala 155:98:@20181.4]
  wire [31:0] _T_201; // @[Bitwise.scala 72:12:@20183.4]
  wire [31:0] _T_203; // @[NV_NVDLA_CDMA_cvt.scala 155:22:@20184.4]
  reg  _T_206; // @[NV_NVDLA_CDMA_cvt.scala 160:27:@20185.4]
  reg [31:0] _RAND_7;
  reg  _T_209; // @[NV_NVDLA_CDMA_cvt.scala 161:29:@20186.4]
  reg [31:0] _RAND_8;
  reg  _T_212; // @[NV_NVDLA_CDMA_cvt.scala 162:29:@20187.4]
  reg [31:0] _RAND_9;
  reg [511:0] _T_214; // @[NV_NVDLA_CDMA_cvt.scala 163:30:@20188.4]
  reg [511:0] _RAND_10;
  reg [255:0] _T_216; // @[NV_NVDLA_CDMA_cvt.scala 164:25:@20189.4]
  reg [255:0] _RAND_11;
  reg [31:0] _T_219; // @[NV_NVDLA_CDMA_cvt.scala 165:29:@20190.4]
  reg [31:0] _RAND_12;
  reg  _T_222; // @[NV_NVDLA_CDMA_cvt.scala 166:29:@20191.4]
  reg [31:0] _RAND_13;
  reg  _T_225; // @[NV_NVDLA_CDMA_cvt.scala 167:33:@20192.4]
  reg [31:0] _RAND_14;
  reg [16:0] _T_228; // @[NV_NVDLA_CDMA_cvt.scala 168:30:@20193.4]
  reg [31:0] _RAND_15;
  reg [3:0] _T_231; // @[NV_NVDLA_CDMA_cvt.scala 169:33:@20194.4]
  reg [31:0] _RAND_16;
  reg [31:0] _T_234; // @[NV_NVDLA_CDMA_cvt.scala 170:34:@20195.4]
  reg [31:0] _RAND_17;
  reg [1:0] _T_237; // @[NV_NVDLA_CDMA_cvt.scala 172:34:@20196.4]
  reg [31:0] _RAND_18;
  wire [511:0] _GEN_15; // @[NV_NVDLA_CDMA_cvt.scala 184:22:@20204.6]
  wire  _GEN_16; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  wire  _GEN_17; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  wire [16:0] _GEN_18; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  wire [3:0] _GEN_19; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  wire  _T_241; // @[NV_NVDLA_CDMA_cvt.scala 189:16:@20209.4]
  wire [31:0] _GEN_22; // @[NV_NVDLA_CDMA_cvt.scala 189:31:@20210.4]
  wire [31:0] _GEN_23; // @[NV_NVDLA_CDMA_cvt.scala 194:35:@20215.4]
  wire [1:0] _GEN_24; // @[NV_NVDLA_CDMA_cvt.scala 198:20:@20218.4]
  reg [16:0] _T_245_0; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_19;
  reg [16:0] _T_245_1; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_20;
  reg [16:0] _T_245_2; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_21;
  reg [16:0] _T_245_3; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_22;
  reg [16:0] _T_245_4; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_23;
  reg [16:0] _T_245_5; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_24;
  reg [16:0] _T_245_6; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_25;
  reg [16:0] _T_245_7; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_26;
  reg [16:0] _T_245_8; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_27;
  reg [16:0] _T_245_9; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_28;
  reg [16:0] _T_245_10; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_29;
  reg [16:0] _T_245_11; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_30;
  reg [16:0] _T_245_12; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_31;
  reg [16:0] _T_245_13; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_32;
  reg [16:0] _T_245_14; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_33;
  reg [16:0] _T_245_15; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_34;
  reg [16:0] _T_245_16; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_35;
  reg [16:0] _T_245_17; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_36;
  reg [16:0] _T_245_18; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_37;
  reg [16:0] _T_245_19; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_38;
  reg [16:0] _T_245_20; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_39;
  reg [16:0] _T_245_21; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_40;
  reg [16:0] _T_245_22; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_41;
  reg [16:0] _T_245_23; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_42;
  reg [16:0] _T_245_24; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_43;
  reg [16:0] _T_245_25; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_44;
  reg [16:0] _T_245_26; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_45;
  reg [16:0] _T_245_27; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_46;
  reg [16:0] _T_245_28; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_47;
  reg [16:0] _T_245_29; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_48;
  reg [16:0] _T_245_30; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_49;
  reg [16:0] _T_245_31; // @[NV_NVDLA_CDMA_cvt.scala 207:22:@20222.4]
  reg [31:0] _RAND_50;
  reg [15:0] _T_283_0; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_51;
  reg [15:0] _T_283_1; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_52;
  reg [15:0] _T_283_2; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_53;
  reg [15:0] _T_283_3; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_54;
  reg [15:0] _T_283_4; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_55;
  reg [15:0] _T_283_5; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_56;
  reg [15:0] _T_283_6; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_57;
  reg [15:0] _T_283_7; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_58;
  reg [15:0] _T_283_8; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_59;
  reg [15:0] _T_283_9; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_60;
  reg [15:0] _T_283_10; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_61;
  reg [15:0] _T_283_11; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_62;
  reg [15:0] _T_283_12; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_63;
  reg [15:0] _T_283_13; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_64;
  reg [15:0] _T_283_14; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_65;
  reg [15:0] _T_283_15; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_66;
  reg [15:0] _T_283_16; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_67;
  reg [15:0] _T_283_17; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_68;
  reg [15:0] _T_283_18; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_69;
  reg [15:0] _T_283_19; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_70;
  reg [15:0] _T_283_20; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_71;
  reg [15:0] _T_283_21; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_72;
  reg [15:0] _T_283_22; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_73;
  reg [15:0] _T_283_23; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_74;
  reg [15:0] _T_283_24; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_75;
  reg [15:0] _T_283_25; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_76;
  reg [15:0] _T_283_26; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_77;
  reg [15:0] _T_283_27; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_283_28; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_283_29; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_283_30; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_81;
  reg [15:0] _T_283_31; // @[NV_NVDLA_CDMA_cvt.scala 208:22:@20223.4]
  reg [31:0] _RAND_82;
  wire  _T_432; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20227.4]
  wire  _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:69:@20228.4]
  wire  _T_434; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20229.4]
  wire [8:0] _T_438; // @[Bitwise.scala 72:12:@20232.4]
  wire [7:0] _T_439; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20233.4]
  wire [16:0] _T_440; // @[Cat.scala 30:58:@20234.4]
  wire [15:0] _T_441; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20236.4]
  wire [15:0] _T_443; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20238.4]
  wire  _T_444; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20240.4]
  wire  _T_445; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20245.4]
  wire  _T_447; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20247.4]
  wire [8:0] _T_451; // @[Bitwise.scala 72:12:@20250.4]
  wire [7:0] _T_452; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20251.4]
  wire [16:0] _T_453; // @[Cat.scala 30:58:@20252.4]
  wire [15:0] _T_454; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20254.4]
  wire [15:0] _T_456; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20256.4]
  wire  _T_457; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20258.4]
  wire  _T_458; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20263.4]
  wire  _T_460; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20265.4]
  wire [8:0] _T_464; // @[Bitwise.scala 72:12:@20268.4]
  wire [7:0] _T_465; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20269.4]
  wire [16:0] _T_466; // @[Cat.scala 30:58:@20270.4]
  wire [15:0] _T_467; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20272.4]
  wire [15:0] _T_469; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20274.4]
  wire  _T_470; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20276.4]
  wire  _T_471; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20281.4]
  wire  _T_473; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20283.4]
  wire [8:0] _T_477; // @[Bitwise.scala 72:12:@20286.4]
  wire [7:0] _T_478; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20287.4]
  wire [16:0] _T_479; // @[Cat.scala 30:58:@20288.4]
  wire [15:0] _T_480; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20290.4]
  wire [15:0] _T_482; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20292.4]
  wire  _T_483; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20294.4]
  wire  _T_484; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20299.4]
  wire  _T_486; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20301.4]
  wire [8:0] _T_490; // @[Bitwise.scala 72:12:@20304.4]
  wire [7:0] _T_491; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20305.4]
  wire [16:0] _T_492; // @[Cat.scala 30:58:@20306.4]
  wire [15:0] _T_493; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20308.4]
  wire [15:0] _T_495; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20310.4]
  wire  _T_496; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20312.4]
  wire  _T_497; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20317.4]
  wire  _T_499; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20319.4]
  wire [8:0] _T_503; // @[Bitwise.scala 72:12:@20322.4]
  wire [7:0] _T_504; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20323.4]
  wire [16:0] _T_505; // @[Cat.scala 30:58:@20324.4]
  wire [15:0] _T_506; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20326.4]
  wire [15:0] _T_508; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20328.4]
  wire  _T_509; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20330.4]
  wire  _T_510; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20335.4]
  wire  _T_512; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20337.4]
  wire [8:0] _T_516; // @[Bitwise.scala 72:12:@20340.4]
  wire [7:0] _T_517; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20341.4]
  wire [16:0] _T_518; // @[Cat.scala 30:58:@20342.4]
  wire [15:0] _T_519; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20344.4]
  wire [15:0] _T_521; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20346.4]
  wire  _T_522; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20348.4]
  wire  _T_523; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20353.4]
  wire  _T_525; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20355.4]
  wire [8:0] _T_529; // @[Bitwise.scala 72:12:@20358.4]
  wire [7:0] _T_530; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20359.4]
  wire [16:0] _T_531; // @[Cat.scala 30:58:@20360.4]
  wire [15:0] _T_532; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20362.4]
  wire [15:0] _T_534; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20364.4]
  wire  _T_535; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20366.4]
  wire  _T_536; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20371.4]
  wire  _T_538; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20373.4]
  wire [8:0] _T_542; // @[Bitwise.scala 72:12:@20376.4]
  wire [7:0] _T_543; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20377.4]
  wire [16:0] _T_544; // @[Cat.scala 30:58:@20378.4]
  wire [15:0] _T_545; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20380.4]
  wire [15:0] _T_547; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20382.4]
  wire  _T_548; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20384.4]
  wire  _T_549; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20389.4]
  wire  _T_551; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20391.4]
  wire [8:0] _T_555; // @[Bitwise.scala 72:12:@20394.4]
  wire [7:0] _T_556; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20395.4]
  wire [16:0] _T_557; // @[Cat.scala 30:58:@20396.4]
  wire [15:0] _T_558; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20398.4]
  wire [15:0] _T_560; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20400.4]
  wire  _T_561; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20402.4]
  wire  _T_562; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20407.4]
  wire  _T_564; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20409.4]
  wire [8:0] _T_568; // @[Bitwise.scala 72:12:@20412.4]
  wire [7:0] _T_569; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20413.4]
  wire [16:0] _T_570; // @[Cat.scala 30:58:@20414.4]
  wire [15:0] _T_571; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20416.4]
  wire [15:0] _T_573; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20418.4]
  wire  _T_574; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20420.4]
  wire  _T_575; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20425.4]
  wire  _T_577; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20427.4]
  wire [8:0] _T_581; // @[Bitwise.scala 72:12:@20430.4]
  wire [7:0] _T_582; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20431.4]
  wire [16:0] _T_583; // @[Cat.scala 30:58:@20432.4]
  wire [15:0] _T_584; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20434.4]
  wire [15:0] _T_586; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20436.4]
  wire  _T_587; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20438.4]
  wire  _T_588; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20443.4]
  wire  _T_590; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20445.4]
  wire [8:0] _T_594; // @[Bitwise.scala 72:12:@20448.4]
  wire [7:0] _T_595; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20449.4]
  wire [16:0] _T_596; // @[Cat.scala 30:58:@20450.4]
  wire [15:0] _T_597; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20452.4]
  wire [15:0] _T_599; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20454.4]
  wire  _T_600; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20456.4]
  wire  _T_601; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20461.4]
  wire  _T_603; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20463.4]
  wire [8:0] _T_607; // @[Bitwise.scala 72:12:@20466.4]
  wire [7:0] _T_608; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20467.4]
  wire [16:0] _T_609; // @[Cat.scala 30:58:@20468.4]
  wire [15:0] _T_610; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20470.4]
  wire [15:0] _T_612; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20472.4]
  wire  _T_613; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20474.4]
  wire  _T_614; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20479.4]
  wire  _T_616; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20481.4]
  wire [8:0] _T_620; // @[Bitwise.scala 72:12:@20484.4]
  wire [7:0] _T_621; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20485.4]
  wire [16:0] _T_622; // @[Cat.scala 30:58:@20486.4]
  wire [15:0] _T_623; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20488.4]
  wire [15:0] _T_625; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20490.4]
  wire  _T_626; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20492.4]
  wire  _T_627; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20497.4]
  wire  _T_629; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20499.4]
  wire [8:0] _T_633; // @[Bitwise.scala 72:12:@20502.4]
  wire [7:0] _T_634; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20503.4]
  wire [16:0] _T_635; // @[Cat.scala 30:58:@20504.4]
  wire [15:0] _T_636; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20506.4]
  wire [15:0] _T_638; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20508.4]
  wire  _T_639; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20510.4]
  wire  _T_640; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20515.4]
  wire  _T_642; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20517.4]
  wire [8:0] _T_646; // @[Bitwise.scala 72:12:@20520.4]
  wire [7:0] _T_647; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20521.4]
  wire [16:0] _T_648; // @[Cat.scala 30:58:@20522.4]
  wire [15:0] _T_649; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20524.4]
  wire [15:0] _T_651; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20526.4]
  wire  _T_652; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20528.4]
  wire  _T_653; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20533.4]
  wire  _T_655; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20535.4]
  wire [8:0] _T_659; // @[Bitwise.scala 72:12:@20538.4]
  wire [7:0] _T_660; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20539.4]
  wire [16:0] _T_661; // @[Cat.scala 30:58:@20540.4]
  wire [15:0] _T_662; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20542.4]
  wire [15:0] _T_664; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20544.4]
  wire  _T_665; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20546.4]
  wire  _T_666; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20551.4]
  wire  _T_668; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20553.4]
  wire [8:0] _T_672; // @[Bitwise.scala 72:12:@20556.4]
  wire [7:0] _T_673; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20557.4]
  wire [16:0] _T_674; // @[Cat.scala 30:58:@20558.4]
  wire [15:0] _T_675; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20560.4]
  wire [15:0] _T_677; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20562.4]
  wire  _T_678; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20564.4]
  wire  _T_679; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20569.4]
  wire  _T_681; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20571.4]
  wire [8:0] _T_685; // @[Bitwise.scala 72:12:@20574.4]
  wire [7:0] _T_686; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20575.4]
  wire [16:0] _T_687; // @[Cat.scala 30:58:@20576.4]
  wire [15:0] _T_688; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20578.4]
  wire [15:0] _T_690; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20580.4]
  wire  _T_691; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20582.4]
  wire  _T_692; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20587.4]
  wire  _T_694; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20589.4]
  wire [8:0] _T_698; // @[Bitwise.scala 72:12:@20592.4]
  wire [7:0] _T_699; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20593.4]
  wire [16:0] _T_700; // @[Cat.scala 30:58:@20594.4]
  wire [15:0] _T_701; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20596.4]
  wire [15:0] _T_703; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20598.4]
  wire  _T_704; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20600.4]
  wire  _T_705; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20605.4]
  wire  _T_707; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20607.4]
  wire [8:0] _T_711; // @[Bitwise.scala 72:12:@20610.4]
  wire [7:0] _T_712; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20611.4]
  wire [16:0] _T_713; // @[Cat.scala 30:58:@20612.4]
  wire [15:0] _T_714; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20614.4]
  wire [15:0] _T_716; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20616.4]
  wire  _T_717; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20618.4]
  wire  _T_718; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20623.4]
  wire  _T_720; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20625.4]
  wire [8:0] _T_724; // @[Bitwise.scala 72:12:@20628.4]
  wire [7:0] _T_725; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20629.4]
  wire [16:0] _T_726; // @[Cat.scala 30:58:@20630.4]
  wire [15:0] _T_727; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20632.4]
  wire [15:0] _T_729; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20634.4]
  wire  _T_730; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20636.4]
  wire  _T_731; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20641.4]
  wire  _T_733; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20643.4]
  wire [8:0] _T_737; // @[Bitwise.scala 72:12:@20646.4]
  wire [7:0] _T_738; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20647.4]
  wire [16:0] _T_739; // @[Cat.scala 30:58:@20648.4]
  wire [15:0] _T_740; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20650.4]
  wire [15:0] _T_742; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20652.4]
  wire  _T_743; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20654.4]
  wire  _T_744; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20659.4]
  wire  _T_746; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20661.4]
  wire [8:0] _T_750; // @[Bitwise.scala 72:12:@20664.4]
  wire [7:0] _T_751; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20665.4]
  wire [16:0] _T_752; // @[Cat.scala 30:58:@20666.4]
  wire [15:0] _T_753; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20668.4]
  wire [15:0] _T_755; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20670.4]
  wire  _T_756; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20672.4]
  wire  _T_757; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20677.4]
  wire  _T_759; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20679.4]
  wire [8:0] _T_763; // @[Bitwise.scala 72:12:@20682.4]
  wire [7:0] _T_764; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20683.4]
  wire [16:0] _T_765; // @[Cat.scala 30:58:@20684.4]
  wire [15:0] _T_766; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20686.4]
  wire [15:0] _T_768; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20688.4]
  wire  _T_769; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20690.4]
  wire  _T_770; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20695.4]
  wire  _T_772; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20697.4]
  wire [8:0] _T_776; // @[Bitwise.scala 72:12:@20700.4]
  wire [7:0] _T_777; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20701.4]
  wire [16:0] _T_778; // @[Cat.scala 30:58:@20702.4]
  wire [15:0] _T_779; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20704.4]
  wire [15:0] _T_781; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20706.4]
  wire  _T_782; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20708.4]
  wire  _T_783; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20713.4]
  wire  _T_785; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20715.4]
  wire [8:0] _T_789; // @[Bitwise.scala 72:12:@20718.4]
  wire [7:0] _T_790; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20719.4]
  wire [16:0] _T_791; // @[Cat.scala 30:58:@20720.4]
  wire [15:0] _T_792; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20722.4]
  wire [15:0] _T_794; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20724.4]
  wire  _T_795; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20726.4]
  wire  _T_796; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20731.4]
  wire  _T_798; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20733.4]
  wire [8:0] _T_802; // @[Bitwise.scala 72:12:@20736.4]
  wire [7:0] _T_803; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20737.4]
  wire [16:0] _T_804; // @[Cat.scala 30:58:@20738.4]
  wire [15:0] _T_805; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20740.4]
  wire [15:0] _T_807; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20742.4]
  wire  _T_808; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20744.4]
  wire  _T_809; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20749.4]
  wire  _T_811; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20751.4]
  wire [8:0] _T_815; // @[Bitwise.scala 72:12:@20754.4]
  wire [7:0] _T_816; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20755.4]
  wire [16:0] _T_817; // @[Cat.scala 30:58:@20756.4]
  wire [15:0] _T_818; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20758.4]
  wire [15:0] _T_820; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20760.4]
  wire  _T_821; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20762.4]
  wire  _T_822; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20767.4]
  wire  _T_824; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20769.4]
  wire [8:0] _T_828; // @[Bitwise.scala 72:12:@20772.4]
  wire [7:0] _T_829; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20773.4]
  wire [16:0] _T_830; // @[Cat.scala 30:58:@20774.4]
  wire [15:0] _T_831; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20776.4]
  wire [15:0] _T_833; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20778.4]
  wire  _T_834; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20780.4]
  wire  _T_835; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20785.4]
  wire  _T_837; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20787.4]
  wire [8:0] _T_841; // @[Bitwise.scala 72:12:@20790.4]
  wire [7:0] _T_842; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20791.4]
  wire [16:0] _T_843; // @[Cat.scala 30:58:@20792.4]
  wire [15:0] _T_844; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20794.4]
  wire [15:0] _T_846; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20796.4]
  wire  _T_847; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20798.4]
  reg  _T_850; // @[NV_NVDLA_CDMA_cvt.scala 223:23:@20803.4]
  reg [31:0] _RAND_83;
  reg [31:0] _T_853; // @[NV_NVDLA_CDMA_cvt.scala 224:25:@20804.4]
  reg [31:0] _RAND_84;
  wire  _T_854; // @[NV_NVDLA_CDMA_cvt.scala 227:19:@20806.4]
  wire [31:0] _GEN_89; // @[NV_NVDLA_CDMA_cvt.scala 227:30:@20807.4]
  wire [15:0] _T_858_0; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20918.4]
  wire [7:0] _T_989; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21291.4]
  wire [15:0] _T_858_1; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20930.4]
  wire [7:0] _T_990; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21292.4]
  wire [15:0] _T_858_2; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20942.4]
  wire [7:0] _T_991; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21293.4]
  wire [15:0] _T_858_3; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20954.4]
  wire [7:0] _T_992; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21294.4]
  wire [15:0] _T_858_4; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20966.4]
  wire [7:0] _T_993; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21295.4]
  wire [15:0] _T_858_5; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20978.4]
  wire [7:0] _T_994; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21296.4]
  wire [15:0] _T_858_6; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20990.4]
  wire [7:0] _T_995; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21297.4]
  wire [15:0] _T_858_7; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21002.4]
  wire [7:0] _T_996; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21298.4]
  wire [15:0] _T_858_8; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21014.4]
  wire [7:0] _T_997; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21299.4]
  wire [15:0] _T_858_9; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21026.4]
  wire [7:0] _T_998; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21300.4]
  wire [15:0] _T_858_10; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21038.4]
  wire [7:0] _T_999; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21301.4]
  wire [15:0] _T_858_11; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21050.4]
  wire [7:0] _T_1000; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21302.4]
  wire [15:0] _T_858_12; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21062.4]
  wire [7:0] _T_1001; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21303.4]
  wire [15:0] _T_858_13; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21074.4]
  wire [7:0] _T_1002; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21304.4]
  wire [15:0] _T_858_14; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21086.4]
  wire [7:0] _T_1003; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21305.4]
  wire [15:0] _T_858_15; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21098.4]
  wire [7:0] _T_1004; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21306.4]
  wire [15:0] _T_858_16; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21110.4]
  wire [7:0] _T_1005; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21307.4]
  wire [15:0] _T_858_17; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21122.4]
  wire [7:0] _T_1006; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21308.4]
  wire [15:0] _T_858_18; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21134.4]
  wire [7:0] _T_1007; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21309.4]
  wire [15:0] _T_858_19; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21146.4]
  wire [7:0] _T_1008; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21310.4]
  wire [15:0] _T_858_20; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21158.4]
  wire [7:0] _T_1009; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21311.4]
  wire [15:0] _T_858_21; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21170.4]
  wire [7:0] _T_1010; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21312.4]
  wire [15:0] _T_858_22; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21182.4]
  wire [7:0] _T_1011; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21313.4]
  wire [15:0] _T_858_23; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21194.4]
  wire [7:0] _T_1012; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21314.4]
  wire [15:0] _T_858_24; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21206.4]
  wire [7:0] _T_1013; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21315.4]
  wire [15:0] _T_858_25; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21218.4]
  wire [7:0] _T_1014; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21316.4]
  wire [15:0] _T_858_26; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21230.4]
  wire [7:0] _T_1015; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21317.4]
  wire [15:0] _T_858_27; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21242.4]
  wire [7:0] _T_1016; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21318.4]
  wire [15:0] _T_858_28; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21254.4]
  wire [7:0] _T_1017; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21319.4]
  wire [15:0] _T_858_29; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21266.4]
  wire [7:0] _T_1018; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21320.4]
  wire [15:0] _T_858_30; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21278.4]
  wire [7:0] _T_1019; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21321.4]
  wire [15:0] _T_858_31; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21290.4]
  wire [7:0] _T_1020; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21322.4]
  wire [63:0] _T_1065; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21362.4]
  wire [127:0] _T_1073; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21370.4]
  wire [63:0] _T_1080; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21377.4]
  wire [255:0] _T_1089; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21386.4]
  reg  _T_1094; // @[NV_NVDLA_CDMA_cvt.scala 261:72:@21388.4]
  reg [31:0] _RAND_85;
  reg  _T_1097; // @[NV_NVDLA_CDMA_cvt.scala 261:72:@21389.4]
  reg [31:0] _RAND_86;
  reg  _T_1100; // @[NV_NVDLA_CDMA_cvt.scala 261:72:@21390.4]
  reg [31:0] _RAND_87;
  reg  _T_1108; // @[NV_NVDLA_CDMA_cvt.scala 263:76:@21393.4]
  reg [31:0] _RAND_88;
  reg  _T_1111; // @[NV_NVDLA_CDMA_cvt.scala 263:76:@21394.4]
  reg [31:0] _RAND_89;
  reg  _T_1114; // @[NV_NVDLA_CDMA_cvt.scala 263:76:@21395.4]
  reg [31:0] _RAND_90;
  reg  _T_1117; // @[NV_NVDLA_CDMA_cvt.scala 263:76:@21396.4]
  reg [31:0] _RAND_91;
  reg  _T_1122; // @[NV_NVDLA_CDMA_cvt.scala 265:72:@21398.4]
  reg [31:0] _RAND_92;
  reg  _T_1125; // @[NV_NVDLA_CDMA_cvt.scala 265:72:@21399.4]
  reg [31:0] _RAND_93;
  reg  _T_1128; // @[NV_NVDLA_CDMA_cvt.scala 265:72:@21400.4]
  reg [31:0] _RAND_94;
  reg  _T_1131; // @[NV_NVDLA_CDMA_cvt.scala 265:72:@21401.4]
  reg [31:0] _RAND_95;
  reg [16:0] _T_1150; // @[NV_NVDLA_CDMA_cvt.scala 270:73:@21408.4]
  reg [31:0] _RAND_96;
  reg [16:0] _T_1153; // @[NV_NVDLA_CDMA_cvt.scala 270:73:@21409.4]
  reg [31:0] _RAND_97;
  reg [16:0] _T_1156; // @[NV_NVDLA_CDMA_cvt.scala 270:73:@21410.4]
  reg [31:0] _RAND_98;
  reg [16:0] _T_1159; // @[NV_NVDLA_CDMA_cvt.scala 270:73:@21411.4]
  reg [31:0] _RAND_99;
  reg [3:0] _T_1164; // @[NV_NVDLA_CDMA_cvt.scala 272:76:@21413.4]
  reg [31:0] _RAND_100;
  reg [3:0] _T_1167; // @[NV_NVDLA_CDMA_cvt.scala 272:76:@21414.4]
  reg [31:0] _RAND_101;
  reg [3:0] _T_1170; // @[NV_NVDLA_CDMA_cvt.scala 272:76:@21415.4]
  reg [31:0] _RAND_102;
  reg [3:0] _T_1173; // @[NV_NVDLA_CDMA_cvt.scala 272:76:@21416.4]
  reg [31:0] _RAND_103;
  reg [31:0] _T_1178; // @[NV_NVDLA_CDMA_cvt.scala 274:77:@21418.4]
  reg [31:0] _RAND_104;
  reg [31:0] _T_1181; // @[NV_NVDLA_CDMA_cvt.scala 274:77:@21419.4]
  reg [31:0] _RAND_105;
  reg [31:0] _T_1184; // @[NV_NVDLA_CDMA_cvt.scala 274:77:@21420.4]
  reg [31:0] _RAND_106;
  reg [31:0] _T_1187; // @[NV_NVDLA_CDMA_cvt.scala 274:77:@21421.4]
  reg [31:0] _RAND_107;
  wire  _T_1119; // @[NV_NVDLA_CDMA_cvt.scala 264:61:@21397.4 NV_NVDLA_CDMA_cvt.scala 279:29:@21424.4]
  wire  _GEN_90; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21431.4]
  wire  _GEN_92; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21443.4]
  wire  _GEN_94; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21455.4]
  wire  _GEN_96; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21467.4]
  wire  _T_1192; // @[NV_NVDLA_CDMA_cvt.scala 303:41:@21477.4]
  wire [1:0] _T_1193; // @[NV_NVDLA_CDMA_cvt.scala 303:30:@21478.4]
  wire  _T_1195; // @[NV_NVDLA_CDMA_cvt.scala 305:25:@21480.4]
  wire [16:0] _T_1197; // @[NV_NVDLA_CDMA_cvt.scala 306:26:@21482.4]
  wire  _T_1198; // @[NV_NVDLA_CDMA_cvt.scala 307:40:@21483.4]
  wire [3:0] _T_1199; // @[NV_NVDLA_CDMA_cvt.scala 307:29:@21484.4]
  wire  _T_1200; // @[NV_NVDLA_CDMA_cvt.scala 308:40:@21485.4]
  wire  _T_1201; // @[NV_NVDLA_CDMA_cvt.scala 308:29:@21486.4]
  wire  _T_1202; // @[NV_NVDLA_CDMA_cvt.scala 309:31:@21487.4]
  wire [31:0] _T_1205; // @[NV_NVDLA_CDMA_cvt.scala 310:30:@21489.4]
  wire [31:0] _T_1206; // @[NV_NVDLA_CDMA_cvt.scala 309:30:@21490.4]
  reg [17:0] _T_1213; // @[NV_NVDLA_CDMA_cvt.scala 318:65:@21494.4]
  reg [31:0] _RAND_108;
  wire  _T_1214; // @[NV_NVDLA_CDMA_cvt.scala 320:38:@21495.4]
  wire [255:0] _T_1215; // @[NV_NVDLA_CDMA_cvt.scala 320:27:@21496.4]
  wire  _T_1216; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21497.4]
  wire [7:0] _T_1217; // @[NV_NVDLA_CDMA_cvt.scala 322:49:@21498.4]
  wire [7:0] _T_1218; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21499.4]
  wire [7:0] _T_1219; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21500.4]
  wire  _T_1220; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21501.4]
  wire [7:0] _T_1222; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21503.4]
  wire [7:0] _T_1223; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21504.4]
  wire  _T_1224; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21505.4]
  wire [7:0] _T_1226; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21507.4]
  wire [7:0] _T_1227; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21508.4]
  wire  _T_1228; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21509.4]
  wire [7:0] _T_1230; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21511.4]
  wire [7:0] _T_1231; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21512.4]
  wire  _T_1232; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21513.4]
  wire [7:0] _T_1234; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21515.4]
  wire [7:0] _T_1235; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21516.4]
  wire  _T_1236; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21517.4]
  wire [7:0] _T_1238; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21519.4]
  wire [7:0] _T_1239; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21520.4]
  wire  _T_1240; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21521.4]
  wire [7:0] _T_1242; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21523.4]
  wire [7:0] _T_1243; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21524.4]
  wire  _T_1244; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21525.4]
  wire [7:0] _T_1246; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21527.4]
  wire [7:0] _T_1247; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21528.4]
  wire  _T_1248; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21529.4]
  wire [7:0] _T_1250; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21531.4]
  wire [7:0] _T_1251; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21532.4]
  wire  _T_1252; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21533.4]
  wire [7:0] _T_1254; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21535.4]
  wire [7:0] _T_1255; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21536.4]
  wire  _T_1256; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21537.4]
  wire [7:0] _T_1258; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21539.4]
  wire [7:0] _T_1259; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21540.4]
  wire  _T_1260; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21541.4]
  wire [7:0] _T_1262; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21543.4]
  wire [7:0] _T_1263; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21544.4]
  wire  _T_1264; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21545.4]
  wire [7:0] _T_1266; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21547.4]
  wire [7:0] _T_1267; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21548.4]
  wire  _T_1268; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21549.4]
  wire [7:0] _T_1270; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21551.4]
  wire [7:0] _T_1271; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21552.4]
  wire  _T_1272; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21553.4]
  wire [7:0] _T_1274; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21555.4]
  wire [7:0] _T_1275; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21556.4]
  wire  _T_1276; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21557.4]
  wire [7:0] _T_1278; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21559.4]
  wire [7:0] _T_1279; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21560.4]
  wire  _T_1280; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21561.4]
  wire [7:0] _T_1282; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21563.4]
  wire [7:0] _T_1283; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21564.4]
  wire  _T_1284; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21565.4]
  wire [7:0] _T_1286; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21567.4]
  wire [7:0] _T_1287; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21568.4]
  wire  _T_1288; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21569.4]
  wire [7:0] _T_1290; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21571.4]
  wire [7:0] _T_1291; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21572.4]
  wire  _T_1292; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21573.4]
  wire [7:0] _T_1294; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21575.4]
  wire [7:0] _T_1295; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21576.4]
  wire  _T_1296; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21577.4]
  wire [7:0] _T_1298; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21579.4]
  wire [7:0] _T_1299; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21580.4]
  wire  _T_1300; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21581.4]
  wire [7:0] _T_1302; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21583.4]
  wire [7:0] _T_1303; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21584.4]
  wire  _T_1304; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21585.4]
  wire [7:0] _T_1306; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21587.4]
  wire [7:0] _T_1307; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21588.4]
  wire  _T_1308; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21589.4]
  wire [7:0] _T_1310; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21591.4]
  wire [7:0] _T_1311; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21592.4]
  wire  _T_1312; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21593.4]
  wire [7:0] _T_1314; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21595.4]
  wire [7:0] _T_1315; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21596.4]
  wire  _T_1316; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21597.4]
  wire [7:0] _T_1318; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21599.4]
  wire [7:0] _T_1319; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21600.4]
  wire  _T_1320; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21601.4]
  wire [7:0] _T_1322; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21603.4]
  wire [7:0] _T_1323; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21604.4]
  wire  _T_1324; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21605.4]
  wire [7:0] _T_1326; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21607.4]
  wire [7:0] _T_1327; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21608.4]
  wire  _T_1328; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21609.4]
  wire [7:0] _T_1330; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21611.4]
  wire [7:0] _T_1331; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21612.4]
  wire  _T_1332; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21613.4]
  wire [7:0] _T_1334; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21615.4]
  wire [7:0] _T_1335; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21616.4]
  wire  _T_1336; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21617.4]
  wire [7:0] _T_1338; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21619.4]
  wire [7:0] _T_1339; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21620.4]
  wire  _T_1340; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21621.4]
  wire [7:0] _T_1342; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21623.4]
  wire [7:0] _T_1343; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21624.4]
  wire [63:0] _T_1388; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21664.4]
  wire [127:0] _T_1396; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21672.4]
  wire [63:0] _T_1403; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21679.4]
  wire [255:0] _T_1412; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21688.4]
  wire  _T_1413; // @[NV_NVDLA_CDMA_cvt.scala 323:45:@21689.4]
  wire [255:0] _T_1416; // @[NV_NVDLA_CDMA_cvt.scala 323:26:@21691.4]
  reg [255:0] _T_1419; // @[NV_NVDLA_CDMA_cvt.scala 324:34:@21692.4]
  reg [255:0] _RAND_109;
  wire  _T_1444; // @[NV_NVDLA_CDMA_cvt.scala 343:44:@21716.4]
  wire  _T_1445; // @[NV_NVDLA_CDMA_cvt.scala 343:25:@21717.4]
  wire  _T_1420; // @[NV_NVDLA_CDMA_cvt.scala 325:40:@21694.4]
  wire [16:0] _T_1421; // @[NV_NVDLA_CDMA_cvt.scala 326:70:@21695.4]
  wire [16:0] _T_1422; // @[NV_NVDLA_CDMA_cvt.scala 326:29:@21696.4]
  wire  _T_1423; // @[NV_NVDLA_CDMA_cvt.scala 328:78:@21697.4]
  wire  _T_1425; // @[NV_NVDLA_CDMA_cvt.scala 328:83:@21699.4]
  wire [1:0] _T_1426; // @[Cat.scala 30:58:@21700.4]
  wire  _T_1427; // @[NV_NVDLA_CDMA_cvt.scala 329:47:@21701.4]
  wire  _T_1429; // @[NV_NVDLA_CDMA_cvt.scala 329:52:@21703.4]
  wire [1:0] _T_1430; // @[Cat.scala 30:58:@21704.4]
  wire [1:0] _T_1431; // @[NV_NVDLA_CDMA_cvt.scala 328:33:@21705.4]
  reg [1:0] _T_1434; // @[NV_NVDLA_CDMA_cvt.scala 332:67:@21706.4]
  reg [31:0] _RAND_110;
  reg  _T_1437; // @[NV_NVDLA_CDMA_cvt.scala 335:62:@21708.4]
  reg [31:0] _RAND_111;
  reg [16:0] _T_1440; // @[Reg.scala 19:20:@21710.4]
  reg [31:0] _RAND_112;
  wire [16:0] _GEN_98; // @[Reg.scala 20:19:@21711.4]
  wire [18:0] _T_1442; // @[NV_NVDLA_CDMA_cvt.scala 342:47:@21714.4]
  wire [17:0] _T_1443; // @[NV_NVDLA_CDMA_cvt.scala 342:47:@21715.4]
  wire [17:0] _GEN_99; // @[NV_NVDLA_CDMA_cvt.scala 345:27:@21721.4]
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20811.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_1 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20814.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_1_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_1_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_1_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_1_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_1_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_2 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20817.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_2_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_2_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_2_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_2_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_2_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_3 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20820.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_3_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_3_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_3_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_3_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_3_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_4 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20823.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_4_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_4_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_4_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_4_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_4_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_5 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20826.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_5_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_5_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_5_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_5_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_5_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_6 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20829.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_6_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_6_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_6_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_6_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_6_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_7 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20832.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_7_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_7_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_7_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_7_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_7_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_8 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20835.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_8_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_8_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_8_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_8_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_8_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_9 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20838.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_9_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_9_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_9_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_9_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_9_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_10 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20841.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_10_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_10_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_10_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_10_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_10_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_11 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20844.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_11_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_11_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_11_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_11_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_11_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_12 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20847.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_12_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_12_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_12_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_12_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_12_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_13 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20850.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_13_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_13_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_13_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_13_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_13_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_14 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20853.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_14_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_14_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_14_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_14_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_14_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_15 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20856.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_15_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_15_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_15_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_15_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_15_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_16 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20859.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_16_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_16_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_16_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_16_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_16_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_17 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20862.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_17_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_17_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_17_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_17_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_17_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_18 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20865.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_18_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_18_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_18_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_18_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_18_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_19 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20868.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_19_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_19_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_19_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_19_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_19_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_20 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20871.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_20_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_20_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_20_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_20_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_20_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_21 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20874.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_21_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_21_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_21_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_21_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_21_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_22 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20877.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_22_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_22_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_22_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_22_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_22_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_23 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20880.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_23_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_23_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_23_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_23_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_23_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_24 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20883.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_24_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_24_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_24_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_24_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_24_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_25 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20886.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_25_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_25_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_25_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_25_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_25_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_26 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20889.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_26_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_26_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_26_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_26_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_26_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_27 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20892.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_27_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_27_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_27_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_27_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_27_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_28 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20895.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_28_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_28_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_28_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_28_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_28_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_29 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20898.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_29_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_29_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_29_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_29_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_29_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_30 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20901.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_30_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_30_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_30_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_30_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_30_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_out_rsc_bits)
  );
  NV_NVDLA_CDMA_CVT_cell NV_NVDLA_CDMA_CVT_cell_31 ( // @[NV_NVDLA_CDMA_cvt.scala 236:42:@20904.4]
    .reset(NV_NVDLA_CDMA_CVT_cell_31_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_CVT_cell_31_io_nvdla_core_clk),
    .io_cfg_mul_in_rsc(NV_NVDLA_CDMA_CVT_cell_31_io_cfg_mul_in_rsc),
    .io_cfg_out_precision(NV_NVDLA_CDMA_CVT_cell_31_io_cfg_out_precision),
    .io_cfg_truncate(NV_NVDLA_CDMA_CVT_cell_31_io_cfg_truncate),
    .io_chn_alu_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_valid),
    .io_chn_alu_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_bits),
    .io_chn_data_in_rsc_valid(NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_valid),
    .io_chn_data_in_rsc_bits(NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_bits),
    .io_chn_data_out_rsc_bits(NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_out_rsc_bits)
  );
  assign _T_126 = ~ io_dp2reg_done; // @[NV_NVDLA_CDMA_cvt.scala 91:15:@20110.4]
  assign _T_127 = _T_126 & io_reg2dp_op_en; // @[NV_NVDLA_CDMA_cvt.scala 91:31:@20111.4]
  assign _T_128 = ~ _T_89; // @[NV_NVDLA_CDMA_cvt.scala 92:28:@20112.4]
  assign _T_129 = _T_127 & _T_128; // @[NV_NVDLA_CDMA_cvt.scala 92:26:@20113.4]
  assign _T_140 = io_reg2dp_cvt_en ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12:@20125.6]
  assign _GEN_0 = _T_129 ? io_reg2dp_proc_precision : _T_92; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _GEN_1 = _T_129 ? io_reg2dp_cvt_scale : _T_95; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _GEN_2 = _T_129 ? io_reg2dp_cvt_truncate : _T_98; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _GEN_3 = _T_129 ? io_reg2dp_cvt_offset : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _GEN_4 = _T_129 ? _T_140 : _T_104; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _GEN_7 = _T_129 ? io_reg2dp_pad_value : _T_113; // @[NV_NVDLA_CDMA_cvt.scala 102:17:@20119.4]
  assign _T_153 = io_dc2cvt_dat_wr_addr_valid ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12:@20150.4]
  assign _T_154 = _T_153 & io_dc2cvt_dat_wr_info_pd; // @[NV_NVDLA_CDMA_cvt.scala 127:61:@20151.4]
  assign _T_158 = io_img2cvt_dat_wr_addr_valid ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12:@20153.4]
  assign _T_159 = _T_158 & io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_CDMA_cvt.scala 128:62:@20154.4]
  assign _T_160 = _T_154 | _T_159; // @[NV_NVDLA_CDMA_cvt.scala 127:88:@20155.4]
  assign _T_161 = _T_160[3:0]; // @[NV_NVDLA_CDMA_cvt.scala 130:33:@20156.4]
  assign _T_162 = _T_160[7]; // @[NV_NVDLA_CDMA_cvt.scala 131:33:@20157.4]
  assign _T_163 = _T_160[8]; // @[NV_NVDLA_CDMA_cvt.scala 132:33:@20158.4]
  assign _T_165 = io_dc2cvt_dat_wr_addr_valid | io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_CDMA_cvt.scala 135:46:@20160.4]
  assign _T_167 = io_img2cvt_dat_wr_addr_valid ? io_img2cvt_dat_wr_sel : 1'h0; // @[NV_NVDLA_CDMA_cvt.scala 138:27:@20161.4]
  assign _T_168 = io_dc2cvt_dat_wr_addr_valid ? io_dc2cvt_dat_wr_sel : _T_167; // @[NV_NVDLA_CDMA_cvt.scala 137:27:@20162.4]
  assign _T_170 = io_img2cvt_dat_wr_addr_valid ? io_img2cvt_dat_wr_pad_mask : 32'h0; // @[NV_NVDLA_CDMA_cvt.scala 140:26:@20163.4]
  assign _T_174 = io_dc2cvt_dat_wr_addr_valid ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12:@20165.4]
  assign _T_175 = _T_174 & io_dc2cvt_dat_wr_addr_bits; // @[NV_NVDLA_CDMA_cvt.scala 141:57:@20166.4]
  assign _T_179 = io_img2cvt_dat_wr_addr_valid ? 17'h1ffff : 17'h0; // @[Bitwise.scala 72:12:@20168.4]
  assign _T_180 = _T_179 & io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_CDMA_cvt.scala 142:58:@20169.4]
  assign _T_181 = _T_175 | _T_180; // @[NV_NVDLA_CDMA_cvt.scala 141:86:@20170.4]
  assign _T_185 = io_dc2cvt_dat_wr_addr_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@20172.4]
  assign _T_186 = _T_185 & io_dc2cvt_dat_wr_data; // @[NV_NVDLA_CDMA_cvt.scala 143:79:@20173.4]
  assign _T_190 = io_img2cvt_dat_wr_addr_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@20175.4]
  assign _T_191 = _T_190 & io_img2cvt_dat_wr_data; // @[NV_NVDLA_CDMA_cvt.scala 144:80:@20176.4]
  assign _T_192 = _T_186 | _T_191; // @[NV_NVDLA_CDMA_cvt.scala 143:103:@20177.4]
  assign _T_195 = _T_104[0]; // @[NV_NVDLA_CDMA_cvt.scala 155:45:@20179.4]
  assign _T_196 = _T_165 & _T_195; // @[NV_NVDLA_CDMA_cvt.scala 155:33:@20180.4]
  assign _T_197 = _T_161[0]; // @[NV_NVDLA_CDMA_cvt.scala 155:98:@20181.4]
  assign _T_201 = _T_197 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@20183.4]
  assign _T_203 = _T_196 ? _T_201 : 32'h0; // @[NV_NVDLA_CDMA_cvt.scala 155:22:@20184.4]
  assign _GEN_15 = _T_162 ? io_img2cvt_mn_wr_data : _T_214; // @[NV_NVDLA_CDMA_cvt.scala 184:22:@20204.6]
  assign _GEN_16 = _T_165 ? _T_162 : _T_209; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  assign _GEN_17 = _T_165 ? _T_163 : _T_212; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  assign _GEN_18 = _T_165 ? _T_181 : _T_228; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  assign _GEN_19 = _T_165 ? _T_161 : _T_231; // @[NV_NVDLA_CDMA_cvt.scala 179:16:@20199.4]
  assign _T_241 = _T_165 | _T_206; // @[NV_NVDLA_CDMA_cvt.scala 189:16:@20209.4]
  assign _GEN_22 = _T_241 ? _T_203 : _T_219; // @[NV_NVDLA_CDMA_cvt.scala 189:31:@20210.4]
  assign _GEN_23 = io_img2cvt_dat_wr_addr_valid ? _T_170 : _T_234; // @[NV_NVDLA_CDMA_cvt.scala 194:35:@20215.4]
  assign _GEN_24 = _T_165 ? {{1'd0}, _T_168} : _T_237; // @[NV_NVDLA_CDMA_cvt.scala 198:20:@20218.4]
  assign _T_432 = _T_216[7]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20227.4]
  assign _T_433 = ~ _T_212; // @[NV_NVDLA_CDMA_cvt.scala 214:69:@20228.4]
  assign _T_434 = _T_432 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20229.4]
  assign _T_438 = _T_434 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20232.4]
  assign _T_439 = _T_216[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20233.4]
  assign _T_440 = {_T_438,_T_439}; // @[Cat.scala 30:58:@20234.4]
  assign _T_441 = _T_214[15:0]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20236.4]
  assign _T_443 = _T_209 ? _T_441 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20238.4]
  assign _T_444 = _T_219[0]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20240.4]
  assign _T_445 = _T_216[15]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20245.4]
  assign _T_447 = _T_445 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20247.4]
  assign _T_451 = _T_447 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20250.4]
  assign _T_452 = _T_216[15:8]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20251.4]
  assign _T_453 = {_T_451,_T_452}; // @[Cat.scala 30:58:@20252.4]
  assign _T_454 = _T_214[31:16]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20254.4]
  assign _T_456 = _T_209 ? _T_454 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20256.4]
  assign _T_457 = _T_219[1]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20258.4]
  assign _T_458 = _T_216[23]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20263.4]
  assign _T_460 = _T_458 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20265.4]
  assign _T_464 = _T_460 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20268.4]
  assign _T_465 = _T_216[23:16]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20269.4]
  assign _T_466 = {_T_464,_T_465}; // @[Cat.scala 30:58:@20270.4]
  assign _T_467 = _T_214[47:32]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20272.4]
  assign _T_469 = _T_209 ? _T_467 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20274.4]
  assign _T_470 = _T_219[2]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20276.4]
  assign _T_471 = _T_216[31]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20281.4]
  assign _T_473 = _T_471 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20283.4]
  assign _T_477 = _T_473 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20286.4]
  assign _T_478 = _T_216[31:24]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20287.4]
  assign _T_479 = {_T_477,_T_478}; // @[Cat.scala 30:58:@20288.4]
  assign _T_480 = _T_214[63:48]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20290.4]
  assign _T_482 = _T_209 ? _T_480 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20292.4]
  assign _T_483 = _T_219[3]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20294.4]
  assign _T_484 = _T_216[39]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20299.4]
  assign _T_486 = _T_484 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20301.4]
  assign _T_490 = _T_486 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20304.4]
  assign _T_491 = _T_216[39:32]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20305.4]
  assign _T_492 = {_T_490,_T_491}; // @[Cat.scala 30:58:@20306.4]
  assign _T_493 = _T_214[79:64]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20308.4]
  assign _T_495 = _T_209 ? _T_493 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20310.4]
  assign _T_496 = _T_219[4]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20312.4]
  assign _T_497 = _T_216[47]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20317.4]
  assign _T_499 = _T_497 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20319.4]
  assign _T_503 = _T_499 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20322.4]
  assign _T_504 = _T_216[47:40]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20323.4]
  assign _T_505 = {_T_503,_T_504}; // @[Cat.scala 30:58:@20324.4]
  assign _T_506 = _T_214[95:80]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20326.4]
  assign _T_508 = _T_209 ? _T_506 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20328.4]
  assign _T_509 = _T_219[5]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20330.4]
  assign _T_510 = _T_216[55]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20335.4]
  assign _T_512 = _T_510 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20337.4]
  assign _T_516 = _T_512 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20340.4]
  assign _T_517 = _T_216[55:48]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20341.4]
  assign _T_518 = {_T_516,_T_517}; // @[Cat.scala 30:58:@20342.4]
  assign _T_519 = _T_214[111:96]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20344.4]
  assign _T_521 = _T_209 ? _T_519 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20346.4]
  assign _T_522 = _T_219[6]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20348.4]
  assign _T_523 = _T_216[63]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20353.4]
  assign _T_525 = _T_523 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20355.4]
  assign _T_529 = _T_525 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20358.4]
  assign _T_530 = _T_216[63:56]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20359.4]
  assign _T_531 = {_T_529,_T_530}; // @[Cat.scala 30:58:@20360.4]
  assign _T_532 = _T_214[127:112]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20362.4]
  assign _T_534 = _T_209 ? _T_532 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20364.4]
  assign _T_535 = _T_219[7]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20366.4]
  assign _T_536 = _T_216[71]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20371.4]
  assign _T_538 = _T_536 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20373.4]
  assign _T_542 = _T_538 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20376.4]
  assign _T_543 = _T_216[71:64]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20377.4]
  assign _T_544 = {_T_542,_T_543}; // @[Cat.scala 30:58:@20378.4]
  assign _T_545 = _T_214[143:128]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20380.4]
  assign _T_547 = _T_209 ? _T_545 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20382.4]
  assign _T_548 = _T_219[8]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20384.4]
  assign _T_549 = _T_216[79]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20389.4]
  assign _T_551 = _T_549 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20391.4]
  assign _T_555 = _T_551 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20394.4]
  assign _T_556 = _T_216[79:72]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20395.4]
  assign _T_557 = {_T_555,_T_556}; // @[Cat.scala 30:58:@20396.4]
  assign _T_558 = _T_214[159:144]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20398.4]
  assign _T_560 = _T_209 ? _T_558 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20400.4]
  assign _T_561 = _T_219[9]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20402.4]
  assign _T_562 = _T_216[87]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20407.4]
  assign _T_564 = _T_562 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20409.4]
  assign _T_568 = _T_564 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20412.4]
  assign _T_569 = _T_216[87:80]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20413.4]
  assign _T_570 = {_T_568,_T_569}; // @[Cat.scala 30:58:@20414.4]
  assign _T_571 = _T_214[175:160]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20416.4]
  assign _T_573 = _T_209 ? _T_571 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20418.4]
  assign _T_574 = _T_219[10]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20420.4]
  assign _T_575 = _T_216[95]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20425.4]
  assign _T_577 = _T_575 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20427.4]
  assign _T_581 = _T_577 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20430.4]
  assign _T_582 = _T_216[95:88]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20431.4]
  assign _T_583 = {_T_581,_T_582}; // @[Cat.scala 30:58:@20432.4]
  assign _T_584 = _T_214[191:176]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20434.4]
  assign _T_586 = _T_209 ? _T_584 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20436.4]
  assign _T_587 = _T_219[11]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20438.4]
  assign _T_588 = _T_216[103]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20443.4]
  assign _T_590 = _T_588 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20445.4]
  assign _T_594 = _T_590 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20448.4]
  assign _T_595 = _T_216[103:96]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20449.4]
  assign _T_596 = {_T_594,_T_595}; // @[Cat.scala 30:58:@20450.4]
  assign _T_597 = _T_214[207:192]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20452.4]
  assign _T_599 = _T_209 ? _T_597 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20454.4]
  assign _T_600 = _T_219[12]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20456.4]
  assign _T_601 = _T_216[111]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20461.4]
  assign _T_603 = _T_601 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20463.4]
  assign _T_607 = _T_603 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20466.4]
  assign _T_608 = _T_216[111:104]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20467.4]
  assign _T_609 = {_T_607,_T_608}; // @[Cat.scala 30:58:@20468.4]
  assign _T_610 = _T_214[223:208]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20470.4]
  assign _T_612 = _T_209 ? _T_610 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20472.4]
  assign _T_613 = _T_219[13]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20474.4]
  assign _T_614 = _T_216[119]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20479.4]
  assign _T_616 = _T_614 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20481.4]
  assign _T_620 = _T_616 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20484.4]
  assign _T_621 = _T_216[119:112]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20485.4]
  assign _T_622 = {_T_620,_T_621}; // @[Cat.scala 30:58:@20486.4]
  assign _T_623 = _T_214[239:224]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20488.4]
  assign _T_625 = _T_209 ? _T_623 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20490.4]
  assign _T_626 = _T_219[14]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20492.4]
  assign _T_627 = _T_216[127]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20497.4]
  assign _T_629 = _T_627 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20499.4]
  assign _T_633 = _T_629 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20502.4]
  assign _T_634 = _T_216[127:120]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20503.4]
  assign _T_635 = {_T_633,_T_634}; // @[Cat.scala 30:58:@20504.4]
  assign _T_636 = _T_214[255:240]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20506.4]
  assign _T_638 = _T_209 ? _T_636 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20508.4]
  assign _T_639 = _T_219[15]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20510.4]
  assign _T_640 = _T_216[135]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20515.4]
  assign _T_642 = _T_640 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20517.4]
  assign _T_646 = _T_642 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20520.4]
  assign _T_647 = _T_216[135:128]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20521.4]
  assign _T_648 = {_T_646,_T_647}; // @[Cat.scala 30:58:@20522.4]
  assign _T_649 = _T_214[271:256]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20524.4]
  assign _T_651 = _T_209 ? _T_649 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20526.4]
  assign _T_652 = _T_219[16]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20528.4]
  assign _T_653 = _T_216[143]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20533.4]
  assign _T_655 = _T_653 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20535.4]
  assign _T_659 = _T_655 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20538.4]
  assign _T_660 = _T_216[143:136]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20539.4]
  assign _T_661 = {_T_659,_T_660}; // @[Cat.scala 30:58:@20540.4]
  assign _T_662 = _T_214[287:272]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20542.4]
  assign _T_664 = _T_209 ? _T_662 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20544.4]
  assign _T_665 = _T_219[17]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20546.4]
  assign _T_666 = _T_216[151]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20551.4]
  assign _T_668 = _T_666 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20553.4]
  assign _T_672 = _T_668 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20556.4]
  assign _T_673 = _T_216[151:144]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20557.4]
  assign _T_674 = {_T_672,_T_673}; // @[Cat.scala 30:58:@20558.4]
  assign _T_675 = _T_214[303:288]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20560.4]
  assign _T_677 = _T_209 ? _T_675 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20562.4]
  assign _T_678 = _T_219[18]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20564.4]
  assign _T_679 = _T_216[159]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20569.4]
  assign _T_681 = _T_679 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20571.4]
  assign _T_685 = _T_681 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20574.4]
  assign _T_686 = _T_216[159:152]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20575.4]
  assign _T_687 = {_T_685,_T_686}; // @[Cat.scala 30:58:@20576.4]
  assign _T_688 = _T_214[319:304]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20578.4]
  assign _T_690 = _T_209 ? _T_688 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20580.4]
  assign _T_691 = _T_219[19]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20582.4]
  assign _T_692 = _T_216[167]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20587.4]
  assign _T_694 = _T_692 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20589.4]
  assign _T_698 = _T_694 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20592.4]
  assign _T_699 = _T_216[167:160]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20593.4]
  assign _T_700 = {_T_698,_T_699}; // @[Cat.scala 30:58:@20594.4]
  assign _T_701 = _T_214[335:320]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20596.4]
  assign _T_703 = _T_209 ? _T_701 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20598.4]
  assign _T_704 = _T_219[20]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20600.4]
  assign _T_705 = _T_216[175]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20605.4]
  assign _T_707 = _T_705 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20607.4]
  assign _T_711 = _T_707 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20610.4]
  assign _T_712 = _T_216[175:168]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20611.4]
  assign _T_713 = {_T_711,_T_712}; // @[Cat.scala 30:58:@20612.4]
  assign _T_714 = _T_214[351:336]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20614.4]
  assign _T_716 = _T_209 ? _T_714 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20616.4]
  assign _T_717 = _T_219[21]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20618.4]
  assign _T_718 = _T_216[183]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20623.4]
  assign _T_720 = _T_718 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20625.4]
  assign _T_724 = _T_720 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20628.4]
  assign _T_725 = _T_216[183:176]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20629.4]
  assign _T_726 = {_T_724,_T_725}; // @[Cat.scala 30:58:@20630.4]
  assign _T_727 = _T_214[367:352]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20632.4]
  assign _T_729 = _T_209 ? _T_727 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20634.4]
  assign _T_730 = _T_219[22]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20636.4]
  assign _T_731 = _T_216[191]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20641.4]
  assign _T_733 = _T_731 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20643.4]
  assign _T_737 = _T_733 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20646.4]
  assign _T_738 = _T_216[191:184]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20647.4]
  assign _T_739 = {_T_737,_T_738}; // @[Cat.scala 30:58:@20648.4]
  assign _T_740 = _T_214[383:368]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20650.4]
  assign _T_742 = _T_209 ? _T_740 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20652.4]
  assign _T_743 = _T_219[23]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20654.4]
  assign _T_744 = _T_216[199]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20659.4]
  assign _T_746 = _T_744 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20661.4]
  assign _T_750 = _T_746 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20664.4]
  assign _T_751 = _T_216[199:192]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20665.4]
  assign _T_752 = {_T_750,_T_751}; // @[Cat.scala 30:58:@20666.4]
  assign _T_753 = _T_214[399:384]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20668.4]
  assign _T_755 = _T_209 ? _T_753 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20670.4]
  assign _T_756 = _T_219[24]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20672.4]
  assign _T_757 = _T_216[207]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20677.4]
  assign _T_759 = _T_757 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20679.4]
  assign _T_763 = _T_759 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20682.4]
  assign _T_764 = _T_216[207:200]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20683.4]
  assign _T_765 = {_T_763,_T_764}; // @[Cat.scala 30:58:@20684.4]
  assign _T_766 = _T_214[415:400]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20686.4]
  assign _T_768 = _T_209 ? _T_766 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20688.4]
  assign _T_769 = _T_219[25]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20690.4]
  assign _T_770 = _T_216[215]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20695.4]
  assign _T_772 = _T_770 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20697.4]
  assign _T_776 = _T_772 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20700.4]
  assign _T_777 = _T_216[215:208]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20701.4]
  assign _T_778 = {_T_776,_T_777}; // @[Cat.scala 30:58:@20702.4]
  assign _T_779 = _T_214[431:416]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20704.4]
  assign _T_781 = _T_209 ? _T_779 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20706.4]
  assign _T_782 = _T_219[26]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20708.4]
  assign _T_783 = _T_216[223]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20713.4]
  assign _T_785 = _T_783 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20715.4]
  assign _T_789 = _T_785 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20718.4]
  assign _T_790 = _T_216[223:216]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20719.4]
  assign _T_791 = {_T_789,_T_790}; // @[Cat.scala 30:58:@20720.4]
  assign _T_792 = _T_214[447:432]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20722.4]
  assign _T_794 = _T_209 ? _T_792 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20724.4]
  assign _T_795 = _T_219[27]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20726.4]
  assign _T_796 = _T_216[231]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20731.4]
  assign _T_798 = _T_796 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20733.4]
  assign _T_802 = _T_798 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20736.4]
  assign _T_803 = _T_216[231:224]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20737.4]
  assign _T_804 = {_T_802,_T_803}; // @[Cat.scala 30:58:@20738.4]
  assign _T_805 = _T_214[463:448]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20740.4]
  assign _T_807 = _T_209 ? _T_805 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20742.4]
  assign _T_808 = _T_219[28]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20744.4]
  assign _T_809 = _T_216[239]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20749.4]
  assign _T_811 = _T_809 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20751.4]
  assign _T_815 = _T_811 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20754.4]
  assign _T_816 = _T_216[239:232]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20755.4]
  assign _T_817 = {_T_815,_T_816}; // @[Cat.scala 30:58:@20756.4]
  assign _T_818 = _T_214[479:464]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20758.4]
  assign _T_820 = _T_209 ? _T_818 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20760.4]
  assign _T_821 = _T_219[29]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20762.4]
  assign _T_822 = _T_216[247]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20767.4]
  assign _T_824 = _T_822 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20769.4]
  assign _T_828 = _T_824 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20772.4]
  assign _T_829 = _T_216[247:240]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20773.4]
  assign _T_830 = {_T_828,_T_829}; // @[Cat.scala 30:58:@20774.4]
  assign _T_831 = _T_214[495:480]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20776.4]
  assign _T_833 = _T_209 ? _T_831 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20778.4]
  assign _T_834 = _T_219[30]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20780.4]
  assign _T_835 = _T_216[255]; // @[NV_NVDLA_CDMA_cvt.scala 214:42:@20785.4]
  assign _T_837 = _T_835 & _T_433; // @[NV_NVDLA_CDMA_cvt.scala 214:67:@20787.4]
  assign _T_841 = _T_837 ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12:@20790.4]
  assign _T_842 = _T_216[255:248]; // @[NV_NVDLA_CDMA_cvt.scala 215:90:@20791.4]
  assign _T_843 = {_T_841,_T_842}; // @[Cat.scala 30:58:@20792.4]
  assign _T_844 = _T_214[511:496]; // @[NV_NVDLA_CDMA_cvt.scala 216:63:@20794.4]
  assign _T_846 = _T_209 ? _T_844 : _T_101; // @[NV_NVDLA_CDMA_cvt.scala 216:27:@20796.4]
  assign _T_847 = _T_219[31]; // @[NV_NVDLA_CDMA_cvt.scala 217:24:@20798.4]
  assign _T_854 = _T_206 | _T_850; // @[NV_NVDLA_CDMA_cvt.scala 227:19:@20806.4]
  assign _GEN_89 = _T_854 ? _T_219 : _T_853; // @[NV_NVDLA_CDMA_cvt.scala 227:30:@20807.4]
  assign _T_858_0 = NV_NVDLA_CDMA_CVT_cell_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20918.4]
  assign _T_989 = _T_858_0[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21291.4]
  assign _T_858_1 = NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20930.4]
  assign _T_990 = _T_858_1[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21292.4]
  assign _T_858_2 = NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20942.4]
  assign _T_991 = _T_858_2[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21293.4]
  assign _T_858_3 = NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20954.4]
  assign _T_992 = _T_858_3[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21294.4]
  assign _T_858_4 = NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20966.4]
  assign _T_993 = _T_858_4[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21295.4]
  assign _T_858_5 = NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20978.4]
  assign _T_994 = _T_858_5[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21296.4]
  assign _T_858_6 = NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@20990.4]
  assign _T_995 = _T_858_6[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21297.4]
  assign _T_858_7 = NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21002.4]
  assign _T_996 = _T_858_7[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21298.4]
  assign _T_858_8 = NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21014.4]
  assign _T_997 = _T_858_8[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21299.4]
  assign _T_858_9 = NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21026.4]
  assign _T_998 = _T_858_9[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21300.4]
  assign _T_858_10 = NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21038.4]
  assign _T_999 = _T_858_10[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21301.4]
  assign _T_858_11 = NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21050.4]
  assign _T_1000 = _T_858_11[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21302.4]
  assign _T_858_12 = NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21062.4]
  assign _T_1001 = _T_858_12[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21303.4]
  assign _T_858_13 = NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21074.4]
  assign _T_1002 = _T_858_13[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21304.4]
  assign _T_858_14 = NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21086.4]
  assign _T_1003 = _T_858_14[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21305.4]
  assign _T_858_15 = NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21098.4]
  assign _T_1004 = _T_858_15[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21306.4]
  assign _T_858_16 = NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21110.4]
  assign _T_1005 = _T_858_16[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21307.4]
  assign _T_858_17 = NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21122.4]
  assign _T_1006 = _T_858_17[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21308.4]
  assign _T_858_18 = NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21134.4]
  assign _T_1007 = _T_858_18[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21309.4]
  assign _T_858_19 = NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21146.4]
  assign _T_1008 = _T_858_19[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21310.4]
  assign _T_858_20 = NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21158.4]
  assign _T_1009 = _T_858_20[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21311.4]
  assign _T_858_21 = NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21170.4]
  assign _T_1010 = _T_858_21[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21312.4]
  assign _T_858_22 = NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21182.4]
  assign _T_1011 = _T_858_22[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21313.4]
  assign _T_858_23 = NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21194.4]
  assign _T_1012 = _T_858_23[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21314.4]
  assign _T_858_24 = NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21206.4]
  assign _T_1013 = _T_858_24[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21315.4]
  assign _T_858_25 = NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21218.4]
  assign _T_1014 = _T_858_25[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21316.4]
  assign _T_858_26 = NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21230.4]
  assign _T_1015 = _T_858_26[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21317.4]
  assign _T_858_27 = NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21242.4]
  assign _T_1016 = _T_858_27[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21318.4]
  assign _T_858_28 = NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21254.4]
  assign _T_1017 = _T_858_28[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21319.4]
  assign _T_858_29 = NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21266.4]
  assign _T_1018 = _T_858_29[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21320.4]
  assign _T_858_30 = NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21278.4]
  assign _T_1019 = _T_858_30[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21321.4]
  assign _T_858_31 = NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_out_rsc_bits; // @[NV_NVDLA_CDMA_cvt.scala 234:19:@20810.4 NV_NVDLA_CDMA_cvt.scala 251:16:@21290.4]
  assign _T_1020 = _T_858_31[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 254:69:@21322.4]
  assign _T_1065 = {_T_996,_T_995,_T_994,_T_993,_T_992,_T_991,_T_990,_T_989}; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21362.4]
  assign _T_1073 = {_T_1004,_T_1003,_T_1002,_T_1001,_T_1000,_T_999,_T_998,_T_997,_T_1065}; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21370.4]
  assign _T_1080 = {_T_1012,_T_1011,_T_1010,_T_1009,_T_1008,_T_1007,_T_1006,_T_1005}; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21377.4]
  assign _T_1089 = {_T_1020,_T_1019,_T_1018,_T_1017,_T_1016,_T_1015,_T_1014,_T_1013,_T_1080,_T_1073}; // @[NV_NVDLA_CDMA_cvt.scala 254:93:@21386.4]
  assign _T_1119 = _T_237[0]; // @[NV_NVDLA_CDMA_cvt.scala 264:61:@21397.4 NV_NVDLA_CDMA_cvt.scala 279:29:@21424.4]
  assign _GEN_90 = _T_222 ? _T_1119 : _T_1122; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21431.4]
  assign _GEN_92 = _T_1094 ? _T_1122 : _T_1125; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21443.4]
  assign _GEN_94 = _T_1097 ? _T_1125 : _T_1128; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21455.4]
  assign _GEN_96 = _T_1100 ? _T_1128 : _T_1131; // @[NV_NVDLA_CDMA_cvt.scala 290:34:@21467.4]
  assign _T_1192 = _T_104[1]; // @[NV_NVDLA_CDMA_cvt.scala 303:41:@21477.4]
  assign _T_1193 = _T_1192 ? {{1'd0}, _T_1131} : _T_237; // @[NV_NVDLA_CDMA_cvt.scala 303:30:@21478.4]
  assign _T_1195 = _T_1192 ? _T_1117 : _T_222; // @[NV_NVDLA_CDMA_cvt.scala 305:25:@21480.4]
  assign _T_1197 = _T_1192 ? _T_1159 : _T_228; // @[NV_NVDLA_CDMA_cvt.scala 306:26:@21482.4]
  assign _T_1198 = _T_104[2]; // @[NV_NVDLA_CDMA_cvt.scala 307:40:@21483.4]
  assign _T_1199 = _T_1198 ? _T_1173 : _T_231; // @[NV_NVDLA_CDMA_cvt.scala 307:29:@21484.4]
  assign _T_1200 = _T_104[3]; // @[NV_NVDLA_CDMA_cvt.scala 308:40:@21485.4]
  assign _T_1201 = _T_1200 ? _T_1117 : _T_225; // @[NV_NVDLA_CDMA_cvt.scala 308:29:@21486.4]
  assign _T_1202 = ~ _T_1201; // @[NV_NVDLA_CDMA_cvt.scala 309:31:@21487.4]
  assign _T_1205 = _T_1200 ? _T_1187 : _T_234; // @[NV_NVDLA_CDMA_cvt.scala 310:30:@21489.4]
  assign _T_1206 = _T_1202 ? 32'h0 : _T_1205; // @[NV_NVDLA_CDMA_cvt.scala 309:30:@21490.4]
  assign _T_1214 = _T_104[5]; // @[NV_NVDLA_CDMA_cvt.scala 320:38:@21495.4]
  assign _T_1215 = _T_1214 ? _T_1089 : _T_216; // @[NV_NVDLA_CDMA_cvt.scala 320:27:@21496.4]
  assign _T_1216 = _T_1206[0]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21497.4]
  assign _T_1217 = _T_113[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 322:49:@21498.4]
  assign _T_1218 = _T_1215[7:0]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21499.4]
  assign _T_1219 = _T_1216 ? _T_1217 : _T_1218; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21500.4]
  assign _T_1220 = _T_1206[1]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21501.4]
  assign _T_1222 = _T_1215[15:8]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21503.4]
  assign _T_1223 = _T_1220 ? _T_1217 : _T_1222; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21504.4]
  assign _T_1224 = _T_1206[2]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21505.4]
  assign _T_1226 = _T_1215[23:16]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21507.4]
  assign _T_1227 = _T_1224 ? _T_1217 : _T_1226; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21508.4]
  assign _T_1228 = _T_1206[3]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21509.4]
  assign _T_1230 = _T_1215[31:24]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21511.4]
  assign _T_1231 = _T_1228 ? _T_1217 : _T_1230; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21512.4]
  assign _T_1232 = _T_1206[4]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21513.4]
  assign _T_1234 = _T_1215[39:32]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21515.4]
  assign _T_1235 = _T_1232 ? _T_1217 : _T_1234; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21516.4]
  assign _T_1236 = _T_1206[5]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21517.4]
  assign _T_1238 = _T_1215[47:40]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21519.4]
  assign _T_1239 = _T_1236 ? _T_1217 : _T_1238; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21520.4]
  assign _T_1240 = _T_1206[6]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21521.4]
  assign _T_1242 = _T_1215[55:48]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21523.4]
  assign _T_1243 = _T_1240 ? _T_1217 : _T_1242; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21524.4]
  assign _T_1244 = _T_1206[7]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21525.4]
  assign _T_1246 = _T_1215[63:56]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21527.4]
  assign _T_1247 = _T_1244 ? _T_1217 : _T_1246; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21528.4]
  assign _T_1248 = _T_1206[8]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21529.4]
  assign _T_1250 = _T_1215[71:64]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21531.4]
  assign _T_1251 = _T_1248 ? _T_1217 : _T_1250; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21532.4]
  assign _T_1252 = _T_1206[9]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21533.4]
  assign _T_1254 = _T_1215[79:72]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21535.4]
  assign _T_1255 = _T_1252 ? _T_1217 : _T_1254; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21536.4]
  assign _T_1256 = _T_1206[10]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21537.4]
  assign _T_1258 = _T_1215[87:80]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21539.4]
  assign _T_1259 = _T_1256 ? _T_1217 : _T_1258; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21540.4]
  assign _T_1260 = _T_1206[11]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21541.4]
  assign _T_1262 = _T_1215[95:88]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21543.4]
  assign _T_1263 = _T_1260 ? _T_1217 : _T_1262; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21544.4]
  assign _T_1264 = _T_1206[12]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21545.4]
  assign _T_1266 = _T_1215[103:96]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21547.4]
  assign _T_1267 = _T_1264 ? _T_1217 : _T_1266; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21548.4]
  assign _T_1268 = _T_1206[13]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21549.4]
  assign _T_1270 = _T_1215[111:104]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21551.4]
  assign _T_1271 = _T_1268 ? _T_1217 : _T_1270; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21552.4]
  assign _T_1272 = _T_1206[14]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21553.4]
  assign _T_1274 = _T_1215[119:112]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21555.4]
  assign _T_1275 = _T_1272 ? _T_1217 : _T_1274; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21556.4]
  assign _T_1276 = _T_1206[15]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21557.4]
  assign _T_1278 = _T_1215[127:120]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21559.4]
  assign _T_1279 = _T_1276 ? _T_1217 : _T_1278; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21560.4]
  assign _T_1280 = _T_1206[16]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21561.4]
  assign _T_1282 = _T_1215[135:128]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21563.4]
  assign _T_1283 = _T_1280 ? _T_1217 : _T_1282; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21564.4]
  assign _T_1284 = _T_1206[17]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21565.4]
  assign _T_1286 = _T_1215[143:136]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21567.4]
  assign _T_1287 = _T_1284 ? _T_1217 : _T_1286; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21568.4]
  assign _T_1288 = _T_1206[18]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21569.4]
  assign _T_1290 = _T_1215[151:144]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21571.4]
  assign _T_1291 = _T_1288 ? _T_1217 : _T_1290; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21572.4]
  assign _T_1292 = _T_1206[19]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21573.4]
  assign _T_1294 = _T_1215[159:152]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21575.4]
  assign _T_1295 = _T_1292 ? _T_1217 : _T_1294; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21576.4]
  assign _T_1296 = _T_1206[20]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21577.4]
  assign _T_1298 = _T_1215[167:160]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21579.4]
  assign _T_1299 = _T_1296 ? _T_1217 : _T_1298; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21580.4]
  assign _T_1300 = _T_1206[21]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21581.4]
  assign _T_1302 = _T_1215[175:168]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21583.4]
  assign _T_1303 = _T_1300 ? _T_1217 : _T_1302; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21584.4]
  assign _T_1304 = _T_1206[22]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21585.4]
  assign _T_1306 = _T_1215[183:176]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21587.4]
  assign _T_1307 = _T_1304 ? _T_1217 : _T_1306; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21588.4]
  assign _T_1308 = _T_1206[23]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21589.4]
  assign _T_1310 = _T_1215[191:184]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21591.4]
  assign _T_1311 = _T_1308 ? _T_1217 : _T_1310; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21592.4]
  assign _T_1312 = _T_1206[24]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21593.4]
  assign _T_1314 = _T_1215[199:192]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21595.4]
  assign _T_1315 = _T_1312 ? _T_1217 : _T_1314; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21596.4]
  assign _T_1316 = _T_1206[25]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21597.4]
  assign _T_1318 = _T_1215[207:200]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21599.4]
  assign _T_1319 = _T_1316 ? _T_1217 : _T_1318; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21600.4]
  assign _T_1320 = _T_1206[26]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21601.4]
  assign _T_1322 = _T_1215[215:208]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21603.4]
  assign _T_1323 = _T_1320 ? _T_1217 : _T_1322; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21604.4]
  assign _T_1324 = _T_1206[27]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21605.4]
  assign _T_1326 = _T_1215[223:216]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21607.4]
  assign _T_1327 = _T_1324 ? _T_1217 : _T_1326; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21608.4]
  assign _T_1328 = _T_1206[28]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21609.4]
  assign _T_1330 = _T_1215[231:224]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21611.4]
  assign _T_1331 = _T_1328 ? _T_1217 : _T_1330; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21612.4]
  assign _T_1332 = _T_1206[29]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21613.4]
  assign _T_1334 = _T_1215[239:232]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21615.4]
  assign _T_1335 = _T_1332 ? _T_1217 : _T_1334; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21616.4]
  assign _T_1336 = _T_1206[30]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21617.4]
  assign _T_1338 = _T_1215[247:240]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21619.4]
  assign _T_1339 = _T_1336 ? _T_1217 : _T_1338; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21620.4]
  assign _T_1340 = _T_1206[31]; // @[NV_NVDLA_CDMA_cvt.scala 322:31:@21621.4]
  assign _T_1342 = _T_1215[255:248]; // @[NV_NVDLA_CDMA_cvt.scala 322:88:@21623.4]
  assign _T_1343 = _T_1340 ? _T_1217 : _T_1342; // @[NV_NVDLA_CDMA_cvt.scala 322:11:@21624.4]
  assign _T_1388 = {_T_1247,_T_1243,_T_1239,_T_1235,_T_1231,_T_1227,_T_1223,_T_1219}; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21664.4]
  assign _T_1396 = {_T_1279,_T_1275,_T_1271,_T_1267,_T_1263,_T_1259,_T_1255,_T_1251,_T_1388}; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21672.4]
  assign _T_1403 = {_T_1311,_T_1307,_T_1303,_T_1299,_T_1295,_T_1291,_T_1287,_T_1283}; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21679.4]
  assign _T_1412 = {_T_1343,_T_1339,_T_1335,_T_1331,_T_1327,_T_1323,_T_1319,_T_1315,_T_1403,_T_1396}; // @[NV_NVDLA_CDMA_cvt.scala 322:134:@21688.4]
  assign _T_1413 = _T_1199[0]; // @[NV_NVDLA_CDMA_cvt.scala 323:45:@21689.4]
  assign _T_1416 = _T_1413 ? _T_1412 : 256'h0; // @[NV_NVDLA_CDMA_cvt.scala 323:26:@21691.4]
  assign _T_1444 = _T_1213[13]; // @[NV_NVDLA_CDMA_cvt.scala 343:44:@21716.4]
  assign _T_1445 = ~ _T_1444; // @[NV_NVDLA_CDMA_cvt.scala 343:25:@21717.4]
  assign _T_1420 = _T_1195 | _T_1445; // @[NV_NVDLA_CDMA_cvt.scala 325:40:@21694.4]
  assign _T_1421 = _T_1213[17:1]; // @[NV_NVDLA_CDMA_cvt.scala 326:70:@21695.4]
  assign _T_1422 = _T_1445 ? _T_1421 : _T_1197; // @[NV_NVDLA_CDMA_cvt.scala 326:29:@21696.4]
  assign _T_1423 = _T_1213[0]; // @[NV_NVDLA_CDMA_cvt.scala 328:78:@21697.4]
  assign _T_1425 = ~ _T_1423; // @[NV_NVDLA_CDMA_cvt.scala 328:83:@21699.4]
  assign _T_1426 = {_T_1423,_T_1425}; // @[Cat.scala 30:58:@21700.4]
  assign _T_1427 = _T_1193[0]; // @[NV_NVDLA_CDMA_cvt.scala 329:47:@21701.4]
  assign _T_1429 = ~ _T_1427; // @[NV_NVDLA_CDMA_cvt.scala 329:52:@21703.4]
  assign _T_1430 = {_T_1427,_T_1429}; // @[Cat.scala 30:58:@21704.4]
  assign _T_1431 = _T_1445 ? _T_1426 : _T_1430; // @[NV_NVDLA_CDMA_cvt.scala 328:33:@21705.4]
  assign _GEN_98 = _T_1420 ? _T_1422 : _T_1440; // @[Reg.scala 20:19:@21711.4]
  assign _T_1442 = _T_1213 + 18'h1; // @[NV_NVDLA_CDMA_cvt.scala 342:47:@21714.4]
  assign _T_1443 = _T_1213 + 18'h1; // @[NV_NVDLA_CDMA_cvt.scala 342:47:@21715.4]
  assign _GEN_99 = _T_1445 ? _T_1443 : _T_1213; // @[NV_NVDLA_CDMA_cvt.scala 345:27:@21721.4]
  assign io_cdma2buf_dat_wr_sel = _T_1434; // @[NV_NVDLA_CDMA_cvt.scala 357:32:@21726.4]
  assign io_cdma2buf_dat_wr_addr_valid = _T_1437; // @[NV_NVDLA_CDMA_cvt.scala 354:31:@21724.4]
  assign io_cdma2buf_dat_wr_addr_bits = _T_1440; // @[NV_NVDLA_CDMA_cvt.scala 355:30:@21725.4]
  assign io_cdma2buf_dat_wr_data = _T_1419; // @[NV_NVDLA_CDMA_cvt.scala 359:25:@21727.4]
  assign io_dp2reg_dat_flush_done = _T_1213[13]; // @[NV_NVDLA_CDMA_cvt.scala 344:26:@21720.4]
  assign NV_NVDLA_CDMA_CVT_cell_reset = reset; // @[:@20813.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20907.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20914.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20915.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20916.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_valid = _T_853[0]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20913.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_chn_alu_in_rsc_bits = _T_283_0; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20911.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_valid = _T_853[0]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20910.4]
  assign NV_NVDLA_CDMA_CVT_cell_io_chn_data_in_rsc_bits = _T_245_0; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20908.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_reset = reset; // @[:@20816.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20919.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20926.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20927.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20928.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_valid = _T_853[1]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20925.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_chn_alu_in_rsc_bits = _T_283_1; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20923.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_valid = _T_853[1]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20922.4]
  assign NV_NVDLA_CDMA_CVT_cell_1_io_chn_data_in_rsc_bits = _T_245_1; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20920.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_reset = reset; // @[:@20819.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20931.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20938.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20939.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20940.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_valid = _T_853[2]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20937.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_chn_alu_in_rsc_bits = _T_283_2; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20935.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_valid = _T_853[2]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20934.4]
  assign NV_NVDLA_CDMA_CVT_cell_2_io_chn_data_in_rsc_bits = _T_245_2; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20932.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_reset = reset; // @[:@20822.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20943.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20950.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20951.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20952.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_valid = _T_853[3]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20949.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_chn_alu_in_rsc_bits = _T_283_3; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20947.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_valid = _T_853[3]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20946.4]
  assign NV_NVDLA_CDMA_CVT_cell_3_io_chn_data_in_rsc_bits = _T_245_3; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20944.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_reset = reset; // @[:@20825.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20955.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20962.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20963.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20964.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_valid = _T_853[4]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20961.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_chn_alu_in_rsc_bits = _T_283_4; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20959.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_valid = _T_853[4]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20958.4]
  assign NV_NVDLA_CDMA_CVT_cell_4_io_chn_data_in_rsc_bits = _T_245_4; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20956.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_reset = reset; // @[:@20828.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20967.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20974.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20975.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20976.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_valid = _T_853[5]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20973.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_chn_alu_in_rsc_bits = _T_283_5; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20971.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_valid = _T_853[5]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20970.4]
  assign NV_NVDLA_CDMA_CVT_cell_5_io_chn_data_in_rsc_bits = _T_245_5; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20968.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_reset = reset; // @[:@20831.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20979.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20986.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20987.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@20988.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_valid = _T_853[6]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20985.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_chn_alu_in_rsc_bits = _T_283_6; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20983.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_valid = _T_853[6]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20982.4]
  assign NV_NVDLA_CDMA_CVT_cell_6_io_chn_data_in_rsc_bits = _T_245_6; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20980.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_reset = reset; // @[:@20834.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@20991.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@20998.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@20999.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21000.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_valid = _T_853[7]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@20997.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_chn_alu_in_rsc_bits = _T_283_7; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@20995.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_valid = _T_853[7]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@20994.4]
  assign NV_NVDLA_CDMA_CVT_cell_7_io_chn_data_in_rsc_bits = _T_245_7; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@20992.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_reset = reset; // @[:@20837.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21003.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21010.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21011.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21012.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_valid = _T_853[8]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21009.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_chn_alu_in_rsc_bits = _T_283_8; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21007.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_valid = _T_853[8]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21006.4]
  assign NV_NVDLA_CDMA_CVT_cell_8_io_chn_data_in_rsc_bits = _T_245_8; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21004.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_reset = reset; // @[:@20840.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21015.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21022.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21023.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21024.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_valid = _T_853[9]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21021.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_chn_alu_in_rsc_bits = _T_283_9; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21019.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_valid = _T_853[9]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21018.4]
  assign NV_NVDLA_CDMA_CVT_cell_9_io_chn_data_in_rsc_bits = _T_245_9; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21016.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_reset = reset; // @[:@20843.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21027.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21034.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21035.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21036.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_valid = _T_853[10]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21033.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_chn_alu_in_rsc_bits = _T_283_10; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21031.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_valid = _T_853[10]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21030.4]
  assign NV_NVDLA_CDMA_CVT_cell_10_io_chn_data_in_rsc_bits = _T_245_10; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21028.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_reset = reset; // @[:@20846.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21039.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21046.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21047.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21048.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_valid = _T_853[11]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21045.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_chn_alu_in_rsc_bits = _T_283_11; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21043.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_valid = _T_853[11]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21042.4]
  assign NV_NVDLA_CDMA_CVT_cell_11_io_chn_data_in_rsc_bits = _T_245_11; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21040.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_reset = reset; // @[:@20849.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21051.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21058.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21059.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21060.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_valid = _T_853[12]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21057.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_chn_alu_in_rsc_bits = _T_283_12; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21055.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_valid = _T_853[12]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21054.4]
  assign NV_NVDLA_CDMA_CVT_cell_12_io_chn_data_in_rsc_bits = _T_245_12; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21052.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_reset = reset; // @[:@20852.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21063.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21070.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21071.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21072.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_valid = _T_853[13]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21069.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_chn_alu_in_rsc_bits = _T_283_13; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21067.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_valid = _T_853[13]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21066.4]
  assign NV_NVDLA_CDMA_CVT_cell_13_io_chn_data_in_rsc_bits = _T_245_13; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21064.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_reset = reset; // @[:@20855.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21075.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21082.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21083.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21084.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_valid = _T_853[14]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21081.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_chn_alu_in_rsc_bits = _T_283_14; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21079.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_valid = _T_853[14]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21078.4]
  assign NV_NVDLA_CDMA_CVT_cell_14_io_chn_data_in_rsc_bits = _T_245_14; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21076.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_reset = reset; // @[:@20858.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21087.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21094.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21095.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21096.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_valid = _T_853[15]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21093.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_chn_alu_in_rsc_bits = _T_283_15; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21091.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_valid = _T_853[15]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21090.4]
  assign NV_NVDLA_CDMA_CVT_cell_15_io_chn_data_in_rsc_bits = _T_245_15; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21088.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_reset = reset; // @[:@20861.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21099.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21106.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21107.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21108.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_valid = _T_853[16]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21105.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_chn_alu_in_rsc_bits = _T_283_16; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21103.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_valid = _T_853[16]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21102.4]
  assign NV_NVDLA_CDMA_CVT_cell_16_io_chn_data_in_rsc_bits = _T_245_16; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21100.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_reset = reset; // @[:@20864.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21111.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21118.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21119.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21120.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_valid = _T_853[17]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21117.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_chn_alu_in_rsc_bits = _T_283_17; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21115.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_valid = _T_853[17]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21114.4]
  assign NV_NVDLA_CDMA_CVT_cell_17_io_chn_data_in_rsc_bits = _T_245_17; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21112.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_reset = reset; // @[:@20867.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21123.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21130.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21131.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21132.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_valid = _T_853[18]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21129.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_chn_alu_in_rsc_bits = _T_283_18; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21127.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_valid = _T_853[18]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21126.4]
  assign NV_NVDLA_CDMA_CVT_cell_18_io_chn_data_in_rsc_bits = _T_245_18; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21124.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_reset = reset; // @[:@20870.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21135.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21142.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21143.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21144.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_valid = _T_853[19]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21141.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_chn_alu_in_rsc_bits = _T_283_19; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21139.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_valid = _T_853[19]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21138.4]
  assign NV_NVDLA_CDMA_CVT_cell_19_io_chn_data_in_rsc_bits = _T_245_19; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21136.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_reset = reset; // @[:@20873.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21147.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21154.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21155.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21156.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_valid = _T_853[20]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21153.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_chn_alu_in_rsc_bits = _T_283_20; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21151.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_valid = _T_853[20]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21150.4]
  assign NV_NVDLA_CDMA_CVT_cell_20_io_chn_data_in_rsc_bits = _T_245_20; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21148.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_reset = reset; // @[:@20876.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21159.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21166.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21167.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21168.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_valid = _T_853[21]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21165.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_chn_alu_in_rsc_bits = _T_283_21; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21163.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_valid = _T_853[21]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21162.4]
  assign NV_NVDLA_CDMA_CVT_cell_21_io_chn_data_in_rsc_bits = _T_245_21; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21160.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_reset = reset; // @[:@20879.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21171.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21178.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21179.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21180.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_valid = _T_853[22]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21177.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_chn_alu_in_rsc_bits = _T_283_22; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21175.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_valid = _T_853[22]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21174.4]
  assign NV_NVDLA_CDMA_CVT_cell_22_io_chn_data_in_rsc_bits = _T_245_22; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21172.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_reset = reset; // @[:@20882.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21183.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21190.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21191.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21192.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_valid = _T_853[23]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21189.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_chn_alu_in_rsc_bits = _T_283_23; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21187.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_valid = _T_853[23]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21186.4]
  assign NV_NVDLA_CDMA_CVT_cell_23_io_chn_data_in_rsc_bits = _T_245_23; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21184.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_reset = reset; // @[:@20885.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21195.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21202.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21203.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21204.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_valid = _T_853[24]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21201.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_chn_alu_in_rsc_bits = _T_283_24; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21199.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_valid = _T_853[24]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21198.4]
  assign NV_NVDLA_CDMA_CVT_cell_24_io_chn_data_in_rsc_bits = _T_245_24; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21196.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_reset = reset; // @[:@20888.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21207.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21214.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21215.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21216.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_valid = _T_853[25]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21213.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_chn_alu_in_rsc_bits = _T_283_25; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21211.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_valid = _T_853[25]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21210.4]
  assign NV_NVDLA_CDMA_CVT_cell_25_io_chn_data_in_rsc_bits = _T_245_25; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21208.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_reset = reset; // @[:@20891.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21219.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21226.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21227.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21228.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_valid = _T_853[26]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21225.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_chn_alu_in_rsc_bits = _T_283_26; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21223.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_valid = _T_853[26]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21222.4]
  assign NV_NVDLA_CDMA_CVT_cell_26_io_chn_data_in_rsc_bits = _T_245_26; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21220.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_reset = reset; // @[:@20894.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21231.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21238.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21239.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21240.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_valid = _T_853[27]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21237.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_chn_alu_in_rsc_bits = _T_283_27; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21235.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_valid = _T_853[27]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21234.4]
  assign NV_NVDLA_CDMA_CVT_cell_27_io_chn_data_in_rsc_bits = _T_245_27; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21232.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_reset = reset; // @[:@20897.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21243.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21250.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21251.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21252.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_valid = _T_853[28]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21249.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_chn_alu_in_rsc_bits = _T_283_28; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21247.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_valid = _T_853[28]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21246.4]
  assign NV_NVDLA_CDMA_CVT_cell_28_io_chn_data_in_rsc_bits = _T_245_28; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21244.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_reset = reset; // @[:@20900.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21255.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21262.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21263.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21264.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_valid = _T_853[29]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21261.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_chn_alu_in_rsc_bits = _T_283_29; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21259.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_valid = _T_853[29]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21258.4]
  assign NV_NVDLA_CDMA_CVT_cell_29_io_chn_data_in_rsc_bits = _T_245_29; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21256.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_reset = reset; // @[:@20903.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21267.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21274.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21275.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21276.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_valid = _T_853[30]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21273.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_chn_alu_in_rsc_bits = _T_283_30; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21271.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_valid = _T_853[30]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21270.4]
  assign NV_NVDLA_CDMA_CVT_cell_30_io_chn_data_in_rsc_bits = _T_245_30; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21268.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_reset = reset; // @[:@20906.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_nvdla_core_clk = io_nvdla_hls_clk; // @[NV_NVDLA_CDMA_cvt.scala 238:33:@21279.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_cfg_mul_in_rsc = _T_95; // @[NV_NVDLA_CDMA_cvt.scala 246:33:@21286.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_cfg_out_precision = _T_92; // @[NV_NVDLA_CDMA_cvt.scala 247:36:@21287.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_cfg_truncate = _T_98; // @[NV_NVDLA_CDMA_cvt.scala 248:31:@21288.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_valid = _T_853[31]; // @[NV_NVDLA_CDMA_cvt.scala 244:39:@21285.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_chn_alu_in_rsc_bits = _T_283_31; // @[NV_NVDLA_CDMA_cvt.scala 243:38:@21283.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_valid = _T_853[31]; // @[NV_NVDLA_CDMA_cvt.scala 241:40:@21282.4]
  assign NV_NVDLA_CDMA_CVT_cell_31_io_chn_data_in_rsc_bits = _T_245_31; // @[NV_NVDLA_CDMA_cvt.scala 240:39:@21280.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_89 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_92 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_95 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_98 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_101 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_104 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_113 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_206 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_209 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_212 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {16{`RANDOM}};
  _T_214 = _RAND_10[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {8{`RANDOM}};
  _T_216 = _RAND_11[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_219 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_222 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_225 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_228 = _RAND_15[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_231 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_234 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_237 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_245_0 = _RAND_19[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_245_1 = _RAND_20[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_245_2 = _RAND_21[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_245_3 = _RAND_22[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_245_4 = _RAND_23[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_245_5 = _RAND_24[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_245_6 = _RAND_25[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_245_7 = _RAND_26[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_245_8 = _RAND_27[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_245_9 = _RAND_28[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_245_10 = _RAND_29[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_245_11 = _RAND_30[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_245_12 = _RAND_31[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_245_13 = _RAND_32[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_245_14 = _RAND_33[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_245_15 = _RAND_34[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_245_16 = _RAND_35[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_245_17 = _RAND_36[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_245_18 = _RAND_37[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_245_19 = _RAND_38[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_245_20 = _RAND_39[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_245_21 = _RAND_40[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_245_22 = _RAND_41[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_245_23 = _RAND_42[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_245_24 = _RAND_43[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_245_25 = _RAND_44[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_245_26 = _RAND_45[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_245_27 = _RAND_46[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_245_28 = _RAND_47[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_245_29 = _RAND_48[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_245_30 = _RAND_49[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_245_31 = _RAND_50[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_283_0 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_283_1 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_283_2 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_283_3 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_283_4 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_283_5 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_283_6 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_283_7 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_283_8 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_283_9 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_283_10 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_283_11 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_283_12 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_283_13 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_283_14 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_283_15 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_283_16 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_283_17 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_283_18 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_283_19 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_283_20 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_283_21 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_283_22 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_283_23 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_283_24 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_283_25 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_283_26 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_283_27 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_283_28 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_283_29 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_283_30 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_283_31 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_850 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_853 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1094 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1097 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1100 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1108 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1111 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1114 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1117 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1122 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1125 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1128 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1131 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1150 = _RAND_96[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1153 = _RAND_97[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1156 = _RAND_98[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1159 = _RAND_99[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1164 = _RAND_100[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1167 = _RAND_101[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1170 = _RAND_102[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1173 = _RAND_103[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1178 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1181 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1184 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1187 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1213 = _RAND_108[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {8{`RANDOM}};
  _T_1419 = _RAND_109[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1434 = _RAND_110[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1437 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1440 = _RAND_112[16:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_89 <= 1'h0;
    end else begin
      _T_89 <= _T_127;
    end
    if (reset) begin
      _T_92 <= 2'h0;
    end else begin
      if (_T_129) begin
        _T_92 <= io_reg2dp_proc_precision;
      end
    end
    if (reset) begin
      _T_95 <= 16'h0;
    end else begin
      if (_T_129) begin
        _T_95 <= io_reg2dp_cvt_scale;
      end
    end
    if (reset) begin
      _T_98 <= 6'h0;
    end else begin
      if (_T_129) begin
        _T_98 <= io_reg2dp_cvt_truncate;
      end
    end
    if (reset) begin
      _T_101 <= 16'h0;
    end else begin
      if (_T_129) begin
        _T_101 <= io_reg2dp_cvt_offset;
      end
    end
    if (reset) begin
      _T_104 <= 6'h0;
    end else begin
      if (_T_129) begin
        if (io_reg2dp_cvt_en) begin
          _T_104 <= 6'h3f;
        end else begin
          _T_104 <= 6'h0;
        end
      end
    end
    if (reset) begin
      _T_113 <= 16'h0;
    end else begin
      if (_T_129) begin
        _T_113 <= io_reg2dp_pad_value;
      end
    end
    if (reset) begin
      _T_206 <= 1'h0;
    end else begin
      _T_206 <= _T_165;
    end
    if (reset) begin
      _T_209 <= 1'h0;
    end else begin
      if (_T_165) begin
        _T_209 <= _T_162;
      end
    end
    if (reset) begin
      _T_212 <= 1'h0;
    end else begin
      if (_T_165) begin
        _T_212 <= _T_163;
      end
    end
    if (_T_165) begin
      if (_T_162) begin
        _T_214 <= io_img2cvt_mn_wr_data;
      end
    end
    if (_T_165) begin
      _T_216 <= _T_192;
    end
    if (reset) begin
      _T_219 <= 32'h0;
    end else begin
      if (_T_241) begin
        if (_T_196) begin
          if (_T_197) begin
            _T_219 <= 32'hffffffff;
          end else begin
            _T_219 <= 32'h0;
          end
        end else begin
          _T_219 <= 32'h0;
        end
      end
    end
    if (reset) begin
      _T_222 <= 1'h0;
    end else begin
      _T_222 <= _T_165;
    end
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= io_img2cvt_dat_wr_addr_valid;
    end
    if (reset) begin
      _T_228 <= 17'h0;
    end else begin
      if (_T_165) begin
        _T_228 <= _T_181;
      end
    end
    if (reset) begin
      _T_231 <= 4'h0;
    end else begin
      if (_T_165) begin
        _T_231 <= _T_161;
      end
    end
    if (reset) begin
      _T_234 <= 32'h0;
    end else begin
      if (io_img2cvt_dat_wr_addr_valid) begin
        if (io_img2cvt_dat_wr_addr_valid) begin
          _T_234 <= io_img2cvt_dat_wr_pad_mask;
        end else begin
          _T_234 <= 32'h0;
        end
      end
    end
    if (reset) begin
      _T_237 <= 2'h0;
    end else begin
      if (_T_165) begin
        _T_237 <= {{1'd0}, _T_168};
      end
    end
    if (_T_444) begin
      _T_245_0 <= _T_440;
    end
    if (_T_457) begin
      _T_245_1 <= _T_453;
    end
    if (_T_470) begin
      _T_245_2 <= _T_466;
    end
    if (_T_483) begin
      _T_245_3 <= _T_479;
    end
    if (_T_496) begin
      _T_245_4 <= _T_492;
    end
    if (_T_509) begin
      _T_245_5 <= _T_505;
    end
    if (_T_522) begin
      _T_245_6 <= _T_518;
    end
    if (_T_535) begin
      _T_245_7 <= _T_531;
    end
    if (_T_548) begin
      _T_245_8 <= _T_544;
    end
    if (_T_561) begin
      _T_245_9 <= _T_557;
    end
    if (_T_574) begin
      _T_245_10 <= _T_570;
    end
    if (_T_587) begin
      _T_245_11 <= _T_583;
    end
    if (_T_600) begin
      _T_245_12 <= _T_596;
    end
    if (_T_613) begin
      _T_245_13 <= _T_609;
    end
    if (_T_626) begin
      _T_245_14 <= _T_622;
    end
    if (_T_639) begin
      _T_245_15 <= _T_635;
    end
    if (_T_652) begin
      _T_245_16 <= _T_648;
    end
    if (_T_665) begin
      _T_245_17 <= _T_661;
    end
    if (_T_678) begin
      _T_245_18 <= _T_674;
    end
    if (_T_691) begin
      _T_245_19 <= _T_687;
    end
    if (_T_704) begin
      _T_245_20 <= _T_700;
    end
    if (_T_717) begin
      _T_245_21 <= _T_713;
    end
    if (_T_730) begin
      _T_245_22 <= _T_726;
    end
    if (_T_743) begin
      _T_245_23 <= _T_739;
    end
    if (_T_756) begin
      _T_245_24 <= _T_752;
    end
    if (_T_769) begin
      _T_245_25 <= _T_765;
    end
    if (_T_782) begin
      _T_245_26 <= _T_778;
    end
    if (_T_795) begin
      _T_245_27 <= _T_791;
    end
    if (_T_808) begin
      _T_245_28 <= _T_804;
    end
    if (_T_821) begin
      _T_245_29 <= _T_817;
    end
    if (_T_834) begin
      _T_245_30 <= _T_830;
    end
    if (_T_847) begin
      _T_245_31 <= _T_843;
    end
    if (_T_444) begin
      if (_T_209) begin
        _T_283_0 <= _T_441;
      end else begin
        _T_283_0 <= _T_101;
      end
    end
    if (_T_457) begin
      if (_T_209) begin
        _T_283_1 <= _T_454;
      end else begin
        _T_283_1 <= _T_101;
      end
    end
    if (_T_470) begin
      if (_T_209) begin
        _T_283_2 <= _T_467;
      end else begin
        _T_283_2 <= _T_101;
      end
    end
    if (_T_483) begin
      if (_T_209) begin
        _T_283_3 <= _T_480;
      end else begin
        _T_283_3 <= _T_101;
      end
    end
    if (_T_496) begin
      if (_T_209) begin
        _T_283_4 <= _T_493;
      end else begin
        _T_283_4 <= _T_101;
      end
    end
    if (_T_509) begin
      if (_T_209) begin
        _T_283_5 <= _T_506;
      end else begin
        _T_283_5 <= _T_101;
      end
    end
    if (_T_522) begin
      if (_T_209) begin
        _T_283_6 <= _T_519;
      end else begin
        _T_283_6 <= _T_101;
      end
    end
    if (_T_535) begin
      if (_T_209) begin
        _T_283_7 <= _T_532;
      end else begin
        _T_283_7 <= _T_101;
      end
    end
    if (_T_548) begin
      if (_T_209) begin
        _T_283_8 <= _T_545;
      end else begin
        _T_283_8 <= _T_101;
      end
    end
    if (_T_561) begin
      if (_T_209) begin
        _T_283_9 <= _T_558;
      end else begin
        _T_283_9 <= _T_101;
      end
    end
    if (_T_574) begin
      if (_T_209) begin
        _T_283_10 <= _T_571;
      end else begin
        _T_283_10 <= _T_101;
      end
    end
    if (_T_587) begin
      if (_T_209) begin
        _T_283_11 <= _T_584;
      end else begin
        _T_283_11 <= _T_101;
      end
    end
    if (_T_600) begin
      if (_T_209) begin
        _T_283_12 <= _T_597;
      end else begin
        _T_283_12 <= _T_101;
      end
    end
    if (_T_613) begin
      if (_T_209) begin
        _T_283_13 <= _T_610;
      end else begin
        _T_283_13 <= _T_101;
      end
    end
    if (_T_626) begin
      if (_T_209) begin
        _T_283_14 <= _T_623;
      end else begin
        _T_283_14 <= _T_101;
      end
    end
    if (_T_639) begin
      if (_T_209) begin
        _T_283_15 <= _T_636;
      end else begin
        _T_283_15 <= _T_101;
      end
    end
    if (_T_652) begin
      if (_T_209) begin
        _T_283_16 <= _T_649;
      end else begin
        _T_283_16 <= _T_101;
      end
    end
    if (_T_665) begin
      if (_T_209) begin
        _T_283_17 <= _T_662;
      end else begin
        _T_283_17 <= _T_101;
      end
    end
    if (_T_678) begin
      if (_T_209) begin
        _T_283_18 <= _T_675;
      end else begin
        _T_283_18 <= _T_101;
      end
    end
    if (_T_691) begin
      if (_T_209) begin
        _T_283_19 <= _T_688;
      end else begin
        _T_283_19 <= _T_101;
      end
    end
    if (_T_704) begin
      if (_T_209) begin
        _T_283_20 <= _T_701;
      end else begin
        _T_283_20 <= _T_101;
      end
    end
    if (_T_717) begin
      if (_T_209) begin
        _T_283_21 <= _T_714;
      end else begin
        _T_283_21 <= _T_101;
      end
    end
    if (_T_730) begin
      if (_T_209) begin
        _T_283_22 <= _T_727;
      end else begin
        _T_283_22 <= _T_101;
      end
    end
    if (_T_743) begin
      if (_T_209) begin
        _T_283_23 <= _T_740;
      end else begin
        _T_283_23 <= _T_101;
      end
    end
    if (_T_756) begin
      if (_T_209) begin
        _T_283_24 <= _T_753;
      end else begin
        _T_283_24 <= _T_101;
      end
    end
    if (_T_769) begin
      if (_T_209) begin
        _T_283_25 <= _T_766;
      end else begin
        _T_283_25 <= _T_101;
      end
    end
    if (_T_782) begin
      if (_T_209) begin
        _T_283_26 <= _T_779;
      end else begin
        _T_283_26 <= _T_101;
      end
    end
    if (_T_795) begin
      if (_T_209) begin
        _T_283_27 <= _T_792;
      end else begin
        _T_283_27 <= _T_101;
      end
    end
    if (_T_808) begin
      if (_T_209) begin
        _T_283_28 <= _T_805;
      end else begin
        _T_283_28 <= _T_101;
      end
    end
    if (_T_821) begin
      if (_T_209) begin
        _T_283_29 <= _T_818;
      end else begin
        _T_283_29 <= _T_101;
      end
    end
    if (_T_834) begin
      if (_T_209) begin
        _T_283_30 <= _T_831;
      end else begin
        _T_283_30 <= _T_101;
      end
    end
    if (_T_847) begin
      if (_T_209) begin
        _T_283_31 <= _T_844;
      end else begin
        _T_283_31 <= _T_101;
      end
    end
    if (reset) begin
      _T_850 <= 1'h0;
    end else begin
      _T_850 <= _T_206;
    end
    if (reset) begin
      _T_853 <= 32'h0;
    end else begin
      if (_T_854) begin
        _T_853 <= _T_219;
      end
    end
    if (reset) begin
      _T_1094 <= 1'h0;
    end else begin
      _T_1094 <= _T_222;
    end
    if (reset) begin
      _T_1097 <= 1'h0;
    end else begin
      _T_1097 <= _T_1094;
    end
    if (reset) begin
      _T_1100 <= 1'h0;
    end else begin
      _T_1100 <= _T_1097;
    end
    if (reset) begin
      _T_1108 <= 1'h0;
    end else begin
      _T_1108 <= _T_225;
    end
    if (reset) begin
      _T_1111 <= 1'h0;
    end else begin
      _T_1111 <= _T_1108;
    end
    if (reset) begin
      _T_1114 <= 1'h0;
    end else begin
      _T_1114 <= _T_1111;
    end
    if (reset) begin
      _T_1117 <= 1'h0;
    end else begin
      _T_1117 <= _T_1114;
    end
    if (reset) begin
      _T_1122 <= 1'h0;
    end else begin
      if (_T_222) begin
        _T_1122 <= _T_1119;
      end
    end
    if (reset) begin
      _T_1125 <= 1'h0;
    end else begin
      if (_T_1094) begin
        _T_1125 <= _T_1122;
      end
    end
    if (reset) begin
      _T_1128 <= 1'h0;
    end else begin
      if (_T_1097) begin
        _T_1128 <= _T_1125;
      end
    end
    if (reset) begin
      _T_1131 <= 1'h0;
    end else begin
      if (_T_1100) begin
        _T_1131 <= _T_1128;
      end
    end
    if (reset) begin
      _T_1150 <= 17'h0;
    end else begin
      _T_1150 <= _T_228;
    end
    if (reset) begin
      _T_1153 <= 17'h0;
    end else begin
      _T_1153 <= _T_1150;
    end
    if (reset) begin
      _T_1156 <= 17'h0;
    end else begin
      _T_1156 <= _T_1153;
    end
    if (reset) begin
      _T_1159 <= 17'h0;
    end else begin
      _T_1159 <= _T_1156;
    end
    if (reset) begin
      _T_1164 <= 4'h0;
    end else begin
      _T_1164 <= _T_231;
    end
    if (reset) begin
      _T_1167 <= 4'h0;
    end else begin
      _T_1167 <= _T_1164;
    end
    if (reset) begin
      _T_1170 <= 4'h0;
    end else begin
      _T_1170 <= _T_1167;
    end
    if (reset) begin
      _T_1173 <= 4'h0;
    end else begin
      _T_1173 <= _T_1170;
    end
    if (reset) begin
      _T_1178 <= 32'h0;
    end else begin
      _T_1178 <= _T_234;
    end
    if (reset) begin
      _T_1181 <= 32'h0;
    end else begin
      _T_1181 <= _T_1178;
    end
    if (reset) begin
      _T_1184 <= 32'h0;
    end else begin
      _T_1184 <= _T_1181;
    end
    if (reset) begin
      _T_1187 <= 32'h0;
    end else begin
      _T_1187 <= _T_1184;
    end
    if (reset) begin
      _T_1419 <= 256'h0;
    end else begin
      if (_T_1413) begin
        _T_1419 <= _T_1412;
      end else begin
        _T_1419 <= 256'h0;
      end
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_1213 <= 18'h0;
    end else begin
      if (_T_1445) begin
        _T_1213 <= _T_1443;
      end
    end
    if (reset) begin
      _T_1434 <= 2'h0;
    end else begin
      if (_T_1445) begin
        _T_1434 <= _T_1426;
      end else begin
        _T_1434 <= _T_1430;
      end
    end
    if (reset) begin
      _T_1437 <= 1'h0;
    end else begin
      _T_1437 <= _T_1420;
    end
    if (reset) begin
      _T_1440 <= 17'h0;
    end else begin
      if (_T_1420) begin
        if (_T_1445) begin
          _T_1440 <= _T_1421;
        end else begin
          if (_T_1192) begin
            _T_1440 <= _T_1159;
          end else begin
            _T_1440 <= _T_228;
          end
        end
      end
    end
  end
endmodule
module NV_NVDLA_slcg_5( // @[:@21738.2]
  input   io_nvdla_clock_nvdla_core_clk, // @[:@21741.4]
  output  io_nvdla_core_gated_clk // @[:@21741.4]
);
  assign io_nvdla_core_gated_clk = io_nvdla_clock_nvdla_core_clk; // @[slcg.scala 23:31:@21743.4]
endmodule
module nv_ram_rws( // @[:@21745.2]
  input          io_clk, // @[:@21748.4]
  input          io_re, // @[:@21748.4]
  input          io_we, // @[:@21748.4]
  input  [3:0]   io_ra, // @[:@21748.4]
  input  [3:0]   io_wa, // @[:@21748.4]
  input  [255:0] io_di, // @[:@21748.4]
  output [255:0] io_dout // @[:@21748.4]
);
  reg [255:0] _T_22_0; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_0;
  reg [255:0] _T_22_1; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_1;
  reg [255:0] _T_22_2; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_2;
  reg [255:0] _T_22_3; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_3;
  reg [255:0] _T_22_4; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_4;
  reg [255:0] _T_22_5; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_5;
  reg [255:0] _T_22_6; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_6;
  reg [255:0] _T_22_7; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_7;
  reg [255:0] _T_22_8; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_8;
  reg [255:0] _T_22_9; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_9;
  reg [255:0] _T_22_10; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_10;
  reg [255:0] _T_22_11; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_11;
  reg [255:0] _T_22_12; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_12;
  reg [255:0] _T_22_13; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_13;
  reg [255:0] _T_22_14; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_14;
  reg [255:0] _T_22_15; // @[nv_ram_rws.scala 27:18:@21750.4]
  reg [255:0] _RAND_15;
  reg [3:0] _T_42; // @[nv_ram_rws.scala 28:19:@21751.4]
  reg [31:0] _RAND_16;
  wire [255:0] _GEN_0; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_1; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_2; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_3; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_4; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_5; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_6; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_7; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_8; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_9; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_10; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_11; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_12; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_13; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_14; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_15; // @[nv_ram_rws.scala 31:20:@21753.6]
  wire [255:0] _GEN_34; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_35; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_36; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_37; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_38; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_39; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_40; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_41; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_42; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_43; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_44; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_45; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_46; // @[nv_ram_rws.scala 36:13:@21758.4]
  wire [255:0] _GEN_47; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_0 = 4'h0 == io_wa ? io_di : _T_22_0; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_1 = 4'h1 == io_wa ? io_di : _T_22_1; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_2 = 4'h2 == io_wa ? io_di : _T_22_2; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_3 = 4'h3 == io_wa ? io_di : _T_22_3; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_4 = 4'h4 == io_wa ? io_di : _T_22_4; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_5 = 4'h5 == io_wa ? io_di : _T_22_5; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_6 = 4'h6 == io_wa ? io_di : _T_22_6; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_7 = 4'h7 == io_wa ? io_di : _T_22_7; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_8 = 4'h8 == io_wa ? io_di : _T_22_8; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_9 = 4'h9 == io_wa ? io_di : _T_22_9; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_10 = 4'ha == io_wa ? io_di : _T_22_10; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_11 = 4'hb == io_wa ? io_di : _T_22_11; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_12 = 4'hc == io_wa ? io_di : _T_22_12; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_13 = 4'hd == io_wa ? io_di : _T_22_13; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_14 = 4'he == io_wa ? io_di : _T_22_14; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_15 = 4'hf == io_wa ? io_di : _T_22_15; // @[nv_ram_rws.scala 31:20:@21753.6]
  assign _GEN_34 = 4'h1 == _T_42 ? _T_22_1 : _T_22_0; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_35 = 4'h2 == _T_42 ? _T_22_2 : _GEN_34; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_36 = 4'h3 == _T_42 ? _T_22_3 : _GEN_35; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_37 = 4'h4 == _T_42 ? _T_22_4 : _GEN_36; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_38 = 4'h5 == _T_42 ? _T_22_5 : _GEN_37; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_39 = 4'h6 == _T_42 ? _T_22_6 : _GEN_38; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_40 = 4'h7 == _T_42 ? _T_22_7 : _GEN_39; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_41 = 4'h8 == _T_42 ? _T_22_8 : _GEN_40; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_42 = 4'h9 == _T_42 ? _T_22_9 : _GEN_41; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_43 = 4'ha == _T_42 ? _T_22_10 : _GEN_42; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_44 = 4'hb == _T_42 ? _T_22_11 : _GEN_43; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_45 = 4'hc == _T_42 ? _T_22_12 : _GEN_44; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_46 = 4'hd == _T_42 ? _T_22_13 : _GEN_45; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign _GEN_47 = 4'he == _T_42 ? _T_22_14 : _GEN_46; // @[nv_ram_rws.scala 36:13:@21758.4]
  assign io_dout = 4'hf == _T_42 ? _T_22_15 : _GEN_47; // @[nv_ram_rws.scala 36:13:@21758.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  _T_22_0 = _RAND_0[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {8{`RANDOM}};
  _T_22_1 = _RAND_1[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {8{`RANDOM}};
  _T_22_2 = _RAND_2[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {8{`RANDOM}};
  _T_22_3 = _RAND_3[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {8{`RANDOM}};
  _T_22_4 = _RAND_4[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {8{`RANDOM}};
  _T_22_5 = _RAND_5[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {8{`RANDOM}};
  _T_22_6 = _RAND_6[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {8{`RANDOM}};
  _T_22_7 = _RAND_7[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {8{`RANDOM}};
  _T_22_8 = _RAND_8[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {8{`RANDOM}};
  _T_22_9 = _RAND_9[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {8{`RANDOM}};
  _T_22_10 = _RAND_10[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {8{`RANDOM}};
  _T_22_11 = _RAND_11[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {8{`RANDOM}};
  _T_22_12 = _RAND_12[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {8{`RANDOM}};
  _T_22_13 = _RAND_13[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {8{`RANDOM}};
  _T_22_14 = _RAND_14[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {8{`RANDOM}};
  _T_22_15 = _RAND_15[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_42 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (4'h0 == io_wa) begin
        _T_22_0 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h1 == io_wa) begin
        _T_22_1 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h2 == io_wa) begin
        _T_22_2 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h3 == io_wa) begin
        _T_22_3 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h4 == io_wa) begin
        _T_22_4 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h5 == io_wa) begin
        _T_22_5 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h6 == io_wa) begin
        _T_22_6 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h7 == io_wa) begin
        _T_22_7 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h8 == io_wa) begin
        _T_22_8 <= io_di;
      end
    end
    if (io_we) begin
      if (4'h9 == io_wa) begin
        _T_22_9 <= io_di;
      end
    end
    if (io_we) begin
      if (4'ha == io_wa) begin
        _T_22_10 <= io_di;
      end
    end
    if (io_we) begin
      if (4'hb == io_wa) begin
        _T_22_11 <= io_di;
      end
    end
    if (io_we) begin
      if (4'hc == io_wa) begin
        _T_22_12 <= io_di;
      end
    end
    if (io_we) begin
      if (4'hd == io_wa) begin
        _T_22_13 <= io_di;
      end
    end
    if (io_we) begin
      if (4'he == io_wa) begin
        _T_22_14 <= io_di;
      end
    end
    if (io_we) begin
      if (4'hf == io_wa) begin
        _T_22_15 <= io_di;
      end
    end
    if (io_re) begin
      _T_42 <= io_ra;
    end
  end
endmodule
module NV_NVDLA_CDMA_shared_buffer( // @[:@21985.2]
  input          reset, // @[:@21987.4]
  input          io_nvdla_core_clk, // @[:@21988.4]
  input          io_dc2sbuf_p_wr_0_addr_valid, // @[:@21988.4]
  input  [7:0]   io_dc2sbuf_p_wr_0_addr_bits, // @[:@21988.4]
  input  [255:0] io_dc2sbuf_p_wr_0_data, // @[:@21988.4]
  input          io_img2sbuf_p_wr_0_addr_valid, // @[:@21988.4]
  input  [7:0]   io_img2sbuf_p_wr_0_addr_bits, // @[:@21988.4]
  input  [255:0] io_img2sbuf_p_wr_0_data, // @[:@21988.4]
  input          io_dc2sbuf_p_rd_0_addr_valid, // @[:@21988.4]
  input  [7:0]   io_dc2sbuf_p_rd_0_addr_bits, // @[:@21988.4]
  output [255:0] io_dc2sbuf_p_rd_0_data, // @[:@21988.4]
  input          io_img2sbuf_p_rd_0_addr_valid, // @[:@21988.4]
  input  [7:0]   io_img2sbuf_p_rd_0_addr_bits, // @[:@21988.4]
  output [255:0] io_img2sbuf_p_rd_0_data // @[:@21988.4]
);
  wire  nv_ram_rws_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire  nv_ram_rws_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire  nv_ram_rws_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire [3:0] nv_ram_rws_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire [3:0] nv_ram_rws_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire [255:0] nv_ram_rws_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire [255:0] nv_ram_rws_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
  wire  nv_ram_rws_1_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire  nv_ram_rws_1_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire  nv_ram_rws_1_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire [3:0] nv_ram_rws_1_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire [3:0] nv_ram_rws_1_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire [255:0] nv_ram_rws_1_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire [255:0] nv_ram_rws_1_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
  wire  nv_ram_rws_2_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire  nv_ram_rws_2_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire  nv_ram_rws_2_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire [3:0] nv_ram_rws_2_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire [3:0] nv_ram_rws_2_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire [255:0] nv_ram_rws_2_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire [255:0] nv_ram_rws_2_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
  wire  nv_ram_rws_3_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire  nv_ram_rws_3_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire  nv_ram_rws_3_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire [3:0] nv_ram_rws_3_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire [3:0] nv_ram_rws_3_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire [255:0] nv_ram_rws_3_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire [255:0] nv_ram_rws_3_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
  wire  nv_ram_rws_4_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire  nv_ram_rws_4_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire  nv_ram_rws_4_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire [3:0] nv_ram_rws_4_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire [3:0] nv_ram_rws_4_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire [255:0] nv_ram_rws_4_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire [255:0] nv_ram_rws_4_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
  wire  nv_ram_rws_5_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire  nv_ram_rws_5_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire  nv_ram_rws_5_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire [3:0] nv_ram_rws_5_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire [3:0] nv_ram_rws_5_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire [255:0] nv_ram_rws_5_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire [255:0] nv_ram_rws_5_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
  wire  nv_ram_rws_6_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire  nv_ram_rws_6_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire  nv_ram_rws_6_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire [3:0] nv_ram_rws_6_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire [3:0] nv_ram_rws_6_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire [255:0] nv_ram_rws_6_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire [255:0] nv_ram_rws_6_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
  wire  nv_ram_rws_7_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire  nv_ram_rws_7_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire  nv_ram_rws_7_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire [3:0] nv_ram_rws_7_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire [3:0] nv_ram_rws_7_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire [255:0] nv_ram_rws_7_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire [255:0] nv_ram_rws_7_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
  wire  nv_ram_rws_8_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire  nv_ram_rws_8_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire  nv_ram_rws_8_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire [3:0] nv_ram_rws_8_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire [3:0] nv_ram_rws_8_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire [255:0] nv_ram_rws_8_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire [255:0] nv_ram_rws_8_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
  wire  nv_ram_rws_9_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire  nv_ram_rws_9_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire  nv_ram_rws_9_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire [3:0] nv_ram_rws_9_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire [3:0] nv_ram_rws_9_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire [255:0] nv_ram_rws_9_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire [255:0] nv_ram_rws_9_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
  wire  nv_ram_rws_10_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire  nv_ram_rws_10_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire  nv_ram_rws_10_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire [3:0] nv_ram_rws_10_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire [3:0] nv_ram_rws_10_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire [255:0] nv_ram_rws_10_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire [255:0] nv_ram_rws_10_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
  wire  nv_ram_rws_11_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire  nv_ram_rws_11_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire  nv_ram_rws_11_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire [3:0] nv_ram_rws_11_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire [3:0] nv_ram_rws_11_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire [255:0] nv_ram_rws_11_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire [255:0] nv_ram_rws_11_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
  wire  nv_ram_rws_12_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire  nv_ram_rws_12_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire  nv_ram_rws_12_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire [3:0] nv_ram_rws_12_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire [3:0] nv_ram_rws_12_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire [255:0] nv_ram_rws_12_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire [255:0] nv_ram_rws_12_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
  wire  nv_ram_rws_13_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire  nv_ram_rws_13_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire  nv_ram_rws_13_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire [3:0] nv_ram_rws_13_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire [3:0] nv_ram_rws_13_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire [255:0] nv_ram_rws_13_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire [255:0] nv_ram_rws_13_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
  wire  nv_ram_rws_14_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire  nv_ram_rws_14_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire  nv_ram_rws_14_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire [3:0] nv_ram_rws_14_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire [3:0] nv_ram_rws_14_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire [255:0] nv_ram_rws_14_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire [255:0] nv_ram_rws_14_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
  wire  nv_ram_rws_15_io_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire  nv_ram_rws_15_io_re; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire  nv_ram_rws_15_io_we; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire [3:0] nv_ram_rws_15_io_ra; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire [3:0] nv_ram_rws_15_io_wa; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire [255:0] nv_ram_rws_15_io_di; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire [255:0] nv_ram_rws_15_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
  wire [3:0] _T_153; // @[NV_NVDLA_CDMA_shared_buffer.scala 56:54:@21990.4]
  wire [3:0] _T_154; // @[NV_NVDLA_CDMA_shared_buffer.scala 57:56:@21991.4]
  wire  _T_158; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21994.4]
  wire  _T_159; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21995.4]
  wire  _T_161; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21996.4]
  wire  _T_162; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21997.4]
  wire  _T_164; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21998.4]
  wire  _T_165; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21999.4]
  wire  _T_167; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22000.4]
  wire  _T_168; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22001.4]
  wire  _T_170; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22002.4]
  wire  _T_171; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22003.4]
  wire  _T_173; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22004.4]
  wire  _T_174; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22005.4]
  wire  _T_176; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22006.4]
  wire  _T_177; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22007.4]
  wire  _T_179; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22008.4]
  wire  _T_180; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22009.4]
  wire  _T_182; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22010.4]
  wire  _T_183; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22011.4]
  wire  _T_185; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22012.4]
  wire  _T_186; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22013.4]
  wire  _T_188; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22014.4]
  wire  _T_189; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22015.4]
  wire  _T_191; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22016.4]
  wire  _T_192; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22017.4]
  wire  _T_194; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22018.4]
  wire  _T_195; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22019.4]
  wire  _T_197; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22020.4]
  wire  _T_198; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22021.4]
  wire  _T_200; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22022.4]
  wire  _T_201; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22023.4]
  wire  _T_203; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22024.4]
  wire  _T_204; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22025.4]
  wire  _T_298; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22092.4]
  wire  _T_299; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22093.4]
  wire  _T_301; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22094.4]
  wire  _T_302; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22095.4]
  wire  _T_304; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22096.4]
  wire  _T_305; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22097.4]
  wire  _T_307; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22098.4]
  wire  _T_308; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22099.4]
  wire  _T_310; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22100.4]
  wire  _T_311; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22101.4]
  wire  _T_313; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22102.4]
  wire  _T_314; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22103.4]
  wire  _T_316; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22104.4]
  wire  _T_317; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22105.4]
  wire  _T_319; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22106.4]
  wire  _T_320; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22107.4]
  wire  _T_322; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22108.4]
  wire  _T_323; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22109.4]
  wire  _T_325; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22110.4]
  wire  _T_326; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22111.4]
  wire  _T_328; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22112.4]
  wire  _T_329; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22113.4]
  wire  _T_331; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22114.4]
  wire  _T_332; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22115.4]
  wire  _T_334; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22116.4]
  wire  _T_335; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22117.4]
  wire  _T_337; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22118.4]
  wire  _T_338; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22119.4]
  wire  _T_340; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22120.4]
  wire  _T_341; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22121.4]
  wire  _T_343; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22122.4]
  wire  _T_344; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22123.4]
  wire [7:0] _T_510; // @[Bitwise.scala 72:12:@22256.4]
  wire [3:0] _T_511; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:86:@22257.4]
  wire [7:0] _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22258.4]
  wire [7:0] _T_512; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22258.4]
  wire [7:0] _T_523; // @[Bitwise.scala 72:12:@22265.4]
  wire [3:0] _T_524; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:88:@22266.4]
  wire [7:0] _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22267.4]
  wire [7:0] _T_525; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22267.4]
  wire [7:0] _T_526; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22268.4]
  wire [7:0] _T_537; // @[Bitwise.scala 72:12:@22275.4]
  wire [7:0] _T_539; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22277.4]
  wire [7:0] _T_550; // @[Bitwise.scala 72:12:@22284.4]
  wire [7:0] _T_552; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22286.4]
  wire [7:0] _T_553; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22287.4]
  wire [7:0] _T_564; // @[Bitwise.scala 72:12:@22294.4]
  wire [7:0] _T_566; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22296.4]
  wire [7:0] _T_577; // @[Bitwise.scala 72:12:@22303.4]
  wire [7:0] _T_579; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22305.4]
  wire [7:0] _T_580; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22306.4]
  wire [7:0] _T_591; // @[Bitwise.scala 72:12:@22313.4]
  wire [7:0] _T_593; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22315.4]
  wire [7:0] _T_604; // @[Bitwise.scala 72:12:@22322.4]
  wire [7:0] _T_606; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22324.4]
  wire [7:0] _T_607; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22325.4]
  wire [7:0] _T_618; // @[Bitwise.scala 72:12:@22332.4]
  wire [7:0] _T_620; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22334.4]
  wire [7:0] _T_631; // @[Bitwise.scala 72:12:@22341.4]
  wire [7:0] _T_633; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22343.4]
  wire [7:0] _T_634; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22344.4]
  wire [7:0] _T_645; // @[Bitwise.scala 72:12:@22351.4]
  wire [7:0] _T_647; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22353.4]
  wire [7:0] _T_658; // @[Bitwise.scala 72:12:@22360.4]
  wire [7:0] _T_660; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22362.4]
  wire [7:0] _T_661; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22363.4]
  wire [7:0] _T_672; // @[Bitwise.scala 72:12:@22370.4]
  wire [7:0] _T_674; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22372.4]
  wire [7:0] _T_685; // @[Bitwise.scala 72:12:@22379.4]
  wire [7:0] _T_687; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22381.4]
  wire [7:0] _T_688; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22382.4]
  wire [7:0] _T_699; // @[Bitwise.scala 72:12:@22389.4]
  wire [7:0] _T_701; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22391.4]
  wire [7:0] _T_712; // @[Bitwise.scala 72:12:@22398.4]
  wire [7:0] _T_714; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22400.4]
  wire [7:0] _T_715; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22401.4]
  wire [7:0] _T_726; // @[Bitwise.scala 72:12:@22408.4]
  wire [7:0] _T_728; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22410.4]
  wire [7:0] _T_739; // @[Bitwise.scala 72:12:@22417.4]
  wire [7:0] _T_741; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22419.4]
  wire [7:0] _T_742; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22420.4]
  wire [7:0] _T_753; // @[Bitwise.scala 72:12:@22427.4]
  wire [7:0] _T_755; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22429.4]
  wire [7:0] _T_766; // @[Bitwise.scala 72:12:@22436.4]
  wire [7:0] _T_768; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22438.4]
  wire [7:0] _T_769; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22439.4]
  wire [7:0] _T_780; // @[Bitwise.scala 72:12:@22446.4]
  wire [7:0] _T_782; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22448.4]
  wire [7:0] _T_793; // @[Bitwise.scala 72:12:@22455.4]
  wire [7:0] _T_795; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22457.4]
  wire [7:0] _T_796; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22458.4]
  wire [7:0] _T_807; // @[Bitwise.scala 72:12:@22465.4]
  wire [7:0] _T_809; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22467.4]
  wire [7:0] _T_820; // @[Bitwise.scala 72:12:@22474.4]
  wire [7:0] _T_822; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22476.4]
  wire [7:0] _T_823; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22477.4]
  wire [7:0] _T_834; // @[Bitwise.scala 72:12:@22484.4]
  wire [7:0] _T_836; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22486.4]
  wire [7:0] _T_847; // @[Bitwise.scala 72:12:@22493.4]
  wire [7:0] _T_849; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22495.4]
  wire [7:0] _T_850; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22496.4]
  wire [7:0] _T_861; // @[Bitwise.scala 72:12:@22503.4]
  wire [7:0] _T_863; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22505.4]
  wire [7:0] _T_874; // @[Bitwise.scala 72:12:@22512.4]
  wire [7:0] _T_876; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22514.4]
  wire [7:0] _T_877; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22515.4]
  wire [7:0] _T_888; // @[Bitwise.scala 72:12:@22522.4]
  wire [7:0] _T_890; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22524.4]
  wire [7:0] _T_901; // @[Bitwise.scala 72:12:@22531.4]
  wire [7:0] _T_903; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22533.4]
  wire [7:0] _T_904; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22534.4]
  wire [7:0] _T_915; // @[Bitwise.scala 72:12:@22541.4]
  wire [7:0] _T_917; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22543.4]
  wire [7:0] _T_928; // @[Bitwise.scala 72:12:@22550.4]
  wire [7:0] _T_930; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22552.4]
  wire [7:0] _T_931; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22553.4]
  wire [255:0] _T_964; // @[Bitwise.scala 72:12:@22577.4]
  wire [255:0] _T_965; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22578.4]
  wire [255:0] _T_975; // @[Bitwise.scala 72:12:@22584.4]
  wire [255:0] _T_976; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22585.4]
  wire [255:0] _T_987; // @[Bitwise.scala 72:12:@22592.4]
  wire [255:0] _T_988; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22593.4]
  wire [255:0] _T_998; // @[Bitwise.scala 72:12:@22599.4]
  wire [255:0] _T_999; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22600.4]
  wire [255:0] _T_1010; // @[Bitwise.scala 72:12:@22607.4]
  wire [255:0] _T_1011; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22608.4]
  wire [255:0] _T_1021; // @[Bitwise.scala 72:12:@22614.4]
  wire [255:0] _T_1022; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22615.4]
  wire [255:0] _T_1033; // @[Bitwise.scala 72:12:@22622.4]
  wire [255:0] _T_1034; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22623.4]
  wire [255:0] _T_1044; // @[Bitwise.scala 72:12:@22629.4]
  wire [255:0] _T_1045; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22630.4]
  wire [255:0] _T_1056; // @[Bitwise.scala 72:12:@22637.4]
  wire [255:0] _T_1057; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22638.4]
  wire [255:0] _T_1067; // @[Bitwise.scala 72:12:@22644.4]
  wire [255:0] _T_1068; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22645.4]
  wire [255:0] _T_1079; // @[Bitwise.scala 72:12:@22652.4]
  wire [255:0] _T_1080; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22653.4]
  wire [255:0] _T_1090; // @[Bitwise.scala 72:12:@22659.4]
  wire [255:0] _T_1091; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22660.4]
  wire [255:0] _T_1102; // @[Bitwise.scala 72:12:@22667.4]
  wire [255:0] _T_1103; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22668.4]
  wire [255:0] _T_1113; // @[Bitwise.scala 72:12:@22674.4]
  wire [255:0] _T_1114; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22675.4]
  wire [255:0] _T_1125; // @[Bitwise.scala 72:12:@22682.4]
  wire [255:0] _T_1126; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22683.4]
  wire [255:0] _T_1136; // @[Bitwise.scala 72:12:@22689.4]
  wire [255:0] _T_1137; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22690.4]
  wire [255:0] _T_1148; // @[Bitwise.scala 72:12:@22697.4]
  wire [255:0] _T_1149; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22698.4]
  wire [255:0] _T_1159; // @[Bitwise.scala 72:12:@22704.4]
  wire [255:0] _T_1160; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22705.4]
  wire [255:0] _T_1171; // @[Bitwise.scala 72:12:@22712.4]
  wire [255:0] _T_1172; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22713.4]
  wire [255:0] _T_1182; // @[Bitwise.scala 72:12:@22719.4]
  wire [255:0] _T_1183; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22720.4]
  wire [255:0] _T_1194; // @[Bitwise.scala 72:12:@22727.4]
  wire [255:0] _T_1195; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22728.4]
  wire [255:0] _T_1205; // @[Bitwise.scala 72:12:@22734.4]
  wire [255:0] _T_1206; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22735.4]
  wire [255:0] _T_1217; // @[Bitwise.scala 72:12:@22742.4]
  wire [255:0] _T_1218; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22743.4]
  wire [255:0] _T_1228; // @[Bitwise.scala 72:12:@22749.4]
  wire [255:0] _T_1229; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22750.4]
  wire [255:0] _T_1240; // @[Bitwise.scala 72:12:@22757.4]
  wire [255:0] _T_1241; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22758.4]
  wire [255:0] _T_1251; // @[Bitwise.scala 72:12:@22764.4]
  wire [255:0] _T_1252; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22765.4]
  wire [255:0] _T_1263; // @[Bitwise.scala 72:12:@22772.4]
  wire [255:0] _T_1264; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22773.4]
  wire [255:0] _T_1274; // @[Bitwise.scala 72:12:@22779.4]
  wire [255:0] _T_1275; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22780.4]
  wire [255:0] _T_1286; // @[Bitwise.scala 72:12:@22787.4]
  wire [255:0] _T_1287; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22788.4]
  wire [255:0] _T_1297; // @[Bitwise.scala 72:12:@22794.4]
  wire [255:0] _T_1298; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22795.4]
  wire [255:0] _T_1309; // @[Bitwise.scala 72:12:@22802.4]
  wire [255:0] _T_1310; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22803.4]
  wire [255:0] _T_1320; // @[Bitwise.scala 72:12:@22809.4]
  wire [255:0] _T_1321; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22810.4]
  wire [3:0] _T_1351; // @[NV_NVDLA_CDMA_shared_buffer.scala 80:54:@22833.4]
  wire [3:0] _T_1352; // @[NV_NVDLA_CDMA_shared_buffer.scala 81:56:@22834.4]
  wire  _T_1356; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22837.4]
  wire  _T_1357; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22838.4]
  wire  _T_1359; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22839.4]
  wire  _T_1360; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22840.4]
  wire  _T_1362; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22841.4]
  wire  _T_1363; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22842.4]
  wire  _T_1365; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22843.4]
  wire  _T_1366; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22844.4]
  wire  _T_1368; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22845.4]
  wire  _T_1369; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22846.4]
  wire  _T_1371; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22847.4]
  wire  _T_1372; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22848.4]
  wire  _T_1374; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22849.4]
  wire  _T_1375; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22850.4]
  wire  _T_1377; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22851.4]
  wire  _T_1378; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22852.4]
  wire  _T_1380; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22853.4]
  wire  _T_1381; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22854.4]
  wire  _T_1383; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22855.4]
  wire  _T_1384; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22856.4]
  wire  _T_1386; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22857.4]
  wire  _T_1387; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22858.4]
  wire  _T_1389; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22859.4]
  wire  _T_1390; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22860.4]
  wire  _T_1392; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22861.4]
  wire  _T_1393; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22862.4]
  wire  _T_1395; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22863.4]
  wire  _T_1396; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22864.4]
  wire  _T_1398; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22865.4]
  wire  _T_1399; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22866.4]
  wire  _T_1401; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22867.4]
  wire  _T_1402; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22868.4]
  wire  _T_1496; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22935.4]
  wire  _T_1497; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22936.4]
  wire  _T_1499; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22937.4]
  wire  _T_1500; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22938.4]
  wire  _T_1502; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22939.4]
  wire  _T_1503; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22940.4]
  wire  _T_1505; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22941.4]
  wire  _T_1506; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22942.4]
  wire  _T_1508; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22943.4]
  wire  _T_1509; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22944.4]
  wire  _T_1511; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22945.4]
  wire  _T_1512; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22946.4]
  wire  _T_1514; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22947.4]
  wire  _T_1515; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22948.4]
  wire  _T_1517; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22949.4]
  wire  _T_1518; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22950.4]
  wire  _T_1520; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22951.4]
  wire  _T_1521; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22952.4]
  wire  _T_1523; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22953.4]
  wire  _T_1524; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22954.4]
  wire  _T_1526; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22955.4]
  wire  _T_1527; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22956.4]
  wire  _T_1529; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22957.4]
  wire  _T_1530; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22958.4]
  wire  _T_1532; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22959.4]
  wire  _T_1533; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22960.4]
  wire  _T_1535; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22961.4]
  wire  _T_1536; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22962.4]
  wire  _T_1538; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22963.4]
  wire  _T_1539; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22964.4]
  wire  _T_1541; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22965.4]
  wire  _T_1542; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22966.4]
  wire  _T_1635; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23033.4]
  wire  _T_1636; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23034.4]
  wire  _T_1637; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23035.4]
  wire  _T_1638; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23036.4]
  wire  _T_1639; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23037.4]
  wire  _T_1640; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23038.4]
  wire  _T_1641; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23039.4]
  wire  _T_1642; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23040.4]
  wire  _T_1643; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23041.4]
  wire  _T_1644; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23042.4]
  wire  _T_1645; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23043.4]
  wire  _T_1646; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23044.4]
  wire  _T_1647; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23045.4]
  wire  _T_1648; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23046.4]
  wire  _T_1649; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23047.4]
  wire  _T_1650; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23048.4]
  wire [7:0] _T_1752; // @[Bitwise.scala 72:12:@23133.4]
  wire [3:0] _T_1753; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:86:@23134.4]
  wire [7:0] _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23135.4]
  wire [7:0] _T_1754; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23135.4]
  wire [7:0] _T_1765; // @[Bitwise.scala 72:12:@23142.4]
  wire [3:0] _T_1766; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:88:@23143.4]
  wire [7:0] _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23144.4]
  wire [7:0] _T_1767; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23144.4]
  wire [7:0] _T_1768; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23145.4]
  wire [7:0] _T_1779; // @[Bitwise.scala 72:12:@23152.4]
  wire [7:0] _T_1781; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23154.4]
  wire [7:0] _T_1792; // @[Bitwise.scala 72:12:@23161.4]
  wire [7:0] _T_1794; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23163.4]
  wire [7:0] _T_1795; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23164.4]
  wire [7:0] _T_1806; // @[Bitwise.scala 72:12:@23171.4]
  wire [7:0] _T_1808; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23173.4]
  wire [7:0] _T_1819; // @[Bitwise.scala 72:12:@23180.4]
  wire [7:0] _T_1821; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23182.4]
  wire [7:0] _T_1822; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23183.4]
  wire [7:0] _T_1833; // @[Bitwise.scala 72:12:@23190.4]
  wire [7:0] _T_1835; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23192.4]
  wire [7:0] _T_1846; // @[Bitwise.scala 72:12:@23199.4]
  wire [7:0] _T_1848; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23201.4]
  wire [7:0] _T_1849; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23202.4]
  wire [7:0] _T_1860; // @[Bitwise.scala 72:12:@23209.4]
  wire [7:0] _T_1862; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23211.4]
  wire [7:0] _T_1873; // @[Bitwise.scala 72:12:@23218.4]
  wire [7:0] _T_1875; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23220.4]
  wire [7:0] _T_1876; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23221.4]
  wire [7:0] _T_1887; // @[Bitwise.scala 72:12:@23228.4]
  wire [7:0] _T_1889; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23230.4]
  wire [7:0] _T_1900; // @[Bitwise.scala 72:12:@23237.4]
  wire [7:0] _T_1902; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23239.4]
  wire [7:0] _T_1903; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23240.4]
  wire [7:0] _T_1914; // @[Bitwise.scala 72:12:@23247.4]
  wire [7:0] _T_1916; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23249.4]
  wire [7:0] _T_1927; // @[Bitwise.scala 72:12:@23256.4]
  wire [7:0] _T_1929; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23258.4]
  wire [7:0] _T_1930; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23259.4]
  wire [7:0] _T_1941; // @[Bitwise.scala 72:12:@23266.4]
  wire [7:0] _T_1943; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23268.4]
  wire [7:0] _T_1954; // @[Bitwise.scala 72:12:@23275.4]
  wire [7:0] _T_1956; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23277.4]
  wire [7:0] _T_1957; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23278.4]
  wire [7:0] _T_1968; // @[Bitwise.scala 72:12:@23285.4]
  wire [7:0] _T_1970; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23287.4]
  wire [7:0] _T_1981; // @[Bitwise.scala 72:12:@23294.4]
  wire [7:0] _T_1983; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23296.4]
  wire [7:0] _T_1984; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23297.4]
  wire [7:0] _T_1995; // @[Bitwise.scala 72:12:@23304.4]
  wire [7:0] _T_1997; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23306.4]
  wire [7:0] _T_2008; // @[Bitwise.scala 72:12:@23313.4]
  wire [7:0] _T_2010; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23315.4]
  wire [7:0] _T_2011; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23316.4]
  wire [7:0] _T_2022; // @[Bitwise.scala 72:12:@23323.4]
  wire [7:0] _T_2024; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23325.4]
  wire [7:0] _T_2035; // @[Bitwise.scala 72:12:@23332.4]
  wire [7:0] _T_2037; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23334.4]
  wire [7:0] _T_2038; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23335.4]
  wire [7:0] _T_2049; // @[Bitwise.scala 72:12:@23342.4]
  wire [7:0] _T_2051; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23344.4]
  wire [7:0] _T_2062; // @[Bitwise.scala 72:12:@23351.4]
  wire [7:0] _T_2064; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23353.4]
  wire [7:0] _T_2065; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23354.4]
  wire [7:0] _T_2076; // @[Bitwise.scala 72:12:@23361.4]
  wire [7:0] _T_2078; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23363.4]
  wire [7:0] _T_2089; // @[Bitwise.scala 72:12:@23370.4]
  wire [7:0] _T_2091; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23372.4]
  wire [7:0] _T_2092; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23373.4]
  wire [7:0] _T_2103; // @[Bitwise.scala 72:12:@23380.4]
  wire [7:0] _T_2105; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23382.4]
  wire [7:0] _T_2116; // @[Bitwise.scala 72:12:@23389.4]
  wire [7:0] _T_2118; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23391.4]
  wire [7:0] _T_2119; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23392.4]
  wire [7:0] _T_2130; // @[Bitwise.scala 72:12:@23399.4]
  wire [7:0] _T_2132; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23401.4]
  wire [7:0] _T_2143; // @[Bitwise.scala 72:12:@23408.4]
  wire [7:0] _T_2145; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23410.4]
  wire [7:0] _T_2146; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23411.4]
  wire [7:0] _T_2157; // @[Bitwise.scala 72:12:@23418.4]
  wire [7:0] _T_2159; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23420.4]
  wire [7:0] _T_2170; // @[Bitwise.scala 72:12:@23427.4]
  wire [7:0] _T_2172; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23429.4]
  wire [7:0] _T_2173; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23430.4]
  reg  _T_2299_0; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_0;
  reg  _T_2299_1; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_1;
  reg  _T_2299_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_2;
  reg  _T_2299_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_3;
  reg  _T_2299_4; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_4;
  reg  _T_2299_5; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_5;
  reg  _T_2299_6; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_6;
  reg  _T_2299_7; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_7;
  reg  _T_2299_8; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_8;
  reg  _T_2299_9; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_9;
  reg  _T_2299_10; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_10;
  reg  _T_2299_11; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_11;
  reg  _T_2299_12; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_12;
  reg  _T_2299_13; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_13;
  reg  _T_2299_14; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_14;
  reg  _T_2299_15; // @[NV_NVDLA_CDMA_shared_buffer.scala 120:33:@23631.4]
  reg [31:0] _RAND_15;
  wire  _T_2479; // @[NV_NVDLA_CDMA_shared_buffer.scala 127:62:@23682.4]
  reg  _T_2482; // @[NV_NVDLA_CDMA_shared_buffer.scala 127:31:@23683.4]
  reg [31:0] _RAND_16;
  wire [15:0] _T_2490; // @[Bitwise.scala 72:12:@23689.4]
  wire [255:0] _T_2206_0; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23508.4]
  wire [255:0] _GEN_66; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23690.4]
  wire [255:0] _T_2491; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23690.4]
  wire [15:0] _T_2495; // @[Bitwise.scala 72:12:@23692.4]
  wire [255:0] _T_2206_1; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23515.4]
  wire [255:0] _GEN_67; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23693.4]
  wire [255:0] _T_2496; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23693.4]
  wire [15:0] _T_2500; // @[Bitwise.scala 72:12:@23695.4]
  wire [255:0] _T_2206_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23522.4]
  wire [255:0] _GEN_68; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23696.4]
  wire [255:0] _T_2501; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23696.4]
  wire [15:0] _T_2505; // @[Bitwise.scala 72:12:@23698.4]
  wire [255:0] _T_2206_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23529.4]
  wire [255:0] _GEN_69; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23699.4]
  wire [255:0] _T_2506; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23699.4]
  wire [15:0] _T_2510; // @[Bitwise.scala 72:12:@23701.4]
  wire [255:0] _T_2206_4; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23536.4]
  wire [255:0] _GEN_70; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23702.4]
  wire [255:0] _T_2511; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23702.4]
  wire [15:0] _T_2515; // @[Bitwise.scala 72:12:@23704.4]
  wire [255:0] _T_2206_5; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23543.4]
  wire [255:0] _GEN_71; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23705.4]
  wire [255:0] _T_2516; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23705.4]
  wire [15:0] _T_2520; // @[Bitwise.scala 72:12:@23707.4]
  wire [255:0] _T_2206_6; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23550.4]
  wire [255:0] _GEN_72; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23708.4]
  wire [255:0] _T_2521; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23708.4]
  wire [15:0] _T_2525; // @[Bitwise.scala 72:12:@23710.4]
  wire [255:0] _T_2206_7; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23557.4]
  wire [255:0] _GEN_73; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23711.4]
  wire [255:0] _T_2526; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23711.4]
  wire [15:0] _T_2530; // @[Bitwise.scala 72:12:@23713.4]
  wire [255:0] _T_2206_8; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23564.4]
  wire [255:0] _GEN_74; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23714.4]
  wire [255:0] _T_2531; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23714.4]
  wire [15:0] _T_2535; // @[Bitwise.scala 72:12:@23716.4]
  wire [255:0] _T_2206_9; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23571.4]
  wire [255:0] _GEN_75; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23717.4]
  wire [255:0] _T_2536; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23717.4]
  wire [15:0] _T_2540; // @[Bitwise.scala 72:12:@23719.4]
  wire [255:0] _T_2206_10; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23578.4]
  wire [255:0] _GEN_76; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23720.4]
  wire [255:0] _T_2541; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23720.4]
  wire [15:0] _T_2545; // @[Bitwise.scala 72:12:@23722.4]
  wire [255:0] _T_2206_11; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23585.4]
  wire [255:0] _GEN_77; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23723.4]
  wire [255:0] _T_2546; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23723.4]
  wire [15:0] _T_2550; // @[Bitwise.scala 72:12:@23725.4]
  wire [255:0] _T_2206_12; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23592.4]
  wire [255:0] _GEN_78; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23726.4]
  wire [255:0] _T_2551; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23726.4]
  wire [15:0] _T_2555; // @[Bitwise.scala 72:12:@23728.4]
  wire [255:0] _T_2206_13; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23599.4]
  wire [255:0] _GEN_79; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23729.4]
  wire [255:0] _T_2556; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23729.4]
  wire [15:0] _T_2560; // @[Bitwise.scala 72:12:@23731.4]
  wire [255:0] _T_2206_14; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23606.4]
  wire [255:0] _GEN_80; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23732.4]
  wire [255:0] _T_2561; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23732.4]
  wire [15:0] _T_2565; // @[Bitwise.scala 72:12:@23734.4]
  wire [255:0] _T_2206_15; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23613.4]
  wire [255:0] _GEN_81; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23735.4]
  wire [255:0] _T_2566; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23735.4]
  wire [255:0] _T_2589; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23753.4]
  wire [255:0] _T_2590; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23754.4]
  wire [255:0] _T_2591; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23755.4]
  wire [255:0] _T_2592; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23756.4]
  wire [255:0] _T_2593; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23757.4]
  wire [255:0] _T_2594; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23758.4]
  wire [255:0] _T_2595; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23759.4]
  wire [255:0] _T_2596; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23760.4]
  wire [255:0] _T_2597; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23761.4]
  wire [255:0] _T_2598; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23762.4]
  wire [255:0] _T_2599; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23763.4]
  wire [255:0] _T_2600; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23764.4]
  wire [255:0] _T_2601; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23765.4]
  wire [255:0] _T_2602; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23766.4]
  wire [255:0] _T_2603; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23767.4]
  reg [255:0] _T_2722; // @[Reg.scala 11:16:@23848.4]
  reg [255:0] _RAND_17;
  nv_ram_rws nv_ram_rws ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23453.4]
    .io_clk(nv_ram_rws_io_clk),
    .io_re(nv_ram_rws_io_re),
    .io_we(nv_ram_rws_io_we),
    .io_ra(nv_ram_rws_io_ra),
    .io_wa(nv_ram_rws_io_wa),
    .io_di(nv_ram_rws_io_di),
    .io_dout(nv_ram_rws_io_dout)
  );
  nv_ram_rws nv_ram_rws_1 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23456.4]
    .io_clk(nv_ram_rws_1_io_clk),
    .io_re(nv_ram_rws_1_io_re),
    .io_we(nv_ram_rws_1_io_we),
    .io_ra(nv_ram_rws_1_io_ra),
    .io_wa(nv_ram_rws_1_io_wa),
    .io_di(nv_ram_rws_1_io_di),
    .io_dout(nv_ram_rws_1_io_dout)
  );
  nv_ram_rws nv_ram_rws_2 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23459.4]
    .io_clk(nv_ram_rws_2_io_clk),
    .io_re(nv_ram_rws_2_io_re),
    .io_we(nv_ram_rws_2_io_we),
    .io_ra(nv_ram_rws_2_io_ra),
    .io_wa(nv_ram_rws_2_io_wa),
    .io_di(nv_ram_rws_2_io_di),
    .io_dout(nv_ram_rws_2_io_dout)
  );
  nv_ram_rws nv_ram_rws_3 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23462.4]
    .io_clk(nv_ram_rws_3_io_clk),
    .io_re(nv_ram_rws_3_io_re),
    .io_we(nv_ram_rws_3_io_we),
    .io_ra(nv_ram_rws_3_io_ra),
    .io_wa(nv_ram_rws_3_io_wa),
    .io_di(nv_ram_rws_3_io_di),
    .io_dout(nv_ram_rws_3_io_dout)
  );
  nv_ram_rws nv_ram_rws_4 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23465.4]
    .io_clk(nv_ram_rws_4_io_clk),
    .io_re(nv_ram_rws_4_io_re),
    .io_we(nv_ram_rws_4_io_we),
    .io_ra(nv_ram_rws_4_io_ra),
    .io_wa(nv_ram_rws_4_io_wa),
    .io_di(nv_ram_rws_4_io_di),
    .io_dout(nv_ram_rws_4_io_dout)
  );
  nv_ram_rws nv_ram_rws_5 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23468.4]
    .io_clk(nv_ram_rws_5_io_clk),
    .io_re(nv_ram_rws_5_io_re),
    .io_we(nv_ram_rws_5_io_we),
    .io_ra(nv_ram_rws_5_io_ra),
    .io_wa(nv_ram_rws_5_io_wa),
    .io_di(nv_ram_rws_5_io_di),
    .io_dout(nv_ram_rws_5_io_dout)
  );
  nv_ram_rws nv_ram_rws_6 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23471.4]
    .io_clk(nv_ram_rws_6_io_clk),
    .io_re(nv_ram_rws_6_io_re),
    .io_we(nv_ram_rws_6_io_we),
    .io_ra(nv_ram_rws_6_io_ra),
    .io_wa(nv_ram_rws_6_io_wa),
    .io_di(nv_ram_rws_6_io_di),
    .io_dout(nv_ram_rws_6_io_dout)
  );
  nv_ram_rws nv_ram_rws_7 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23474.4]
    .io_clk(nv_ram_rws_7_io_clk),
    .io_re(nv_ram_rws_7_io_re),
    .io_we(nv_ram_rws_7_io_we),
    .io_ra(nv_ram_rws_7_io_ra),
    .io_wa(nv_ram_rws_7_io_wa),
    .io_di(nv_ram_rws_7_io_di),
    .io_dout(nv_ram_rws_7_io_dout)
  );
  nv_ram_rws nv_ram_rws_8 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23477.4]
    .io_clk(nv_ram_rws_8_io_clk),
    .io_re(nv_ram_rws_8_io_re),
    .io_we(nv_ram_rws_8_io_we),
    .io_ra(nv_ram_rws_8_io_ra),
    .io_wa(nv_ram_rws_8_io_wa),
    .io_di(nv_ram_rws_8_io_di),
    .io_dout(nv_ram_rws_8_io_dout)
  );
  nv_ram_rws nv_ram_rws_9 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23480.4]
    .io_clk(nv_ram_rws_9_io_clk),
    .io_re(nv_ram_rws_9_io_re),
    .io_we(nv_ram_rws_9_io_we),
    .io_ra(nv_ram_rws_9_io_ra),
    .io_wa(nv_ram_rws_9_io_wa),
    .io_di(nv_ram_rws_9_io_di),
    .io_dout(nv_ram_rws_9_io_dout)
  );
  nv_ram_rws nv_ram_rws_10 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23483.4]
    .io_clk(nv_ram_rws_10_io_clk),
    .io_re(nv_ram_rws_10_io_re),
    .io_we(nv_ram_rws_10_io_we),
    .io_ra(nv_ram_rws_10_io_ra),
    .io_wa(nv_ram_rws_10_io_wa),
    .io_di(nv_ram_rws_10_io_di),
    .io_dout(nv_ram_rws_10_io_dout)
  );
  nv_ram_rws nv_ram_rws_11 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23486.4]
    .io_clk(nv_ram_rws_11_io_clk),
    .io_re(nv_ram_rws_11_io_re),
    .io_we(nv_ram_rws_11_io_we),
    .io_ra(nv_ram_rws_11_io_ra),
    .io_wa(nv_ram_rws_11_io_wa),
    .io_di(nv_ram_rws_11_io_di),
    .io_dout(nv_ram_rws_11_io_dout)
  );
  nv_ram_rws nv_ram_rws_12 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23489.4]
    .io_clk(nv_ram_rws_12_io_clk),
    .io_re(nv_ram_rws_12_io_re),
    .io_we(nv_ram_rws_12_io_we),
    .io_ra(nv_ram_rws_12_io_ra),
    .io_wa(nv_ram_rws_12_io_wa),
    .io_di(nv_ram_rws_12_io_di),
    .io_dout(nv_ram_rws_12_io_dout)
  );
  nv_ram_rws nv_ram_rws_13 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23492.4]
    .io_clk(nv_ram_rws_13_io_clk),
    .io_re(nv_ram_rws_13_io_re),
    .io_we(nv_ram_rws_13_io_we),
    .io_ra(nv_ram_rws_13_io_ra),
    .io_wa(nv_ram_rws_13_io_wa),
    .io_di(nv_ram_rws_13_io_di),
    .io_dout(nv_ram_rws_13_io_dout)
  );
  nv_ram_rws nv_ram_rws_14 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23495.4]
    .io_clk(nv_ram_rws_14_io_clk),
    .io_re(nv_ram_rws_14_io_re),
    .io_we(nv_ram_rws_14_io_we),
    .io_ra(nv_ram_rws_14_io_ra),
    .io_wa(nv_ram_rws_14_io_wa),
    .io_di(nv_ram_rws_14_io_di),
    .io_dout(nv_ram_rws_14_io_dout)
  );
  nv_ram_rws nv_ram_rws_15 ( // @[NV_NVDLA_CDMA_shared_buffer.scala 105:63:@23498.4]
    .io_clk(nv_ram_rws_15_io_clk),
    .io_re(nv_ram_rws_15_io_re),
    .io_we(nv_ram_rws_15_io_we),
    .io_ra(nv_ram_rws_15_io_ra),
    .io_wa(nv_ram_rws_15_io_wa),
    .io_di(nv_ram_rws_15_io_di),
    .io_dout(nv_ram_rws_15_io_dout)
  );
  assign _T_153 = io_dc2sbuf_p_wr_0_addr_bits[7:4]; // @[NV_NVDLA_CDMA_shared_buffer.scala 56:54:@21990.4]
  assign _T_154 = io_img2sbuf_p_wr_0_addr_bits[7:4]; // @[NV_NVDLA_CDMA_shared_buffer.scala 57:56:@21991.4]
  assign _T_158 = _T_153 == 4'h0; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21994.4]
  assign _T_159 = _T_158 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21995.4]
  assign _T_161 = _T_153 == 4'h1; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21996.4]
  assign _T_162 = _T_161 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21997.4]
  assign _T_164 = _T_153 == 4'h2; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@21998.4]
  assign _T_165 = _T_164 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@21999.4]
  assign _T_167 = _T_153 == 4'h3; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22000.4]
  assign _T_168 = _T_167 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22001.4]
  assign _T_170 = _T_153 == 4'h4; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22002.4]
  assign _T_171 = _T_170 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22003.4]
  assign _T_173 = _T_153 == 4'h5; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22004.4]
  assign _T_174 = _T_173 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22005.4]
  assign _T_176 = _T_153 == 4'h6; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22006.4]
  assign _T_177 = _T_176 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22007.4]
  assign _T_179 = _T_153 == 4'h7; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22008.4]
  assign _T_180 = _T_179 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22009.4]
  assign _T_182 = _T_153 == 4'h8; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22010.4]
  assign _T_183 = _T_182 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22011.4]
  assign _T_185 = _T_153 == 4'h9; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22012.4]
  assign _T_186 = _T_185 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22013.4]
  assign _T_188 = _T_153 == 4'ha; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22014.4]
  assign _T_189 = _T_188 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22015.4]
  assign _T_191 = _T_153 == 4'hb; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22016.4]
  assign _T_192 = _T_191 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22017.4]
  assign _T_194 = _T_153 == 4'hc; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22018.4]
  assign _T_195 = _T_194 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22019.4]
  assign _T_197 = _T_153 == 4'hd; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22020.4]
  assign _T_198 = _T_197 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22021.4]
  assign _T_200 = _T_153 == 4'he; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22022.4]
  assign _T_201 = _T_200 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22023.4]
  assign _T_203 = _T_153 == 4'hf; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:94:@22024.4]
  assign _T_204 = _T_203 & io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 61:102:@22025.4]
  assign _T_298 = _T_154 == 4'h0; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22092.4]
  assign _T_299 = _T_298 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22093.4]
  assign _T_301 = _T_154 == 4'h1; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22094.4]
  assign _T_302 = _T_301 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22095.4]
  assign _T_304 = _T_154 == 4'h2; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22096.4]
  assign _T_305 = _T_304 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22097.4]
  assign _T_307 = _T_154 == 4'h3; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22098.4]
  assign _T_308 = _T_307 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22099.4]
  assign _T_310 = _T_154 == 4'h4; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22100.4]
  assign _T_311 = _T_310 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22101.4]
  assign _T_313 = _T_154 == 4'h5; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22102.4]
  assign _T_314 = _T_313 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22103.4]
  assign _T_316 = _T_154 == 4'h6; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22104.4]
  assign _T_317 = _T_316 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22105.4]
  assign _T_319 = _T_154 == 4'h7; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22106.4]
  assign _T_320 = _T_319 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22107.4]
  assign _T_322 = _T_154 == 4'h8; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22108.4]
  assign _T_323 = _T_322 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22109.4]
  assign _T_325 = _T_154 == 4'h9; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22110.4]
  assign _T_326 = _T_325 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22111.4]
  assign _T_328 = _T_154 == 4'ha; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22112.4]
  assign _T_329 = _T_328 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22113.4]
  assign _T_331 = _T_154 == 4'hb; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22114.4]
  assign _T_332 = _T_331 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22115.4]
  assign _T_334 = _T_154 == 4'hc; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22116.4]
  assign _T_335 = _T_334 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22117.4]
  assign _T_337 = _T_154 == 4'hd; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22118.4]
  assign _T_338 = _T_337 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22119.4]
  assign _T_340 = _T_154 == 4'he; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22120.4]
  assign _T_341 = _T_340 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22121.4]
  assign _T_343 = _T_154 == 4'hf; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:96:@22122.4]
  assign _T_344 = _T_343 & io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 63:104:@22123.4]
  assign _T_510 = _T_159 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22256.4]
  assign _T_511 = io_dc2sbuf_p_wr_0_addr_bits[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:86:@22257.4]
  assign _GEN_2 = {{4'd0}, _T_511}; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22258.4]
  assign _T_512 = _T_510 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22258.4]
  assign _T_523 = _T_299 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22265.4]
  assign _T_524 = io_img2sbuf_p_wr_0_addr_bits[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:88:@22266.4]
  assign _GEN_3 = {{4'd0}, _T_524}; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22267.4]
  assign _T_525 = _T_523 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22267.4]
  assign _T_526 = _T_512 | _T_525; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22268.4]
  assign _T_537 = _T_162 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22275.4]
  assign _T_539 = _T_537 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22277.4]
  assign _T_550 = _T_302 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22284.4]
  assign _T_552 = _T_550 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22286.4]
  assign _T_553 = _T_539 | _T_552; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22287.4]
  assign _T_564 = _T_165 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22294.4]
  assign _T_566 = _T_564 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22296.4]
  assign _T_577 = _T_305 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22303.4]
  assign _T_579 = _T_577 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22305.4]
  assign _T_580 = _T_566 | _T_579; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22306.4]
  assign _T_591 = _T_168 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22313.4]
  assign _T_593 = _T_591 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22315.4]
  assign _T_604 = _T_308 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22322.4]
  assign _T_606 = _T_604 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22324.4]
  assign _T_607 = _T_593 | _T_606; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22325.4]
  assign _T_618 = _T_171 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22332.4]
  assign _T_620 = _T_618 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22334.4]
  assign _T_631 = _T_311 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22341.4]
  assign _T_633 = _T_631 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22343.4]
  assign _T_634 = _T_620 | _T_633; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22344.4]
  assign _T_645 = _T_174 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22351.4]
  assign _T_647 = _T_645 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22353.4]
  assign _T_658 = _T_314 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22360.4]
  assign _T_660 = _T_658 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22362.4]
  assign _T_661 = _T_647 | _T_660; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22363.4]
  assign _T_672 = _T_177 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22370.4]
  assign _T_674 = _T_672 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22372.4]
  assign _T_685 = _T_317 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22379.4]
  assign _T_687 = _T_685 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22381.4]
  assign _T_688 = _T_674 | _T_687; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22382.4]
  assign _T_699 = _T_180 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22389.4]
  assign _T_701 = _T_699 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22391.4]
  assign _T_712 = _T_320 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22398.4]
  assign _T_714 = _T_712 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22400.4]
  assign _T_715 = _T_701 | _T_714; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22401.4]
  assign _T_726 = _T_183 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22408.4]
  assign _T_728 = _T_726 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22410.4]
  assign _T_739 = _T_323 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22417.4]
  assign _T_741 = _T_739 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22419.4]
  assign _T_742 = _T_728 | _T_741; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22420.4]
  assign _T_753 = _T_186 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22427.4]
  assign _T_755 = _T_753 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22429.4]
  assign _T_766 = _T_326 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22436.4]
  assign _T_768 = _T_766 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22438.4]
  assign _T_769 = _T_755 | _T_768; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22439.4]
  assign _T_780 = _T_189 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22446.4]
  assign _T_782 = _T_780 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22448.4]
  assign _T_793 = _T_329 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22455.4]
  assign _T_795 = _T_793 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22457.4]
  assign _T_796 = _T_782 | _T_795; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22458.4]
  assign _T_807 = _T_192 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22465.4]
  assign _T_809 = _T_807 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22467.4]
  assign _T_820 = _T_332 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22474.4]
  assign _T_822 = _T_820 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22476.4]
  assign _T_823 = _T_809 | _T_822; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22477.4]
  assign _T_834 = _T_195 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22484.4]
  assign _T_836 = _T_834 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22486.4]
  assign _T_847 = _T_335 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22493.4]
  assign _T_849 = _T_847 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22495.4]
  assign _T_850 = _T_836 | _T_849; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22496.4]
  assign _T_861 = _T_198 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22503.4]
  assign _T_863 = _T_861 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22505.4]
  assign _T_874 = _T_338 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22512.4]
  assign _T_876 = _T_874 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22514.4]
  assign _T_877 = _T_863 | _T_876; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22515.4]
  assign _T_888 = _T_201 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22522.4]
  assign _T_890 = _T_888 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22524.4]
  assign _T_901 = _T_341 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22531.4]
  assign _T_903 = _T_901 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22533.4]
  assign _T_904 = _T_890 | _T_903; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22534.4]
  assign _T_915 = _T_204 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22541.4]
  assign _T_917 = _T_915 & _GEN_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 68:57:@22543.4]
  assign _T_928 = _T_344 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@22550.4]
  assign _T_930 = _T_928 & _GEN_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 70:58:@22552.4]
  assign _T_931 = _T_917 | _T_930; // @[NV_NVDLA_CDMA_shared_buffer.scala 69:96:@22553.4]
  assign _T_964 = _T_159 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22577.4]
  assign _T_965 = _T_964 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22578.4]
  assign _T_975 = _T_299 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22584.4]
  assign _T_976 = _T_975 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22585.4]
  assign _T_987 = _T_162 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22592.4]
  assign _T_988 = _T_987 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22593.4]
  assign _T_998 = _T_302 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22599.4]
  assign _T_999 = _T_998 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22600.4]
  assign _T_1010 = _T_165 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22607.4]
  assign _T_1011 = _T_1010 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22608.4]
  assign _T_1021 = _T_305 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22614.4]
  assign _T_1022 = _T_1021 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22615.4]
  assign _T_1033 = _T_168 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22622.4]
  assign _T_1034 = _T_1033 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22623.4]
  assign _T_1044 = _T_308 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22629.4]
  assign _T_1045 = _T_1044 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22630.4]
  assign _T_1056 = _T_171 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22637.4]
  assign _T_1057 = _T_1056 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22638.4]
  assign _T_1067 = _T_311 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22644.4]
  assign _T_1068 = _T_1067 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22645.4]
  assign _T_1079 = _T_174 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22652.4]
  assign _T_1080 = _T_1079 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22653.4]
  assign _T_1090 = _T_314 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22659.4]
  assign _T_1091 = _T_1090 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22660.4]
  assign _T_1102 = _T_177 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22667.4]
  assign _T_1103 = _T_1102 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22668.4]
  assign _T_1113 = _T_317 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22674.4]
  assign _T_1114 = _T_1113 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22675.4]
  assign _T_1125 = _T_180 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22682.4]
  assign _T_1126 = _T_1125 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22683.4]
  assign _T_1136 = _T_320 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22689.4]
  assign _T_1137 = _T_1136 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22690.4]
  assign _T_1148 = _T_183 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22697.4]
  assign _T_1149 = _T_1148 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22698.4]
  assign _T_1159 = _T_323 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22704.4]
  assign _T_1160 = _T_1159 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22705.4]
  assign _T_1171 = _T_186 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22712.4]
  assign _T_1172 = _T_1171 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22713.4]
  assign _T_1182 = _T_326 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22719.4]
  assign _T_1183 = _T_1182 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22720.4]
  assign _T_1194 = _T_189 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22727.4]
  assign _T_1195 = _T_1194 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22728.4]
  assign _T_1205 = _T_329 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22734.4]
  assign _T_1206 = _T_1205 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22735.4]
  assign _T_1217 = _T_192 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22742.4]
  assign _T_1218 = _T_1217 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22743.4]
  assign _T_1228 = _T_332 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22749.4]
  assign _T_1229 = _T_1228 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22750.4]
  assign _T_1240 = _T_195 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22757.4]
  assign _T_1241 = _T_1240 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22758.4]
  assign _T_1251 = _T_335 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22764.4]
  assign _T_1252 = _T_1251 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22765.4]
  assign _T_1263 = _T_198 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22772.4]
  assign _T_1264 = _T_1263 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22773.4]
  assign _T_1274 = _T_338 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22779.4]
  assign _T_1275 = _T_1274 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22780.4]
  assign _T_1286 = _T_201 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22787.4]
  assign _T_1287 = _T_1286 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22788.4]
  assign _T_1297 = _T_341 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22794.4]
  assign _T_1298 = _T_1297 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22795.4]
  assign _T_1309 = _T_204 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22802.4]
  assign _T_1310 = _T_1309 & io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 74:80:@22803.4]
  assign _T_1320 = _T_344 ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12:@22809.4]
  assign _T_1321 = _T_1320 & io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_CDMA_shared_buffer.scala 76:81:@22810.4]
  assign _T_1351 = io_dc2sbuf_p_rd_0_addr_bits[7:4]; // @[NV_NVDLA_CDMA_shared_buffer.scala 80:54:@22833.4]
  assign _T_1352 = io_img2sbuf_p_rd_0_addr_bits[7:4]; // @[NV_NVDLA_CDMA_shared_buffer.scala 81:56:@22834.4]
  assign _T_1356 = _T_1351 == 4'h0; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22837.4]
  assign _T_1357 = _T_1356 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22838.4]
  assign _T_1359 = _T_1351 == 4'h1; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22839.4]
  assign _T_1360 = _T_1359 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22840.4]
  assign _T_1362 = _T_1351 == 4'h2; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22841.4]
  assign _T_1363 = _T_1362 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22842.4]
  assign _T_1365 = _T_1351 == 4'h3; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22843.4]
  assign _T_1366 = _T_1365 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22844.4]
  assign _T_1368 = _T_1351 == 4'h4; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22845.4]
  assign _T_1369 = _T_1368 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22846.4]
  assign _T_1371 = _T_1351 == 4'h5; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22847.4]
  assign _T_1372 = _T_1371 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22848.4]
  assign _T_1374 = _T_1351 == 4'h6; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22849.4]
  assign _T_1375 = _T_1374 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22850.4]
  assign _T_1377 = _T_1351 == 4'h7; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22851.4]
  assign _T_1378 = _T_1377 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22852.4]
  assign _T_1380 = _T_1351 == 4'h8; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22853.4]
  assign _T_1381 = _T_1380 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22854.4]
  assign _T_1383 = _T_1351 == 4'h9; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22855.4]
  assign _T_1384 = _T_1383 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22856.4]
  assign _T_1386 = _T_1351 == 4'ha; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22857.4]
  assign _T_1387 = _T_1386 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22858.4]
  assign _T_1389 = _T_1351 == 4'hb; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22859.4]
  assign _T_1390 = _T_1389 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22860.4]
  assign _T_1392 = _T_1351 == 4'hc; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22861.4]
  assign _T_1393 = _T_1392 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22862.4]
  assign _T_1395 = _T_1351 == 4'hd; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22863.4]
  assign _T_1396 = _T_1395 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22864.4]
  assign _T_1398 = _T_1351 == 4'he; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22865.4]
  assign _T_1399 = _T_1398 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22866.4]
  assign _T_1401 = _T_1351 == 4'hf; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:94:@22867.4]
  assign _T_1402 = _T_1401 & io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 85:102:@22868.4]
  assign _T_1496 = _T_1352 == 4'h0; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22935.4]
  assign _T_1497 = _T_1496 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22936.4]
  assign _T_1499 = _T_1352 == 4'h1; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22937.4]
  assign _T_1500 = _T_1499 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22938.4]
  assign _T_1502 = _T_1352 == 4'h2; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22939.4]
  assign _T_1503 = _T_1502 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22940.4]
  assign _T_1505 = _T_1352 == 4'h3; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22941.4]
  assign _T_1506 = _T_1505 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22942.4]
  assign _T_1508 = _T_1352 == 4'h4; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22943.4]
  assign _T_1509 = _T_1508 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22944.4]
  assign _T_1511 = _T_1352 == 4'h5; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22945.4]
  assign _T_1512 = _T_1511 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22946.4]
  assign _T_1514 = _T_1352 == 4'h6; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22947.4]
  assign _T_1515 = _T_1514 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22948.4]
  assign _T_1517 = _T_1352 == 4'h7; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22949.4]
  assign _T_1518 = _T_1517 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22950.4]
  assign _T_1520 = _T_1352 == 4'h8; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22951.4]
  assign _T_1521 = _T_1520 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22952.4]
  assign _T_1523 = _T_1352 == 4'h9; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22953.4]
  assign _T_1524 = _T_1523 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22954.4]
  assign _T_1526 = _T_1352 == 4'ha; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22955.4]
  assign _T_1527 = _T_1526 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22956.4]
  assign _T_1529 = _T_1352 == 4'hb; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22957.4]
  assign _T_1530 = _T_1529 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22958.4]
  assign _T_1532 = _T_1352 == 4'hc; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22959.4]
  assign _T_1533 = _T_1532 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22960.4]
  assign _T_1535 = _T_1352 == 4'hd; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22961.4]
  assign _T_1536 = _T_1535 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22962.4]
  assign _T_1538 = _T_1352 == 4'he; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22963.4]
  assign _T_1539 = _T_1538 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22964.4]
  assign _T_1541 = _T_1352 == 4'hf; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:96:@22965.4]
  assign _T_1542 = _T_1541 & io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 87:104:@22966.4]
  assign _T_1635 = _T_1357 | _T_1497; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23033.4]
  assign _T_1636 = _T_1360 | _T_1500; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23034.4]
  assign _T_1637 = _T_1363 | _T_1503; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23035.4]
  assign _T_1638 = _T_1366 | _T_1506; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23036.4]
  assign _T_1639 = _T_1369 | _T_1509; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23037.4]
  assign _T_1640 = _T_1372 | _T_1512; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23038.4]
  assign _T_1641 = _T_1375 | _T_1515; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23039.4]
  assign _T_1642 = _T_1378 | _T_1518; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23040.4]
  assign _T_1643 = _T_1381 | _T_1521; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23041.4]
  assign _T_1644 = _T_1384 | _T_1524; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23042.4]
  assign _T_1645 = _T_1387 | _T_1527; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23043.4]
  assign _T_1646 = _T_1390 | _T_1530; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23044.4]
  assign _T_1647 = _T_1393 | _T_1533; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23045.4]
  assign _T_1648 = _T_1396 | _T_1536; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23046.4]
  assign _T_1649 = _T_1399 | _T_1539; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23047.4]
  assign _T_1650 = _T_1402 | _T_1542; // @[NV_NVDLA_CDMA_shared_buffer.scala 90:87:@23048.4]
  assign _T_1752 = _T_1357 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23133.4]
  assign _T_1753 = io_dc2sbuf_p_rd_0_addr_bits[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:86:@23134.4]
  assign _GEN_34 = {{4'd0}, _T_1753}; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23135.4]
  assign _T_1754 = _T_1752 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23135.4]
  assign _T_1765 = _T_1497 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23142.4]
  assign _T_1766 = io_img2sbuf_p_rd_0_addr_bits[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:88:@23143.4]
  assign _GEN_35 = {{4'd0}, _T_1766}; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23144.4]
  assign _T_1767 = _T_1765 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23144.4]
  assign _T_1768 = _T_1754 | _T_1767; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23145.4]
  assign _T_1779 = _T_1360 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23152.4]
  assign _T_1781 = _T_1779 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23154.4]
  assign _T_1792 = _T_1500 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23161.4]
  assign _T_1794 = _T_1792 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23163.4]
  assign _T_1795 = _T_1781 | _T_1794; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23164.4]
  assign _T_1806 = _T_1363 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23171.4]
  assign _T_1808 = _T_1806 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23173.4]
  assign _T_1819 = _T_1503 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23180.4]
  assign _T_1821 = _T_1819 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23182.4]
  assign _T_1822 = _T_1808 | _T_1821; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23183.4]
  assign _T_1833 = _T_1366 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23190.4]
  assign _T_1835 = _T_1833 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23192.4]
  assign _T_1846 = _T_1506 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23199.4]
  assign _T_1848 = _T_1846 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23201.4]
  assign _T_1849 = _T_1835 | _T_1848; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23202.4]
  assign _T_1860 = _T_1369 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23209.4]
  assign _T_1862 = _T_1860 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23211.4]
  assign _T_1873 = _T_1509 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23218.4]
  assign _T_1875 = _T_1873 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23220.4]
  assign _T_1876 = _T_1862 | _T_1875; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23221.4]
  assign _T_1887 = _T_1372 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23228.4]
  assign _T_1889 = _T_1887 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23230.4]
  assign _T_1900 = _T_1512 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23237.4]
  assign _T_1902 = _T_1900 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23239.4]
  assign _T_1903 = _T_1889 | _T_1902; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23240.4]
  assign _T_1914 = _T_1375 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23247.4]
  assign _T_1916 = _T_1914 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23249.4]
  assign _T_1927 = _T_1515 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23256.4]
  assign _T_1929 = _T_1927 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23258.4]
  assign _T_1930 = _T_1916 | _T_1929; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23259.4]
  assign _T_1941 = _T_1378 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23266.4]
  assign _T_1943 = _T_1941 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23268.4]
  assign _T_1954 = _T_1518 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23275.4]
  assign _T_1956 = _T_1954 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23277.4]
  assign _T_1957 = _T_1943 | _T_1956; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23278.4]
  assign _T_1968 = _T_1381 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23285.4]
  assign _T_1970 = _T_1968 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23287.4]
  assign _T_1981 = _T_1521 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23294.4]
  assign _T_1983 = _T_1981 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23296.4]
  assign _T_1984 = _T_1970 | _T_1983; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23297.4]
  assign _T_1995 = _T_1384 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23304.4]
  assign _T_1997 = _T_1995 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23306.4]
  assign _T_2008 = _T_1524 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23313.4]
  assign _T_2010 = _T_2008 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23315.4]
  assign _T_2011 = _T_1997 | _T_2010; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23316.4]
  assign _T_2022 = _T_1387 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23323.4]
  assign _T_2024 = _T_2022 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23325.4]
  assign _T_2035 = _T_1527 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23332.4]
  assign _T_2037 = _T_2035 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23334.4]
  assign _T_2038 = _T_2024 | _T_2037; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23335.4]
  assign _T_2049 = _T_1390 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23342.4]
  assign _T_2051 = _T_2049 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23344.4]
  assign _T_2062 = _T_1530 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23351.4]
  assign _T_2064 = _T_2062 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23353.4]
  assign _T_2065 = _T_2051 | _T_2064; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23354.4]
  assign _T_2076 = _T_1393 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23361.4]
  assign _T_2078 = _T_2076 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23363.4]
  assign _T_2089 = _T_1533 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23370.4]
  assign _T_2091 = _T_2089 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23372.4]
  assign _T_2092 = _T_2078 | _T_2091; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23373.4]
  assign _T_2103 = _T_1396 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23380.4]
  assign _T_2105 = _T_2103 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23382.4]
  assign _T_2116 = _T_1536 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23389.4]
  assign _T_2118 = _T_2116 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23391.4]
  assign _T_2119 = _T_2105 | _T_2118; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23392.4]
  assign _T_2130 = _T_1399 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23399.4]
  assign _T_2132 = _T_2130 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23401.4]
  assign _T_2143 = _T_1539 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23408.4]
  assign _T_2145 = _T_2143 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23410.4]
  assign _T_2146 = _T_2132 | _T_2145; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23411.4]
  assign _T_2157 = _T_1402 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23418.4]
  assign _T_2159 = _T_2157 & _GEN_34; // @[NV_NVDLA_CDMA_shared_buffer.scala 95:57:@23420.4]
  assign _T_2170 = _T_1542 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@23427.4]
  assign _T_2172 = _T_2170 & _GEN_35; // @[NV_NVDLA_CDMA_shared_buffer.scala 97:58:@23429.4]
  assign _T_2173 = _T_2159 | _T_2172; // @[NV_NVDLA_CDMA_shared_buffer.scala 96:96:@23430.4]
  assign _T_2479 = io_dc2sbuf_p_rd_0_addr_valid | io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_CDMA_shared_buffer.scala 127:62:@23682.4]
  assign _T_2490 = _T_2299_0 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23689.4]
  assign _T_2206_0 = nv_ram_rws_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23508.4]
  assign _GEN_66 = {{240'd0}, _T_2490}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23690.4]
  assign _T_2491 = _GEN_66 & _T_2206_0; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23690.4]
  assign _T_2495 = _T_2299_1 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23692.4]
  assign _T_2206_1 = nv_ram_rws_1_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23515.4]
  assign _GEN_67 = {{240'd0}, _T_2495}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23693.4]
  assign _T_2496 = _GEN_67 & _T_2206_1; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23693.4]
  assign _T_2500 = _T_2299_2 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23695.4]
  assign _T_2206_2 = nv_ram_rws_2_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23522.4]
  assign _GEN_68 = {{240'd0}, _T_2500}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23696.4]
  assign _T_2501 = _GEN_68 & _T_2206_2; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23696.4]
  assign _T_2505 = _T_2299_3 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23698.4]
  assign _T_2206_3 = nv_ram_rws_3_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23529.4]
  assign _GEN_69 = {{240'd0}, _T_2505}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23699.4]
  assign _T_2506 = _GEN_69 & _T_2206_3; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23699.4]
  assign _T_2510 = _T_2299_4 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23701.4]
  assign _T_2206_4 = nv_ram_rws_4_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23536.4]
  assign _GEN_70 = {{240'd0}, _T_2510}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23702.4]
  assign _T_2511 = _GEN_70 & _T_2206_4; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23702.4]
  assign _T_2515 = _T_2299_5 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23704.4]
  assign _T_2206_5 = nv_ram_rws_5_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23543.4]
  assign _GEN_71 = {{240'd0}, _T_2515}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23705.4]
  assign _T_2516 = _GEN_71 & _T_2206_5; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23705.4]
  assign _T_2520 = _T_2299_6 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23707.4]
  assign _T_2206_6 = nv_ram_rws_6_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23550.4]
  assign _GEN_72 = {{240'd0}, _T_2520}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23708.4]
  assign _T_2521 = _GEN_72 & _T_2206_6; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23708.4]
  assign _T_2525 = _T_2299_7 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23710.4]
  assign _T_2206_7 = nv_ram_rws_7_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23557.4]
  assign _GEN_73 = {{240'd0}, _T_2525}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23711.4]
  assign _T_2526 = _GEN_73 & _T_2206_7; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23711.4]
  assign _T_2530 = _T_2299_8 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23713.4]
  assign _T_2206_8 = nv_ram_rws_8_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23564.4]
  assign _GEN_74 = {{240'd0}, _T_2530}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23714.4]
  assign _T_2531 = _GEN_74 & _T_2206_8; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23714.4]
  assign _T_2535 = _T_2299_9 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23716.4]
  assign _T_2206_9 = nv_ram_rws_9_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23571.4]
  assign _GEN_75 = {{240'd0}, _T_2535}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23717.4]
  assign _T_2536 = _GEN_75 & _T_2206_9; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23717.4]
  assign _T_2540 = _T_2299_10 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23719.4]
  assign _T_2206_10 = nv_ram_rws_10_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23578.4]
  assign _GEN_76 = {{240'd0}, _T_2540}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23720.4]
  assign _T_2541 = _GEN_76 & _T_2206_10; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23720.4]
  assign _T_2545 = _T_2299_11 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23722.4]
  assign _T_2206_11 = nv_ram_rws_11_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23585.4]
  assign _GEN_77 = {{240'd0}, _T_2545}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23723.4]
  assign _T_2546 = _GEN_77 & _T_2206_11; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23723.4]
  assign _T_2550 = _T_2299_12 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23725.4]
  assign _T_2206_12 = nv_ram_rws_12_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23592.4]
  assign _GEN_78 = {{240'd0}, _T_2550}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23726.4]
  assign _T_2551 = _GEN_78 & _T_2206_12; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23726.4]
  assign _T_2555 = _T_2299_13 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23728.4]
  assign _T_2206_13 = nv_ram_rws_13_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23599.4]
  assign _GEN_79 = {{240'd0}, _T_2555}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23729.4]
  assign _T_2556 = _GEN_79 & _T_2206_13; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23729.4]
  assign _T_2560 = _T_2299_14 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23731.4]
  assign _T_2206_14 = nv_ram_rws_14_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23606.4]
  assign _GEN_80 = {{240'd0}, _T_2560}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23732.4]
  assign _T_2561 = _GEN_80 & _T_2206_14; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23732.4]
  assign _T_2565 = _T_2299_15 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@23734.4]
  assign _T_2206_15 = nv_ram_rws_15_io_dout; // @[NV_NVDLA_CDMA_shared_buffer.scala 106:21:@23501.4 NV_NVDLA_CDMA_shared_buffer.scala 114:18:@23613.4]
  assign _GEN_81 = {{240'd0}, _T_2565}; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23735.4]
  assign _T_2566 = _GEN_81 & _T_2206_15; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:80:@23735.4]
  assign _T_2589 = _T_2491 | _T_2496; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23753.4]
  assign _T_2590 = _T_2589 | _T_2501; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23754.4]
  assign _T_2591 = _T_2590 | _T_2506; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23755.4]
  assign _T_2592 = _T_2591 | _T_2511; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23756.4]
  assign _T_2593 = _T_2592 | _T_2516; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23757.4]
  assign _T_2594 = _T_2593 | _T_2521; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23758.4]
  assign _T_2595 = _T_2594 | _T_2526; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23759.4]
  assign _T_2596 = _T_2595 | _T_2531; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23760.4]
  assign _T_2597 = _T_2596 | _T_2536; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23761.4]
  assign _T_2598 = _T_2597 | _T_2541; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23762.4]
  assign _T_2599 = _T_2598 | _T_2546; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23763.4]
  assign _T_2600 = _T_2599 | _T_2551; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23764.4]
  assign _T_2601 = _T_2600 | _T_2556; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23765.4]
  assign _T_2602 = _T_2601 | _T_2561; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23766.4]
  assign _T_2603 = _T_2602 | _T_2566; // @[NV_NVDLA_CDMA_shared_buffer.scala 135:104:@23767.4]
  assign io_dc2sbuf_p_rd_0_data = _T_2722; // @[NV_NVDLA_CDMA_shared_buffer.scala 144:25:@23856.4]
  assign io_img2sbuf_p_rd_0_data = _T_2722; // @[NV_NVDLA_CDMA_shared_buffer.scala 145:26:@23857.4]
  assign nv_ram_rws_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23502.4]
  assign nv_ram_rws_io_re = _T_1357 | _T_1497; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23504.4]
  assign nv_ram_rws_io_we = _T_159 | _T_299; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23506.4]
  assign nv_ram_rws_io_ra = _T_1768[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23503.4]
  assign nv_ram_rws_io_wa = _T_526[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23505.4]
  assign nv_ram_rws_io_di = _T_965 | _T_976; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23507.4]
  assign nv_ram_rws_1_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23509.4]
  assign nv_ram_rws_1_io_re = _T_1360 | _T_1500; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23511.4]
  assign nv_ram_rws_1_io_we = _T_162 | _T_302; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23513.4]
  assign nv_ram_rws_1_io_ra = _T_1795[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23510.4]
  assign nv_ram_rws_1_io_wa = _T_553[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23512.4]
  assign nv_ram_rws_1_io_di = _T_988 | _T_999; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23514.4]
  assign nv_ram_rws_2_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23516.4]
  assign nv_ram_rws_2_io_re = _T_1363 | _T_1503; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23518.4]
  assign nv_ram_rws_2_io_we = _T_165 | _T_305; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23520.4]
  assign nv_ram_rws_2_io_ra = _T_1822[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23517.4]
  assign nv_ram_rws_2_io_wa = _T_580[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23519.4]
  assign nv_ram_rws_2_io_di = _T_1011 | _T_1022; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23521.4]
  assign nv_ram_rws_3_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23523.4]
  assign nv_ram_rws_3_io_re = _T_1366 | _T_1506; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23525.4]
  assign nv_ram_rws_3_io_we = _T_168 | _T_308; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23527.4]
  assign nv_ram_rws_3_io_ra = _T_1849[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23524.4]
  assign nv_ram_rws_3_io_wa = _T_607[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23526.4]
  assign nv_ram_rws_3_io_di = _T_1034 | _T_1045; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23528.4]
  assign nv_ram_rws_4_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23530.4]
  assign nv_ram_rws_4_io_re = _T_1369 | _T_1509; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23532.4]
  assign nv_ram_rws_4_io_we = _T_171 | _T_311; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23534.4]
  assign nv_ram_rws_4_io_ra = _T_1876[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23531.4]
  assign nv_ram_rws_4_io_wa = _T_634[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23533.4]
  assign nv_ram_rws_4_io_di = _T_1057 | _T_1068; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23535.4]
  assign nv_ram_rws_5_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23537.4]
  assign nv_ram_rws_5_io_re = _T_1372 | _T_1512; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23539.4]
  assign nv_ram_rws_5_io_we = _T_174 | _T_314; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23541.4]
  assign nv_ram_rws_5_io_ra = _T_1903[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23538.4]
  assign nv_ram_rws_5_io_wa = _T_661[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23540.4]
  assign nv_ram_rws_5_io_di = _T_1080 | _T_1091; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23542.4]
  assign nv_ram_rws_6_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23544.4]
  assign nv_ram_rws_6_io_re = _T_1375 | _T_1515; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23546.4]
  assign nv_ram_rws_6_io_we = _T_177 | _T_317; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23548.4]
  assign nv_ram_rws_6_io_ra = _T_1930[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23545.4]
  assign nv_ram_rws_6_io_wa = _T_688[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23547.4]
  assign nv_ram_rws_6_io_di = _T_1103 | _T_1114; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23549.4]
  assign nv_ram_rws_7_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23551.4]
  assign nv_ram_rws_7_io_re = _T_1378 | _T_1518; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23553.4]
  assign nv_ram_rws_7_io_we = _T_180 | _T_320; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23555.4]
  assign nv_ram_rws_7_io_ra = _T_1957[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23552.4]
  assign nv_ram_rws_7_io_wa = _T_715[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23554.4]
  assign nv_ram_rws_7_io_di = _T_1126 | _T_1137; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23556.4]
  assign nv_ram_rws_8_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23558.4]
  assign nv_ram_rws_8_io_re = _T_1381 | _T_1521; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23560.4]
  assign nv_ram_rws_8_io_we = _T_183 | _T_323; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23562.4]
  assign nv_ram_rws_8_io_ra = _T_1984[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23559.4]
  assign nv_ram_rws_8_io_wa = _T_742[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23561.4]
  assign nv_ram_rws_8_io_di = _T_1149 | _T_1160; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23563.4]
  assign nv_ram_rws_9_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23565.4]
  assign nv_ram_rws_9_io_re = _T_1384 | _T_1524; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23567.4]
  assign nv_ram_rws_9_io_we = _T_186 | _T_326; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23569.4]
  assign nv_ram_rws_9_io_ra = _T_2011[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23566.4]
  assign nv_ram_rws_9_io_wa = _T_769[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23568.4]
  assign nv_ram_rws_9_io_di = _T_1172 | _T_1183; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23570.4]
  assign nv_ram_rws_10_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23572.4]
  assign nv_ram_rws_10_io_re = _T_1387 | _T_1527; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23574.4]
  assign nv_ram_rws_10_io_we = _T_189 | _T_329; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23576.4]
  assign nv_ram_rws_10_io_ra = _T_2038[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23573.4]
  assign nv_ram_rws_10_io_wa = _T_796[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23575.4]
  assign nv_ram_rws_10_io_di = _T_1195 | _T_1206; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23577.4]
  assign nv_ram_rws_11_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23579.4]
  assign nv_ram_rws_11_io_re = _T_1390 | _T_1530; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23581.4]
  assign nv_ram_rws_11_io_we = _T_192 | _T_332; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23583.4]
  assign nv_ram_rws_11_io_ra = _T_2065[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23580.4]
  assign nv_ram_rws_11_io_wa = _T_823[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23582.4]
  assign nv_ram_rws_11_io_di = _T_1218 | _T_1229; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23584.4]
  assign nv_ram_rws_12_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23586.4]
  assign nv_ram_rws_12_io_re = _T_1393 | _T_1533; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23588.4]
  assign nv_ram_rws_12_io_we = _T_195 | _T_335; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23590.4]
  assign nv_ram_rws_12_io_ra = _T_2092[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23587.4]
  assign nv_ram_rws_12_io_wa = _T_850[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23589.4]
  assign nv_ram_rws_12_io_di = _T_1241 | _T_1252; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23591.4]
  assign nv_ram_rws_13_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23593.4]
  assign nv_ram_rws_13_io_re = _T_1396 | _T_1536; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23595.4]
  assign nv_ram_rws_13_io_we = _T_198 | _T_338; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23597.4]
  assign nv_ram_rws_13_io_ra = _T_2119[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23594.4]
  assign nv_ram_rws_13_io_wa = _T_877[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23596.4]
  assign nv_ram_rws_13_io_di = _T_1264 | _T_1275; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23598.4]
  assign nv_ram_rws_14_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23600.4]
  assign nv_ram_rws_14_io_re = _T_1399 | _T_1539; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23602.4]
  assign nv_ram_rws_14_io_we = _T_201 | _T_341; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23604.4]
  assign nv_ram_rws_14_io_ra = _T_2146[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23601.4]
  assign nv_ram_rws_14_io_wa = _T_904[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23603.4]
  assign nv_ram_rws_14_io_di = _T_1287 | _T_1298; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23605.4]
  assign nv_ram_rws_15_io_clk = io_nvdla_core_clk; // @[NV_NVDLA_CDMA_shared_buffer.scala 108:31:@23607.4]
  assign nv_ram_rws_15_io_re = _T_1402 | _T_1542; // @[NV_NVDLA_CDMA_shared_buffer.scala 110:30:@23609.4]
  assign nv_ram_rws_15_io_we = _T_204 | _T_344; // @[NV_NVDLA_CDMA_shared_buffer.scala 112:30:@23611.4]
  assign nv_ram_rws_15_io_ra = _T_2173[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 109:30:@23608.4]
  assign nv_ram_rws_15_io_wa = _T_931[3:0]; // @[NV_NVDLA_CDMA_shared_buffer.scala 111:30:@23610.4]
  assign nv_ram_rws_15_io_di = _T_1310 | _T_1321; // @[NV_NVDLA_CDMA_shared_buffer.scala 113:30:@23612.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2299_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2299_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2299_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_2299_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_2299_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_2299_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_2299_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_2299_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_2299_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_2299_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2299_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2299_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_2299_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_2299_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_2299_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_2299_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_2482 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {8{`RANDOM}};
  _T_2722 = _RAND_17[255:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_2299_0 <= 1'h0;
    end else begin
      _T_2299_0 <= _T_1635;
    end
    if (reset) begin
      _T_2299_1 <= 1'h0;
    end else begin
      _T_2299_1 <= _T_1636;
    end
    if (reset) begin
      _T_2299_2 <= 1'h0;
    end else begin
      _T_2299_2 <= _T_1637;
    end
    if (reset) begin
      _T_2299_3 <= 1'h0;
    end else begin
      _T_2299_3 <= _T_1638;
    end
    if (reset) begin
      _T_2299_4 <= 1'h0;
    end else begin
      _T_2299_4 <= _T_1639;
    end
    if (reset) begin
      _T_2299_5 <= 1'h0;
    end else begin
      _T_2299_5 <= _T_1640;
    end
    if (reset) begin
      _T_2299_6 <= 1'h0;
    end else begin
      _T_2299_6 <= _T_1641;
    end
    if (reset) begin
      _T_2299_7 <= 1'h0;
    end else begin
      _T_2299_7 <= _T_1642;
    end
    if (reset) begin
      _T_2299_8 <= 1'h0;
    end else begin
      _T_2299_8 <= _T_1643;
    end
    if (reset) begin
      _T_2299_9 <= 1'h0;
    end else begin
      _T_2299_9 <= _T_1644;
    end
    if (reset) begin
      _T_2299_10 <= 1'h0;
    end else begin
      _T_2299_10 <= _T_1645;
    end
    if (reset) begin
      _T_2299_11 <= 1'h0;
    end else begin
      _T_2299_11 <= _T_1646;
    end
    if (reset) begin
      _T_2299_12 <= 1'h0;
    end else begin
      _T_2299_12 <= _T_1647;
    end
    if (reset) begin
      _T_2299_13 <= 1'h0;
    end else begin
      _T_2299_13 <= _T_1648;
    end
    if (reset) begin
      _T_2299_14 <= 1'h0;
    end else begin
      _T_2299_14 <= _T_1649;
    end
    if (reset) begin
      _T_2299_15 <= 1'h0;
    end else begin
      _T_2299_15 <= _T_1650;
    end
    if (reset) begin
      _T_2482 <= 1'h0;
    end else begin
      _T_2482 <= _T_2479;
    end
    if (_T_2482) begin
      _T_2722 <= _T_2603;
    end
  end
endmodule
module NV_NVDLA_CDMA_status( // @[:@23868.2]
  input         reset, // @[:@23870.4]
  input         io_nvdla_core_clk, // @[:@23871.4]
  input         io_dc2status_dat_updt_valid, // @[:@23871.4]
  input  [14:0] io_dc2status_dat_updt_bits_entries, // @[:@23871.4]
  input  [13:0] io_dc2status_dat_updt_bits_slices, // @[:@23871.4]
  input         io_img2status_dat_updt_valid, // @[:@23871.4]
  input  [14:0] io_img2status_dat_updt_bits_entries, // @[:@23871.4]
  input  [13:0] io_img2status_dat_updt_bits_slices, // @[:@23871.4]
  input         io_sc2cdma_dat_updt_valid, // @[:@23871.4]
  input  [14:0] io_sc2cdma_dat_updt_bits_entries, // @[:@23871.4]
  output        io_cdma2sc_dat_updt_valid, // @[:@23871.4]
  output [14:0] io_cdma2sc_dat_updt_bits_entries, // @[:@23871.4]
  output [13:0] io_cdma2sc_dat_updt_bits_slices, // @[:@23871.4]
  output [14:0] io_status2dma_free_entries, // @[:@23871.4]
  output [14:0] io_status2dma_wr_idx, // @[:@23871.4]
  input  [1:0]  io_dc2status_state, // @[:@23871.4]
  input  [1:0]  io_img2status_state, // @[:@23871.4]
  input  [1:0]  io_wt2status_state, // @[:@23871.4]
  input         io_dp2reg_consumer, // @[:@23871.4]
  output        io_dp2reg_done, // @[:@23871.4]
  input         io_reg2dp_op_en, // @[:@23871.4]
  input  [4:0]  io_reg2dp_data_bank, // @[:@23871.4]
  output [1:0]  io_cdma_wt2glb_done_intr_pd, // @[:@23871.4]
  output [1:0]  io_cdma_dat2glb_done_intr_pd, // @[:@23871.4]
  input  [1:0]  io_sc2cdma_dat_pending_req, // @[:@23871.4]
  output [1:0]  io_cdma2sc_dat_pending_ack, // @[:@23871.4]
  output        io_status2dma_fsm_switch // @[:@23871.4]
);
  reg  _T_111; // @[NV_NVDLA_CDMA_status.scala 72:44:@23873.4]
  reg [31:0] _RAND_0;
  reg  _T_114; // @[NV_NVDLA_CDMA_status.scala 73:36:@23874.4]
  reg [31:0] _RAND_1;
  reg  _T_117; // @[NV_NVDLA_CDMA_status.scala 74:37:@23875.4]
  reg [31:0] _RAND_2;
  reg [1:0] _T_120; // @[NV_NVDLA_CDMA_status.scala 75:31:@23876.4]
  reg [31:0] _RAND_3;
  reg [1:0] _T_123; // @[NV_NVDLA_CDMA_status.scala 76:32:@23877.4]
  reg [31:0] _RAND_4;
  wire  _T_125; // @[NV_NVDLA_CDMA_status.scala 78:46:@23878.4]
  wire  _T_127; // @[NV_NVDLA_CDMA_status.scala 79:46:@23879.4]
  wire  _T_129; // @[NV_NVDLA_CDMA_status.scala 80:46:@23880.4]
  wire  _T_131; // @[NV_NVDLA_CDMA_status.scala 81:48:@23881.4]
  wire  _T_133; // @[NV_NVDLA_CDMA_status.scala 82:48:@23882.4]
  wire  _T_134; // @[NV_NVDLA_CDMA_status.scala 83:43:@23883.4]
  wire  _T_135; // @[NV_NVDLA_CDMA_status.scala 84:53:@23884.4]
  wire  _T_136; // @[NV_NVDLA_CDMA_status.scala 84:51:@23885.4]
  wire  _T_137; // @[NV_NVDLA_CDMA_status.scala 84:80:@23886.4]
  wire  _T_138; // @[NV_NVDLA_CDMA_status.scala 84:97:@23887.4]
  wire  _T_139; // @[NV_NVDLA_CDMA_status.scala 86:46:@23888.4]
  wire  _T_140; // @[NV_NVDLA_CDMA_status.scala 86:69:@23889.4]
  wire  _T_141; // @[NV_NVDLA_CDMA_status.scala 86:67:@23890.4]
  wire  _T_142; // @[NV_NVDLA_CDMA_status.scala 86:88:@23891.4]
  wire  _T_143; // @[NV_NVDLA_CDMA_status.scala 87:48:@23892.4]
  wire  _T_144; // @[NV_NVDLA_CDMA_status.scala 87:46:@23893.4]
  wire  _T_146; // @[NV_NVDLA_CDMA_status.scala 87:68:@23895.4]
  wire  _T_147; // @[NV_NVDLA_CDMA_status.scala 87:89:@23896.4]
  wire [1:0] _T_148; // @[Cat.scala 30:58:@23897.4]
  wire  _T_150; // @[NV_NVDLA_CDMA_status.scala 89:70:@23899.4]
  wire  _T_151; // @[NV_NVDLA_CDMA_status.scala 89:68:@23900.4]
  wire  _T_152; // @[NV_NVDLA_CDMA_status.scala 89:90:@23901.4]
  wire  _T_156; // @[NV_NVDLA_CDMA_status.scala 90:68:@23905.4]
  wire  _T_157; // @[NV_NVDLA_CDMA_status.scala 90:90:@23906.4]
  wire [1:0] _T_158; // @[Cat.scala 30:58:@23907.4]
  wire  _T_159; // @[NV_NVDLA_CDMA_status.scala 93:42:@23909.4]
  wire  _T_160; // @[NV_NVDLA_CDMA_status.scala 94:43:@23911.4]
  reg [14:0] _T_166; // @[NV_NVDLA_CDMA_status.scala 107:43:@23920.4]
  reg [31:0] _RAND_5;
  reg [14:0] _T_172; // @[NV_NVDLA_CDMA_status.scala 109:46:@23922.4]
  reg [31:0] _RAND_6;
  reg [14:0] _T_175; // @[NV_NVDLA_CDMA_status.scala 110:40:@23923.4]
  reg [31:0] _RAND_7;
  reg [5:0] _T_178; // @[NV_NVDLA_CDMA_status.scala 111:28:@23924.4]
  reg [31:0] _RAND_8;
  reg  _T_181; // @[NV_NVDLA_CDMA_status.scala 112:30:@23925.4]
  reg [31:0] _RAND_9;
  reg  _T_184; // @[NV_NVDLA_CDMA_status.scala 113:30:@23926.4]
  reg [31:0] _RAND_10;
  wire [5:0] _T_190; // @[NV_NVDLA_CDMA_status.scala 118:43:@23929.4]
  wire  _T_191; // @[NV_NVDLA_CDMA_status.scala 119:60:@23930.4]
  wire  _T_192; // @[NV_NVDLA_CDMA_status.scala 119:44:@23931.4]
  wire  _T_193; // @[NV_NVDLA_CDMA_status.scala 122:60:@23932.4]
  wire  _T_194; // @[NV_NVDLA_CDMA_status.scala 122:42:@23933.4]
  wire  _T_195; // @[NV_NVDLA_CDMA_status.scala 123:50:@23934.4]
  wire  _T_196; // @[NV_NVDLA_CDMA_status.scala 124:33:@23935.4]
  wire  _T_197; // @[NV_NVDLA_CDMA_status.scala 124:76:@23936.4]
  wire  _T_198; // @[NV_NVDLA_CDMA_status.scala 124:61:@23937.4]
  wire [14:0] _T_202; // @[Bitwise.scala 72:12:@23939.4]
  wire [14:0] _T_203; // @[NV_NVDLA_CDMA_status.scala 125:62:@23940.4]
  wire [14:0] _T_207; // @[Bitwise.scala 72:12:@23942.4]
  wire [14:0] _T_208; // @[NV_NVDLA_CDMA_status.scala 126:63:@23943.4]
  wire [14:0] _T_209; // @[NV_NVDLA_CDMA_status.scala 125:99:@23944.4]
  wire [14:0] _T_211; // @[NV_NVDLA_CDMA_status.scala 127:26:@23945.4]
  wire [15:0] _T_214; // @[NV_NVDLA_CDMA_status.scala 128:113:@23947.4]
  wire [14:0] _T_215; // @[NV_NVDLA_CDMA_status.scala 128:113:@23948.4]
  wire [15:0] _T_216; // @[NV_NVDLA_CDMA_status.scala 128:127:@23949.4]
  wire [15:0] _T_217; // @[NV_NVDLA_CDMA_status.scala 128:127:@23950.4]
  wire [14:0] _T_218; // @[NV_NVDLA_CDMA_status.scala 128:127:@23951.4]
  wire [14:0] _T_219; // @[NV_NVDLA_CDMA_status.scala 128:41:@23952.4]
  wire [13:0] _T_223; // @[Bitwise.scala 72:12:@23954.4]
  wire [13:0] _T_224; // @[NV_NVDLA_CDMA_status.scala 129:61:@23955.4]
  wire [13:0] _T_228; // @[Bitwise.scala 72:12:@23957.4]
  wire [13:0] _T_229; // @[NV_NVDLA_CDMA_status.scala 130:62:@23958.4]
  wire [13:0] _T_230; // @[NV_NVDLA_CDMA_status.scala 129:97:@23959.4]
  wire [14:0] _T_242; // @[Cat.scala 30:58:@23968.4]
  wire [15:0] _T_243; // @[NV_NVDLA_CDMA_status.scala 133:105:@23969.4]
  wire [15:0] _T_244; // @[NV_NVDLA_CDMA_status.scala 133:105:@23970.4]
  wire [14:0] _T_245; // @[NV_NVDLA_CDMA_status.scala 133:105:@23971.4]
  wire  _T_246; // @[NV_NVDLA_CDMA_status.scala 134:53:@23972.4]
  wire [15:0] _T_247; // @[NV_NVDLA_CDMA_status.scala 135:55:@23973.4]
  wire [14:0] _T_248; // @[NV_NVDLA_CDMA_status.scala 135:55:@23974.4]
  wire [15:0] _T_253; // @[NV_NVDLA_CDMA_status.scala 136:74:@23978.4]
  wire [15:0] _T_254; // @[NV_NVDLA_CDMA_status.scala 136:74:@23979.4]
  wire [14:0] _T_255; // @[NV_NVDLA_CDMA_status.scala 136:74:@23980.4]
  wire  _T_258; // @[NV_NVDLA_CDMA_status.scala 137:61:@23982.4]
  wire  _T_261; // @[NV_NVDLA_CDMA_status.scala 139:35:@23984.4]
  wire [14:0] _T_262; // @[NV_NVDLA_CDMA_status.scala 140:34:@23985.4]
  wire [14:0] _T_263; // @[NV_NVDLA_CDMA_status.scala 139:34:@23986.4]
  wire [14:0] _T_264; // @[NV_NVDLA_CDMA_status.scala 138:34:@23987.4]
  wire [14:0] _GEN_0; // @[NV_NVDLA_CDMA_status.scala 144:21:@23989.4]
  wire [14:0] _GEN_2; // @[NV_NVDLA_CDMA_status.scala 144:21:@23989.4]
  wire [14:0] _GEN_3; // @[NV_NVDLA_CDMA_status.scala 149:25:@23994.4]
  wire [5:0] _GEN_4; // @[NV_NVDLA_CDMA_status.scala 152:27:@23997.4]
  reg  _T_269; // @[NV_NVDLA_CDMA_status.scala 164:64:@24007.4]
  reg [31:0] _RAND_11;
  reg  _T_272; // @[NV_NVDLA_CDMA_status.scala 164:64:@24008.4]
  reg [31:0] _RAND_12;
  reg  _T_275; // @[NV_NVDLA_CDMA_status.scala 164:64:@24009.4]
  reg [31:0] _RAND_13;
  reg  _T_278; // @[NV_NVDLA_CDMA_status.scala 164:64:@24010.4]
  reg [31:0] _RAND_14;
  reg  _T_281; // @[NV_NVDLA_CDMA_status.scala 164:64:@24011.4]
  reg [31:0] _RAND_15;
  reg  _T_284; // @[NV_NVDLA_CDMA_status.scala 164:64:@24012.4]
  reg [31:0] _RAND_16;
  reg  _T_287; // @[NV_NVDLA_CDMA_status.scala 164:64:@24013.4]
  reg [31:0] _RAND_17;
  reg  _T_290; // @[NV_NVDLA_CDMA_status.scala 164:64:@24014.4]
  reg [31:0] _RAND_18;
  reg  _T_293; // @[NV_NVDLA_CDMA_status.scala 164:64:@24015.4]
  reg [31:0] _RAND_19;
  reg [14:0] _T_298; // @[NV_NVDLA_CDMA_status.scala 166:67:@24017.4]
  reg [31:0] _RAND_20;
  reg [14:0] _T_301; // @[NV_NVDLA_CDMA_status.scala 166:67:@24018.4]
  reg [31:0] _RAND_21;
  reg [14:0] _T_304; // @[NV_NVDLA_CDMA_status.scala 166:67:@24019.4]
  reg [31:0] _RAND_22;
  reg [14:0] _T_307; // @[NV_NVDLA_CDMA_status.scala 166:67:@24020.4]
  reg [31:0] _RAND_23;
  reg [14:0] _T_310; // @[NV_NVDLA_CDMA_status.scala 166:67:@24021.4]
  reg [31:0] _RAND_24;
  reg [14:0] _T_313; // @[NV_NVDLA_CDMA_status.scala 166:67:@24022.4]
  reg [31:0] _RAND_25;
  reg [14:0] _T_316; // @[NV_NVDLA_CDMA_status.scala 166:67:@24023.4]
  reg [31:0] _RAND_26;
  reg [14:0] _T_319; // @[NV_NVDLA_CDMA_status.scala 166:67:@24024.4]
  reg [31:0] _RAND_27;
  reg [14:0] _T_322; // @[NV_NVDLA_CDMA_status.scala 166:67:@24025.4]
  reg [31:0] _RAND_28;
  reg [13:0] _T_327; // @[NV_NVDLA_CDMA_status.scala 168:66:@24027.4]
  reg [31:0] _RAND_29;
  reg [13:0] _T_330; // @[NV_NVDLA_CDMA_status.scala 168:66:@24028.4]
  reg [31:0] _RAND_30;
  reg [13:0] _T_333; // @[NV_NVDLA_CDMA_status.scala 168:66:@24029.4]
  reg [31:0] _RAND_31;
  reg [13:0] _T_336; // @[NV_NVDLA_CDMA_status.scala 168:66:@24030.4]
  reg [31:0] _RAND_32;
  reg [13:0] _T_339; // @[NV_NVDLA_CDMA_status.scala 168:66:@24031.4]
  reg [31:0] _RAND_33;
  reg [13:0] _T_342; // @[NV_NVDLA_CDMA_status.scala 168:66:@24032.4]
  reg [31:0] _RAND_34;
  reg [13:0] _T_345; // @[NV_NVDLA_CDMA_status.scala 168:66:@24033.4]
  reg [31:0] _RAND_35;
  reg [13:0] _T_348; // @[NV_NVDLA_CDMA_status.scala 168:66:@24034.4]
  reg [31:0] _RAND_36;
  reg [13:0] _T_351; // @[NV_NVDLA_CDMA_status.scala 168:66:@24035.4]
  reg [31:0] _RAND_37;
  wire [14:0] _GEN_5; // @[NV_NVDLA_CDMA_status.scala 175:28:@24040.4]
  wire [13:0] _GEN_6; // @[NV_NVDLA_CDMA_status.scala 175:28:@24040.4]
  wire [14:0] _GEN_7; // @[NV_NVDLA_CDMA_status.scala 175:28:@24045.4]
  wire [13:0] _GEN_8; // @[NV_NVDLA_CDMA_status.scala 175:28:@24045.4]
  wire [14:0] _GEN_9; // @[NV_NVDLA_CDMA_status.scala 175:28:@24050.4]
  wire [13:0] _GEN_10; // @[NV_NVDLA_CDMA_status.scala 175:28:@24050.4]
  wire [14:0] _GEN_11; // @[NV_NVDLA_CDMA_status.scala 175:28:@24055.4]
  wire [13:0] _GEN_12; // @[NV_NVDLA_CDMA_status.scala 175:28:@24055.4]
  wire [14:0] _GEN_13; // @[NV_NVDLA_CDMA_status.scala 175:28:@24060.4]
  wire [13:0] _GEN_14; // @[NV_NVDLA_CDMA_status.scala 175:28:@24060.4]
  wire [14:0] _GEN_15; // @[NV_NVDLA_CDMA_status.scala 175:28:@24065.4]
  wire [13:0] _GEN_16; // @[NV_NVDLA_CDMA_status.scala 175:28:@24065.4]
  wire [14:0] _GEN_17; // @[NV_NVDLA_CDMA_status.scala 175:28:@24070.4]
  wire [13:0] _GEN_18; // @[NV_NVDLA_CDMA_status.scala 175:28:@24070.4]
  wire [14:0] _GEN_19; // @[NV_NVDLA_CDMA_status.scala 175:28:@24075.4]
  wire [13:0] _GEN_20; // @[NV_NVDLA_CDMA_status.scala 175:28:@24075.4]
  wire [14:0] _GEN_21; // @[NV_NVDLA_CDMA_status.scala 175:28:@24080.4]
  wire [13:0] _GEN_22; // @[NV_NVDLA_CDMA_status.scala 175:28:@24080.4]
  assign _T_125 = io_wt2status_state == 2'h3; // @[NV_NVDLA_CDMA_status.scala 78:46:@23878.4]
  assign _T_127 = io_dc2status_state == 2'h3; // @[NV_NVDLA_CDMA_status.scala 79:46:@23879.4]
  assign _T_129 = io_dc2status_state == 2'h1; // @[NV_NVDLA_CDMA_status.scala 80:46:@23880.4]
  assign _T_131 = io_img2status_state == 2'h3; // @[NV_NVDLA_CDMA_status.scala 81:48:@23881.4]
  assign _T_133 = io_img2status_state == 2'h1; // @[NV_NVDLA_CDMA_status.scala 82:48:@23882.4]
  assign _T_134 = _T_127 | _T_131; // @[NV_NVDLA_CDMA_status.scala 83:43:@23883.4]
  assign _T_135 = ~ _T_111; // @[NV_NVDLA_CDMA_status.scala 84:53:@23884.4]
  assign _T_136 = io_reg2dp_op_en & _T_135; // @[NV_NVDLA_CDMA_status.scala 84:51:@23885.4]
  assign _T_137 = _T_136 & _T_125; // @[NV_NVDLA_CDMA_status.scala 84:80:@23886.4]
  assign _T_138 = _T_137 & _T_134; // @[NV_NVDLA_CDMA_status.scala 84:97:@23887.4]
  assign _T_139 = io_reg2dp_op_en & io_dp2reg_consumer; // @[NV_NVDLA_CDMA_status.scala 86:46:@23888.4]
  assign _T_140 = ~ _T_114; // @[NV_NVDLA_CDMA_status.scala 86:69:@23889.4]
  assign _T_141 = _T_139 & _T_140; // @[NV_NVDLA_CDMA_status.scala 86:67:@23890.4]
  assign _T_142 = _T_141 & _T_125; // @[NV_NVDLA_CDMA_status.scala 86:88:@23891.4]
  assign _T_143 = ~ io_dp2reg_consumer; // @[NV_NVDLA_CDMA_status.scala 87:48:@23892.4]
  assign _T_144 = io_reg2dp_op_en & _T_143; // @[NV_NVDLA_CDMA_status.scala 87:46:@23893.4]
  assign _T_146 = _T_144 & _T_140; // @[NV_NVDLA_CDMA_status.scala 87:68:@23895.4]
  assign _T_147 = _T_146 & _T_125; // @[NV_NVDLA_CDMA_status.scala 87:89:@23896.4]
  assign _T_148 = {_T_142,_T_147}; // @[Cat.scala 30:58:@23897.4]
  assign _T_150 = ~ _T_117; // @[NV_NVDLA_CDMA_status.scala 89:70:@23899.4]
  assign _T_151 = _T_139 & _T_150; // @[NV_NVDLA_CDMA_status.scala 89:68:@23900.4]
  assign _T_152 = _T_151 & _T_134; // @[NV_NVDLA_CDMA_status.scala 89:90:@23901.4]
  assign _T_156 = _T_144 & _T_150; // @[NV_NVDLA_CDMA_status.scala 90:68:@23905.4]
  assign _T_157 = _T_156 & _T_134; // @[NV_NVDLA_CDMA_status.scala 90:90:@23906.4]
  assign _T_158 = {_T_152,_T_157}; // @[Cat.scala 30:58:@23907.4]
  assign _T_159 = io_reg2dp_op_en & _T_125; // @[NV_NVDLA_CDMA_status.scala 93:42:@23909.4]
  assign _T_160 = io_reg2dp_op_en & _T_134; // @[NV_NVDLA_CDMA_status.scala 94:43:@23911.4]
  assign _T_190 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CDMA_status.scala 118:43:@23929.4]
  assign _T_191 = _T_190 != _T_178; // @[NV_NVDLA_CDMA_status.scala 119:60:@23930.4]
  assign _T_192 = io_reg2dp_op_en & _T_191; // @[NV_NVDLA_CDMA_status.scala 119:44:@23931.4]
  assign _T_193 = _T_129 | _T_133; // @[NV_NVDLA_CDMA_status.scala 122:60:@23932.4]
  assign _T_194 = io_reg2dp_op_en & _T_193; // @[NV_NVDLA_CDMA_status.scala 122:42:@23933.4]
  assign _T_195 = io_dc2status_dat_updt_valid | io_img2status_dat_updt_valid; // @[NV_NVDLA_CDMA_status.scala 123:50:@23934.4]
  assign _T_196 = _T_195 | io_sc2cdma_dat_updt_valid; // @[NV_NVDLA_CDMA_status.scala 124:33:@23935.4]
  assign _T_197 = _T_181 & _T_184; // @[NV_NVDLA_CDMA_status.scala 124:76:@23936.4]
  assign _T_198 = _T_196 | _T_197; // @[NV_NVDLA_CDMA_status.scala 124:61:@23937.4]
  assign _T_202 = io_dc2status_dat_updt_valid ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12:@23939.4]
  assign _T_203 = _T_202 & io_dc2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_status.scala 125:62:@23940.4]
  assign _T_207 = io_img2status_dat_updt_valid ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12:@23942.4]
  assign _T_208 = _T_207 & io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_CDMA_status.scala 126:63:@23943.4]
  assign _T_209 = _T_203 | _T_208; // @[NV_NVDLA_CDMA_status.scala 125:99:@23944.4]
  assign _T_211 = io_sc2cdma_dat_updt_valid ? io_sc2cdma_dat_updt_bits_entries : 15'h0; // @[NV_NVDLA_CDMA_status.scala 127:26:@23945.4]
  assign _T_214 = _T_166 + _T_209; // @[NV_NVDLA_CDMA_status.scala 128:113:@23947.4]
  assign _T_215 = _T_166 + _T_209; // @[NV_NVDLA_CDMA_status.scala 128:113:@23948.4]
  assign _T_216 = _T_215 - _T_211; // @[NV_NVDLA_CDMA_status.scala 128:127:@23949.4]
  assign _T_217 = $unsigned(_T_216); // @[NV_NVDLA_CDMA_status.scala 128:127:@23950.4]
  assign _T_218 = _T_217[14:0]; // @[NV_NVDLA_CDMA_status.scala 128:127:@23951.4]
  assign _T_219 = _T_197 ? 15'h0 : _T_218; // @[NV_NVDLA_CDMA_status.scala 128:41:@23952.4]
  assign _T_223 = io_dc2status_dat_updt_valid ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12:@23954.4]
  assign _T_224 = _T_223 & io_dc2status_dat_updt_bits_slices; // @[NV_NVDLA_CDMA_status.scala 129:61:@23955.4]
  assign _T_228 = io_img2status_dat_updt_valid ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12:@23957.4]
  assign _T_229 = _T_228 & io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_CDMA_status.scala 130:62:@23958.4]
  assign _T_230 = _T_224 | _T_229; // @[NV_NVDLA_CDMA_status.scala 129:97:@23959.4]
  assign _T_242 = {_T_178,9'h0}; // @[Cat.scala 30:58:@23968.4]
  assign _T_243 = _T_242 - _T_219; // @[NV_NVDLA_CDMA_status.scala 133:105:@23969.4]
  assign _T_244 = $unsigned(_T_243); // @[NV_NVDLA_CDMA_status.scala 133:105:@23970.4]
  assign _T_245 = _T_244[14:0]; // @[NV_NVDLA_CDMA_status.scala 133:105:@23971.4]
  assign _T_246 = _T_245 != _T_172; // @[NV_NVDLA_CDMA_status.scala 134:53:@23972.4]
  assign _T_247 = _T_175 + _T_209; // @[NV_NVDLA_CDMA_status.scala 135:55:@23973.4]
  assign _T_248 = _T_175 + _T_209; // @[NV_NVDLA_CDMA_status.scala 135:55:@23974.4]
  assign _T_253 = _T_248 - _T_242; // @[NV_NVDLA_CDMA_status.scala 136:74:@23978.4]
  assign _T_254 = $unsigned(_T_253); // @[NV_NVDLA_CDMA_status.scala 136:74:@23979.4]
  assign _T_255 = _T_254[14:0]; // @[NV_NVDLA_CDMA_status.scala 136:74:@23980.4]
  assign _T_258 = _T_248 >= _T_242; // @[NV_NVDLA_CDMA_status.scala 137:61:@23982.4]
  assign _T_261 = ~ _T_195; // @[NV_NVDLA_CDMA_status.scala 139:35:@23984.4]
  assign _T_262 = _T_258 ? _T_255 : _T_248; // @[NV_NVDLA_CDMA_status.scala 140:34:@23985.4]
  assign _T_263 = _T_261 ? _T_175 : _T_262; // @[NV_NVDLA_CDMA_status.scala 139:34:@23986.4]
  assign _T_264 = _T_197 ? 15'h0 : _T_263; // @[NV_NVDLA_CDMA_status.scala 138:34:@23987.4]
  assign _GEN_0 = _T_198 ? _T_219 : _T_166; // @[NV_NVDLA_CDMA_status.scala 144:21:@23989.4]
  assign _GEN_2 = _T_198 ? _T_264 : _T_175; // @[NV_NVDLA_CDMA_status.scala 144:21:@23989.4]
  assign _GEN_3 = _T_246 ? _T_245 : _T_172; // @[NV_NVDLA_CDMA_status.scala 149:25:@23994.4]
  assign _GEN_4 = _T_192 ? _T_190 : _T_178; // @[NV_NVDLA_CDMA_status.scala 152:27:@23997.4]
  assign _GEN_5 = _T_195 ? _T_209 : _T_298; // @[NV_NVDLA_CDMA_status.scala 175:28:@24040.4]
  assign _GEN_6 = _T_195 ? _T_230 : _T_327; // @[NV_NVDLA_CDMA_status.scala 175:28:@24040.4]
  assign _GEN_7 = _T_269 ? _T_298 : _T_301; // @[NV_NVDLA_CDMA_status.scala 175:28:@24045.4]
  assign _GEN_8 = _T_269 ? _T_327 : _T_330; // @[NV_NVDLA_CDMA_status.scala 175:28:@24045.4]
  assign _GEN_9 = _T_272 ? _T_301 : _T_304; // @[NV_NVDLA_CDMA_status.scala 175:28:@24050.4]
  assign _GEN_10 = _T_272 ? _T_330 : _T_333; // @[NV_NVDLA_CDMA_status.scala 175:28:@24050.4]
  assign _GEN_11 = _T_275 ? _T_304 : _T_307; // @[NV_NVDLA_CDMA_status.scala 175:28:@24055.4]
  assign _GEN_12 = _T_275 ? _T_333 : _T_336; // @[NV_NVDLA_CDMA_status.scala 175:28:@24055.4]
  assign _GEN_13 = _T_278 ? _T_307 : _T_310; // @[NV_NVDLA_CDMA_status.scala 175:28:@24060.4]
  assign _GEN_14 = _T_278 ? _T_336 : _T_339; // @[NV_NVDLA_CDMA_status.scala 175:28:@24060.4]
  assign _GEN_15 = _T_281 ? _T_310 : _T_313; // @[NV_NVDLA_CDMA_status.scala 175:28:@24065.4]
  assign _GEN_16 = _T_281 ? _T_339 : _T_342; // @[NV_NVDLA_CDMA_status.scala 175:28:@24065.4]
  assign _GEN_17 = _T_284 ? _T_313 : _T_316; // @[NV_NVDLA_CDMA_status.scala 175:28:@24070.4]
  assign _GEN_18 = _T_284 ? _T_342 : _T_345; // @[NV_NVDLA_CDMA_status.scala 175:28:@24070.4]
  assign _GEN_19 = _T_287 ? _T_316 : _T_319; // @[NV_NVDLA_CDMA_status.scala 175:28:@24075.4]
  assign _GEN_20 = _T_287 ? _T_345 : _T_348; // @[NV_NVDLA_CDMA_status.scala 175:28:@24075.4]
  assign _GEN_21 = _T_290 ? _T_319 : _T_322; // @[NV_NVDLA_CDMA_status.scala 175:28:@24080.4]
  assign _GEN_22 = _T_290 ? _T_348 : _T_351; // @[NV_NVDLA_CDMA_status.scala 175:28:@24080.4]
  assign io_cdma2sc_dat_updt_valid = _T_293; // @[NV_NVDLA_CDMA_status.scala 181:31:@24084.4]
  assign io_cdma2sc_dat_updt_bits_entries = _T_322; // @[NV_NVDLA_CDMA_status.scala 182:38:@24085.4]
  assign io_cdma2sc_dat_updt_bits_slices = _T_351; // @[NV_NVDLA_CDMA_status.scala 183:37:@24086.4]
  assign io_status2dma_free_entries = _T_172; // @[NV_NVDLA_CDMA_status.scala 159:32:@24003.4]
  assign io_status2dma_wr_idx = _T_175; // @[NV_NVDLA_CDMA_status.scala 161:26:@24005.4]
  assign io_dp2reg_done = io_status2dma_fsm_switch; // @[NV_NVDLA_CDMA_status.scala 99:20:@23916.4]
  assign io_cdma_wt2glb_done_intr_pd = _T_120; // @[NV_NVDLA_CDMA_status.scala 100:33:@23917.4]
  assign io_cdma_dat2glb_done_intr_pd = _T_123; // @[NV_NVDLA_CDMA_status.scala 101:34:@23918.4]
  assign io_cdma2sc_dat_pending_ack = {{1'd0}, _T_181}; // @[NV_NVDLA_CDMA_status.scala 157:32:@24002.4]
  assign io_status2dma_fsm_switch = _T_111; // @[NV_NVDLA_CDMA_status.scala 98:30:@23915.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_111 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_114 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_117 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_120 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_123 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_166 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_172 = _RAND_6[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_175 = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_178 = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_181 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_184 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_269 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_272 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_275 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_278 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_281 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_284 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_287 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_290 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_293 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_298 = _RAND_20[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_301 = _RAND_21[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_304 = _RAND_22[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_307 = _RAND_23[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_310 = _RAND_24[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_313 = _RAND_25[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_316 = _RAND_26[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_319 = _RAND_27[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_322 = _RAND_28[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_327 = _RAND_29[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_330 = _RAND_30[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_333 = _RAND_31[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_336 = _RAND_32[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_339 = _RAND_33[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_342 = _RAND_34[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_345 = _RAND_35[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_348 = _RAND_36[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_351 = _RAND_37[13:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_111 <= 1'h0;
    end else begin
      _T_111 <= _T_138;
    end
    if (reset) begin
      _T_114 <= 1'h0;
    end else begin
      _T_114 <= _T_159;
    end
    if (reset) begin
      _T_117 <= 1'h0;
    end else begin
      _T_117 <= _T_160;
    end
    if (reset) begin
      _T_120 <= 2'h0;
    end else begin
      _T_120 <= _T_148;
    end
    if (reset) begin
      _T_123 <= 2'h0;
    end else begin
      _T_123 <= _T_158;
    end
    if (reset) begin
      _T_166 <= 15'h0;
    end else begin
      if (_T_198) begin
        if (_T_197) begin
          _T_166 <= 15'h0;
        end else begin
          _T_166 <= _T_218;
        end
      end
    end
    if (reset) begin
      _T_172 <= 15'h0;
    end else begin
      if (_T_246) begin
        _T_172 <= _T_245;
      end
    end
    if (reset) begin
      _T_175 <= 15'h0;
    end else begin
      if (_T_198) begin
        if (_T_197) begin
          _T_175 <= 15'h0;
        end else begin
          if (!(_T_261)) begin
            if (_T_258) begin
              _T_175 <= _T_255;
            end else begin
              _T_175 <= _T_248;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_178 <= 6'h0;
    end else begin
      if (_T_192) begin
        _T_178 <= _T_190;
      end
    end
    if (reset) begin
      _T_181 <= 1'h0;
    end else begin
      _T_181 <= _T_194;
    end
    if (reset) begin
      _T_184 <= 1'h0;
    end else begin
      _T_184 <= io_sc2cdma_dat_pending_req[0];
    end
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_195;
    end
    if (reset) begin
      _T_272 <= 1'h0;
    end else begin
      _T_272 <= _T_269;
    end
    if (reset) begin
      _T_275 <= 1'h0;
    end else begin
      _T_275 <= _T_272;
    end
    if (reset) begin
      _T_278 <= 1'h0;
    end else begin
      _T_278 <= _T_275;
    end
    if (reset) begin
      _T_281 <= 1'h0;
    end else begin
      _T_281 <= _T_278;
    end
    if (reset) begin
      _T_284 <= 1'h0;
    end else begin
      _T_284 <= _T_281;
    end
    if (reset) begin
      _T_287 <= 1'h0;
    end else begin
      _T_287 <= _T_284;
    end
    if (reset) begin
      _T_290 <= 1'h0;
    end else begin
      _T_290 <= _T_287;
    end
    if (reset) begin
      _T_293 <= 1'h0;
    end else begin
      _T_293 <= _T_290;
    end
    if (reset) begin
      _T_298 <= 15'h0;
    end else begin
      if (_T_195) begin
        _T_298 <= _T_209;
      end
    end
    if (reset) begin
      _T_301 <= 15'h0;
    end else begin
      if (_T_269) begin
        _T_301 <= _T_298;
      end
    end
    if (reset) begin
      _T_304 <= 15'h0;
    end else begin
      if (_T_272) begin
        _T_304 <= _T_301;
      end
    end
    if (reset) begin
      _T_307 <= 15'h0;
    end else begin
      if (_T_275) begin
        _T_307 <= _T_304;
      end
    end
    if (reset) begin
      _T_310 <= 15'h0;
    end else begin
      if (_T_278) begin
        _T_310 <= _T_307;
      end
    end
    if (reset) begin
      _T_313 <= 15'h0;
    end else begin
      if (_T_281) begin
        _T_313 <= _T_310;
      end
    end
    if (reset) begin
      _T_316 <= 15'h0;
    end else begin
      if (_T_284) begin
        _T_316 <= _T_313;
      end
    end
    if (reset) begin
      _T_319 <= 15'h0;
    end else begin
      if (_T_287) begin
        _T_319 <= _T_316;
      end
    end
    if (reset) begin
      _T_322 <= 15'h0;
    end else begin
      if (_T_290) begin
        _T_322 <= _T_319;
      end
    end
    if (reset) begin
      _T_327 <= 14'h0;
    end else begin
      if (_T_195) begin
        _T_327 <= _T_230;
      end
    end
    if (reset) begin
      _T_330 <= 14'h0;
    end else begin
      if (_T_269) begin
        _T_330 <= _T_327;
      end
    end
    if (reset) begin
      _T_333 <= 14'h0;
    end else begin
      if (_T_272) begin
        _T_333 <= _T_330;
      end
    end
    if (reset) begin
      _T_336 <= 14'h0;
    end else begin
      if (_T_275) begin
        _T_336 <= _T_333;
      end
    end
    if (reset) begin
      _T_339 <= 14'h0;
    end else begin
      if (_T_278) begin
        _T_339 <= _T_336;
      end
    end
    if (reset) begin
      _T_342 <= 14'h0;
    end else begin
      if (_T_281) begin
        _T_342 <= _T_339;
      end
    end
    if (reset) begin
      _T_345 <= 14'h0;
    end else begin
      if (_T_284) begin
        _T_345 <= _T_342;
      end
    end
    if (reset) begin
      _T_348 <= 14'h0;
    end else begin
      if (_T_287) begin
        _T_348 <= _T_345;
      end
    end
    if (reset) begin
      _T_351 <= 14'h0;
    end else begin
      if (_T_290) begin
        _T_351 <= _T_348;
      end
    end
  end
endmodule
module NV_soDLA_cdma( // @[:@24088.2]
  input          clock, // @[:@24089.4]
  input          reset, // @[:@24090.4]
  input          io_nvdla_clock_nvdla_core_clk, // @[:@24091.4]
  input          io_nvdla_clock_dla_clk_ovr_on_sync, // @[:@24091.4]
  input          io_nvdla_clock_global_clk_ovr_on_sync, // @[:@24091.4]
  input          io_nvdla_clock_tmc2slcg_disable_clock_gating, // @[:@24091.4]
  input          io_nvdla_core_rstn, // @[:@24091.4]
  output         io_csb2cdma_req_ready, // @[:@24091.4]
  input          io_csb2cdma_req_valid, // @[:@24091.4]
  input  [62:0]  io_csb2cdma_req_bits, // @[:@24091.4]
  output         io_csb2cdma_resp_valid, // @[:@24091.4]
  output [33:0]  io_csb2cdma_resp_bits, // @[:@24091.4]
  output [1:0]   io_cdma2buf_dat_wr_sel, // @[:@24091.4]
  output         io_cdma2buf_dat_wr_addr_valid, // @[:@24091.4]
  output [16:0]  io_cdma2buf_dat_wr_addr_bits, // @[:@24091.4]
  output [255:0] io_cdma2buf_dat_wr_data, // @[:@24091.4]
  output [1:0]   io_cdma2buf_wt_wr_sel, // @[:@24091.4]
  output         io_cdma2buf_wt_wr_addr_valid, // @[:@24091.4]
  output [16:0]  io_cdma2buf_wt_wr_addr_bits, // @[:@24091.4]
  output [255:0] io_cdma2buf_wt_wr_data, // @[:@24091.4]
  output [1:0]   io_cdma_dat2glb_done_intr_pd, // @[:@24091.4]
  output [1:0]   io_cdma_wt2glb_done_intr_pd, // @[:@24091.4]
  input          io_cdma_dat2cvif_rd_req_pd_ready, // @[:@24091.4]
  output         io_cdma_dat2cvif_rd_req_pd_valid, // @[:@24091.4]
  output [78:0]  io_cdma_dat2cvif_rd_req_pd_bits, // @[:@24091.4]
  output         io_cvif2cdma_dat_rd_rsp_pd_ready, // @[:@24091.4]
  input          io_cvif2cdma_dat_rd_rsp_pd_valid, // @[:@24091.4]
  input  [256:0] io_cvif2cdma_dat_rd_rsp_pd_bits, // @[:@24091.4]
  input          io_cdma_wt2cvif_rd_req_pd_ready, // @[:@24091.4]
  output         io_cdma_wt2cvif_rd_req_pd_valid, // @[:@24091.4]
  output [78:0]  io_cdma_wt2cvif_rd_req_pd_bits, // @[:@24091.4]
  output         io_cvif2cdma_wt_rd_rsp_pd_ready, // @[:@24091.4]
  input          io_cvif2cdma_wt_rd_rsp_pd_valid, // @[:@24091.4]
  input  [256:0] io_cvif2cdma_wt_rd_rsp_pd_bits, // @[:@24091.4]
  input          io_cdma_dat2mcif_rd_req_pd_ready, // @[:@24091.4]
  output         io_cdma_dat2mcif_rd_req_pd_valid, // @[:@24091.4]
  output [78:0]  io_cdma_dat2mcif_rd_req_pd_bits, // @[:@24091.4]
  output         io_mcif2cdma_dat_rd_rsp_pd_ready, // @[:@24091.4]
  input          io_mcif2cdma_dat_rd_rsp_pd_valid, // @[:@24091.4]
  input  [256:0] io_mcif2cdma_dat_rd_rsp_pd_bits, // @[:@24091.4]
  input          io_cdma_wt2mcif_rd_req_pd_ready, // @[:@24091.4]
  output         io_cdma_wt2mcif_rd_req_pd_valid, // @[:@24091.4]
  output [78:0]  io_cdma_wt2mcif_rd_req_pd_bits, // @[:@24091.4]
  output         io_mcif2cdma_wt_rd_rsp_pd_ready, // @[:@24091.4]
  input          io_mcif2cdma_wt_rd_rsp_pd_valid, // @[:@24091.4]
  input  [256:0] io_mcif2cdma_wt_rd_rsp_pd_bits, // @[:@24091.4]
  input          io_sc2cdma_dat_pending_req, // @[:@24091.4]
  input          io_sc2cdma_wt_pending_req, // @[:@24091.4]
  output         io_cdma2sc_dat_pending_ack, // @[:@24091.4]
  output         io_cdma2sc_wt_pending_ack, // @[:@24091.4]
  output         io_cdma2sc_dat_updt_valid, // @[:@24091.4]
  output [14:0]  io_cdma2sc_dat_updt_bits_entries, // @[:@24091.4]
  output [13:0]  io_cdma2sc_dat_updt_bits_slices, // @[:@24091.4]
  input          io_sc2cdma_dat_updt_valid, // @[:@24091.4]
  input  [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@24091.4]
  input  [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@24091.4]
  output         io_cdma2sc_wt_updt_valid, // @[:@24091.4]
  output [14:0]  io_cdma2sc_wt_updt_bits_entries, // @[:@24091.4]
  output [13:0]  io_cdma2sc_wt_updt_bits_kernels, // @[:@24091.4]
  input          io_sc2cdma_wt_updt_valid, // @[:@24091.4]
  input  [14:0]  io_sc2cdma_wt_updt_bits_entries, // @[:@24091.4]
  input  [13:0]  io_sc2cdma_wt_updt_bits_kernels, // @[:@24091.4]
  input  [31:0]  io_pwrbus_ram_pd // @[:@24091.4]
);
  wire  NV_NVDLA_CDMA_regfile_reset; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_csb2cdma_req_valid; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [62:0] NV_NVDLA_CDMA_regfile_io_csb2cdma_req_bits; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_valid; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [33:0] NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_bits; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_dp2reg_done; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_latency; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_stall; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_latency; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_stall; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_dp2reg_dat_flush_done; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_dp2reg_wt_flush_done; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_dp2reg_wt_rd_stall; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_dp2reg_consumer; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [4:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [4:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bank; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [4:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_batches; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_batch_stride; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_en; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [5:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_truncate; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_offset; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_scale; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_0; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_1; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_0; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_1; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_packed; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_packed; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_ram_type; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [5:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_format; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_sign_override; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [12:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_height; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [12:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_width; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [12:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_channel; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [13:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_entries; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [11:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_grains; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_stride; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_uv_line_stride; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_format; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_gu; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ry; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ax; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_bv; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_reuse; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [1:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_proc_precision; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_weight_rls; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_reuse; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_dma_en; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [4:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_x_offset; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_stride; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_high; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_low; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [31:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bytes; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_ram_type; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [17:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_byte_per_kernel; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [12:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_kernel; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [4:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_left; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [5:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_right; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire [15:0] NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_value; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
  wire  NV_NVDLA_CDMA_wt_reset; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_nvdla_core_ng_clk; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [78:0] NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [256:0] NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [78:0] NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [256:0] NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [1:0] NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_sel; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [16:0] NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_bits; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [255:0] NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_data; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [1:0] NV_NVDLA_CDMA_wt_io_wt2status_state; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [14:0] NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_entries; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [13:0] NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_kernels; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_cdma2sc_wt_pending_ack; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_valid; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [14:0] NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_bits_entries; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_sc2cdma_wt_pending_req; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_reg2dp_weight_reuse; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_reg2dp_skip_weight_rls; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [17:0] NV_NVDLA_CDMA_wt_io_reg2dp_byte_per_kernel; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [12:0] NV_NVDLA_CDMA_wt_io_reg2dp_weight_kernel; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_reg2dp_weight_ram_type; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [26:0] NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_low; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [31:0] NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_high; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [31:0] NV_NVDLA_CDMA_wt_io_reg2dp_weight_bytes; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [4:0] NV_NVDLA_CDMA_wt_io_reg2dp_data_bank; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [4:0] NV_NVDLA_CDMA_wt_io_reg2dp_weight_bank; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_reg2dp_dma_en; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_CDMA_wt_io_dp2reg_wt_flush_done; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire [31:0] NV_NVDLA_CDMA_wt_io_dp2reg_wt_rd_stall; // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
  wire  NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 88:27:@24099.4]
  wire  NV_NVDLA_slcg_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 88:27:@24099.4]
  wire  NV_NVDLA_CDMA_dc_reset; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_nvdla_core_ng_clk; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [78:0] NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [256:0] NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [78:0] NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [256:0] NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [16:0] NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [255:0] NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [11:0] NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_conv_mode; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_data_reuse; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_skip_data_rls; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_datain_format; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [12:0] NV_NVDLA_CDMA_dc_io_reg2dp_datain_width; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [12:0] NV_NVDLA_CDMA_dc_io_reg2dp_datain_height; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [12:0] NV_NVDLA_CDMA_dc_io_reg2dp_datain_channel; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_datain_ram_type; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [31:0] NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_high_0; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [26:0] NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_low_0; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [26:0] NV_NVDLA_CDMA_dc_io_reg2dp_line_stride; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [26:0] NV_NVDLA_CDMA_dc_io_reg2dp_surf_stride; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [26:0] NV_NVDLA_CDMA_dc_io_reg2dp_batch_stride; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_line_packed; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_surf_packed; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [4:0] NV_NVDLA_CDMA_dc_io_reg2dp_batches; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [16:0] NV_NVDLA_CDMA_dc_io_reg2dp_entries; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [11:0] NV_NVDLA_CDMA_dc_io_reg2dp_grains; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [4:0] NV_NVDLA_CDMA_dc_io_reg2dp_data_bank; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_reg2dp_dma_en; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [31:0] NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_stall; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [31:0] NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_latency; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [1:0] NV_NVDLA_CDMA_dc_io_dc2status_state; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [14:0] NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [13:0] NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [14:0] NV_NVDLA_CDMA_dc_io_status2dma_free_entries; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [14:0] NV_NVDLA_CDMA_dc_io_status2dma_wr_idx; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [7:0] NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [255:0] NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_data; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [7:0] NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire [255:0] NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_data; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_CDMA_dc_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
  wire  NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 90:27:@24105.4]
  wire  NV_NVDLA_slcg_1_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 90:27:@24105.4]
  wire  NV_NVDLA_CDMA_img_reset; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_nvdla_core_ng_clk; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [78:0] NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [256:0] NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [78:0] NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [256:0] NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [16:0] NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [255:0] NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [511:0] NV_NVDLA_CDMA_img_io_img2cvt_mn_wr_data; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_pad_mask; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [11:0] NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [1:0] NV_NVDLA_CDMA_img_io_img2status_state; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [14:0] NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [13:0] NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [14:0] NV_NVDLA_CDMA_img_io_status2dma_free_entries; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [14:0] NV_NVDLA_CDMA_img_io_status2dma_wr_idx; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [7:0] NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [255:0] NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_data; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [7:0] NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [255:0] NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_data; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_conv_mode; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_data_reuse; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_skip_data_rls; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_datain_format; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [5:0] NV_NVDLA_CDMA_img_io_reg2dp_pixel_format; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_pixel_sign_override; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [12:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_width; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [12:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_height; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [12:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_channel; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [4:0] NV_NVDLA_CDMA_img_io_reg2dp_pixel_x_offset; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_datain_ram_type; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_0; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_0; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_1; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_line_stride; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_uv_line_stride; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_1; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_mean_format; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [15:0] NV_NVDLA_CDMA_img_io_reg2dp_mean_ry; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [15:0] NV_NVDLA_CDMA_img_io_reg2dp_mean_gu; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [15:0] NV_NVDLA_CDMA_img_io_reg2dp_mean_bv; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [15:0] NV_NVDLA_CDMA_img_io_reg2dp_mean_ax; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [13:0] NV_NVDLA_CDMA_img_io_reg2dp_entries; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [4:0] NV_NVDLA_CDMA_img_io_reg2dp_pad_left; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [5:0] NV_NVDLA_CDMA_img_io_reg2dp_pad_right; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [4:0] NV_NVDLA_CDMA_img_io_reg2dp_data_bank; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_CDMA_img_io_reg2dp_dma_en; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_dp2reg_img_rd_stall; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire [31:0] NV_NVDLA_CDMA_img_io_dp2reg_img_rd_latency; // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
  wire  NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 92:28:@24111.4]
  wire  NV_NVDLA_slcg_2_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 92:28:@24111.4]
  wire  NV_NVDLA_CDMA_dma_mux_reset; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [78:0] NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire [256:0] NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
  wire  NV_NVDLA_slcg_3_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 94:28:@24117.4]
  wire  NV_NVDLA_slcg_3_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 94:28:@24117.4]
  wire  NV_NVDLA_CDMA_cvt_reset; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_nvdla_core_ng_clk; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_nvdla_hls_clk; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [16:0] NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [255:0] NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [11:0] NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [16:0] NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [255:0] NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [511:0] NV_NVDLA_CDMA_cvt_io_img2cvt_mn_wr_data; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [31:0] NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_pad_mask; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [11:0] NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [1:0] NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_sel; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [16:0] NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [255:0] NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_data; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [1:0] NV_NVDLA_CDMA_cvt_io_reg2dp_proc_precision; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_en; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [5:0] NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_truncate; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [15:0] NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_offset; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [15:0] NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_scale; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire [15:0] NV_NVDLA_CDMA_cvt_io_reg2dp_pad_value; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_dp2reg_done; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_CDMA_cvt_io_dp2reg_dat_flush_done; // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
  wire  NV_NVDLA_slcg_4_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 96:28:@24123.4]
  wire  NV_NVDLA_slcg_4_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 96:28:@24123.4]
  wire  NV_NVDLA_slcg_5_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 97:28:@24126.4]
  wire  NV_NVDLA_slcg_5_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 97:28:@24126.4]
  wire  NV_NVDLA_CDMA_shared_buffer_reset; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_CDMA_shared_buffer_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [7:0] NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_bits; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [255:0] NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_data; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_valid; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [7:0] NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_bits; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [255:0] NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_data; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [7:0] NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_bits; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [255:0] NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_data; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_valid; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [7:0] NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_bits; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire [255:0] NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_data; // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
  wire  NV_NVDLA_slcg_6_io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 99:31:@24132.4]
  wire  NV_NVDLA_slcg_6_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 99:31:@24132.4]
  wire  NV_NVDLA_CDMA_status_reset; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_dc2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [13:0] NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_img2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [13:0] NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_valid; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_valid; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [13:0] NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_status2dma_free_entries; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [14:0] NV_NVDLA_CDMA_status_io_status2dma_wr_idx; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_dc2status_state; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_img2status_state; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_wt2status_state; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_dp2reg_consumer; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_dp2reg_done; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [4:0] NV_NVDLA_CDMA_status_io_reg2dp_data_bank; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_cdma_wt2glb_done_intr_pd; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_cdma_dat2glb_done_intr_pd; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_sc2cdma_dat_pending_req; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire [1:0] NV_NVDLA_CDMA_status_io_cdma2sc_dat_pending_ack; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  wire  NV_NVDLA_CDMA_status_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
  NV_NVDLA_CDMA_regfile NV_NVDLA_CDMA_regfile ( // @[NV_NVDLA_cdma.scala 86:27:@24093.4]
    .reset(NV_NVDLA_CDMA_regfile_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_regfile_io_nvdla_core_clk),
    .io_csb2cdma_req_valid(NV_NVDLA_CDMA_regfile_io_csb2cdma_req_valid),
    .io_csb2cdma_req_bits(NV_NVDLA_CDMA_regfile_io_csb2cdma_req_bits),
    .io_csb2cdma_resp_valid(NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_valid),
    .io_csb2cdma_resp_bits(NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_bits),
    .io_dp2reg_done(NV_NVDLA_CDMA_regfile_io_dp2reg_done),
    .io_dp2reg_dc_rd_latency(NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_latency),
    .io_dp2reg_dc_rd_stall(NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_stall),
    .io_dp2reg_img_rd_latency(NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_latency),
    .io_dp2reg_img_rd_stall(NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_stall),
    .io_dp2reg_dat_flush_done(NV_NVDLA_CDMA_regfile_io_dp2reg_dat_flush_done),
    .io_dp2reg_wt_flush_done(NV_NVDLA_CDMA_regfile_io_dp2reg_wt_flush_done),
    .io_dp2reg_wt_rd_stall(NV_NVDLA_CDMA_regfile_io_dp2reg_wt_rd_stall),
    .io_dp2reg_consumer(NV_NVDLA_CDMA_regfile_io_dp2reg_consumer),
    .io_reg2dp_field_data_bank(NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank),
    .io_reg2dp_field_weight_bank(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bank),
    .io_reg2dp_field_batches(NV_NVDLA_CDMA_regfile_io_reg2dp_field_batches),
    .io_reg2dp_field_batch_stride(NV_NVDLA_CDMA_regfile_io_reg2dp_field_batch_stride),
    .io_reg2dp_field_cvt_en(NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_en),
    .io_reg2dp_field_cvt_truncate(NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_truncate),
    .io_reg2dp_field_cvt_offset(NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_offset),
    .io_reg2dp_field_cvt_scale(NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_scale),
    .io_reg2dp_field_datain_addr_high_0(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_0),
    .io_reg2dp_field_datain_addr_high_1(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_1),
    .io_reg2dp_field_datain_addr_low_0(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_0),
    .io_reg2dp_field_datain_addr_low_1(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_1),
    .io_reg2dp_field_line_packed(NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_packed),
    .io_reg2dp_field_surf_packed(NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_packed),
    .io_reg2dp_field_datain_ram_type(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_ram_type),
    .io_reg2dp_field_datain_format(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_format),
    .io_reg2dp_field_pixel_format(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_format),
    .io_reg2dp_field_pixel_sign_override(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_sign_override),
    .io_reg2dp_field_datain_height(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_height),
    .io_reg2dp_field_datain_width(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_width),
    .io_reg2dp_field_datain_channel(NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_channel),
    .io_reg2dp_field_entries(NV_NVDLA_CDMA_regfile_io_reg2dp_field_entries),
    .io_reg2dp_field_grains(NV_NVDLA_CDMA_regfile_io_reg2dp_field_grains),
    .io_reg2dp_field_line_stride(NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_stride),
    .io_reg2dp_field_uv_line_stride(NV_NVDLA_CDMA_regfile_io_reg2dp_field_uv_line_stride),
    .io_reg2dp_field_mean_format(NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_format),
    .io_reg2dp_field_mean_gu(NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_gu),
    .io_reg2dp_field_mean_ry(NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ry),
    .io_reg2dp_field_mean_ax(NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ax),
    .io_reg2dp_field_mean_bv(NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_bv),
    .io_reg2dp_field_conv_mode(NV_NVDLA_CDMA_regfile_io_reg2dp_field_conv_mode),
    .io_reg2dp_field_data_reuse(NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_reuse),
    .io_reg2dp_field_proc_precision(NV_NVDLA_CDMA_regfile_io_reg2dp_field_proc_precision),
    .io_reg2dp_field_skip_data_rls(NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_data_rls),
    .io_reg2dp_field_skip_weight_rls(NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_weight_rls),
    .io_reg2dp_field_weight_reuse(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_reuse),
    .io_reg2dp_field_dma_en(NV_NVDLA_CDMA_regfile_io_reg2dp_field_dma_en),
    .io_reg2dp_field_pixel_x_offset(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_x_offset),
    .io_reg2dp_field_surf_stride(NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_stride),
    .io_reg2dp_field_weight_addr_high(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_high),
    .io_reg2dp_field_weight_addr_low(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_low),
    .io_reg2dp_field_weight_bytes(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bytes),
    .io_reg2dp_field_weight_ram_type(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_ram_type),
    .io_reg2dp_field_byte_per_kernel(NV_NVDLA_CDMA_regfile_io_reg2dp_field_byte_per_kernel),
    .io_reg2dp_field_weight_kernel(NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_kernel),
    .io_reg2dp_field_pad_left(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_left),
    .io_reg2dp_field_pad_right(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_right),
    .io_reg2dp_field_pad_value(NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_value),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_regfile_io_reg2dp_op_en)
  );
  NV_NVDLA_CDMA_wt NV_NVDLA_CDMA_wt ( // @[NV_NVDLA_cdma.scala 87:22:@24096.4]
    .reset(NV_NVDLA_CDMA_wt_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_wt_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CDMA_wt_io_nvdla_core_ng_clk),
    .io_cdma_wt2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_ready),
    .io_cdma_wt2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_valid),
    .io_cdma_wt2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_bits),
    .io_mcif2cdma_wt_rd_rsp_pd_ready(NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_ready),
    .io_mcif2cdma_wt_rd_rsp_pd_valid(NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_valid),
    .io_mcif2cdma_wt_rd_rsp_pd_bits(NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_bits),
    .io_cdma_wt2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_ready),
    .io_cdma_wt2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_valid),
    .io_cdma_wt2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_bits),
    .io_cvif2cdma_wt_rd_rsp_pd_ready(NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_ready),
    .io_cvif2cdma_wt_rd_rsp_pd_valid(NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_valid),
    .io_cvif2cdma_wt_rd_rsp_pd_bits(NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_bits),
    .io_cdma2buf_wt_wr_sel(NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_sel),
    .io_cdma2buf_wt_wr_addr_valid(NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_valid),
    .io_cdma2buf_wt_wr_addr_bits(NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_bits),
    .io_cdma2buf_wt_wr_data(NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_data),
    .io_status2dma_fsm_switch(NV_NVDLA_CDMA_wt_io_status2dma_fsm_switch),
    .io_wt2status_state(NV_NVDLA_CDMA_wt_io_wt2status_state),
    .io_cdma2sc_wt_updt_valid(NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_valid),
    .io_cdma2sc_wt_updt_bits_entries(NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_entries),
    .io_cdma2sc_wt_updt_bits_kernels(NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_kernels),
    .io_cdma2sc_wt_pending_ack(NV_NVDLA_CDMA_wt_io_cdma2sc_wt_pending_ack),
    .io_sc2cdma_wt_updt_valid(NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_valid),
    .io_sc2cdma_wt_updt_bits_entries(NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_bits_entries),
    .io_sc2cdma_wt_pending_req(NV_NVDLA_CDMA_wt_io_sc2cdma_wt_pending_req),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_wt_io_reg2dp_op_en),
    .io_reg2dp_weight_reuse(NV_NVDLA_CDMA_wt_io_reg2dp_weight_reuse),
    .io_reg2dp_skip_weight_rls(NV_NVDLA_CDMA_wt_io_reg2dp_skip_weight_rls),
    .io_reg2dp_byte_per_kernel(NV_NVDLA_CDMA_wt_io_reg2dp_byte_per_kernel),
    .io_reg2dp_weight_kernel(NV_NVDLA_CDMA_wt_io_reg2dp_weight_kernel),
    .io_reg2dp_weight_ram_type(NV_NVDLA_CDMA_wt_io_reg2dp_weight_ram_type),
    .io_reg2dp_weight_addr_low(NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_low),
    .io_reg2dp_weight_addr_high(NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_high),
    .io_reg2dp_weight_bytes(NV_NVDLA_CDMA_wt_io_reg2dp_weight_bytes),
    .io_reg2dp_data_bank(NV_NVDLA_CDMA_wt_io_reg2dp_data_bank),
    .io_reg2dp_weight_bank(NV_NVDLA_CDMA_wt_io_reg2dp_weight_bank),
    .io_reg2dp_dma_en(NV_NVDLA_CDMA_wt_io_reg2dp_dma_en),
    .io_dp2reg_wt_flush_done(NV_NVDLA_CDMA_wt_io_dp2reg_wt_flush_done),
    .io_dp2reg_wt_rd_stall(NV_NVDLA_CDMA_wt_io_dp2reg_wt_rd_stall)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg ( // @[NV_NVDLA_cdma.scala 88:27:@24099.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_dc NV_NVDLA_CDMA_dc ( // @[NV_NVDLA_cdma.scala 89:22:@24102.4]
    .reset(NV_NVDLA_CDMA_dc_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_dc_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CDMA_dc_io_nvdla_core_ng_clk),
    .io_dc_dat2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_ready),
    .io_dc_dat2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_valid),
    .io_dc_dat2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_bits),
    .io_mcif2dc_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_ready),
    .io_mcif2dc_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_valid),
    .io_mcif2dc_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_bits),
    .io_dc_dat2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_ready),
    .io_dc_dat2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_valid),
    .io_dc_dat2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_bits),
    .io_cvif2dc_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_ready),
    .io_cvif2dc_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_valid),
    .io_cvif2dc_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_bits),
    .io_dc2cvt_dat_wr_sel(NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_sel),
    .io_dc2cvt_dat_wr_addr_valid(NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_valid),
    .io_dc2cvt_dat_wr_addr_bits(NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_bits),
    .io_dc2cvt_dat_wr_data(NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_data),
    .io_dc2cvt_dat_wr_info_pd(NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_info_pd),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_dc_io_reg2dp_op_en),
    .io_reg2dp_conv_mode(NV_NVDLA_CDMA_dc_io_reg2dp_conv_mode),
    .io_reg2dp_data_reuse(NV_NVDLA_CDMA_dc_io_reg2dp_data_reuse),
    .io_reg2dp_skip_data_rls(NV_NVDLA_CDMA_dc_io_reg2dp_skip_data_rls),
    .io_reg2dp_datain_format(NV_NVDLA_CDMA_dc_io_reg2dp_datain_format),
    .io_reg2dp_datain_width(NV_NVDLA_CDMA_dc_io_reg2dp_datain_width),
    .io_reg2dp_datain_height(NV_NVDLA_CDMA_dc_io_reg2dp_datain_height),
    .io_reg2dp_datain_channel(NV_NVDLA_CDMA_dc_io_reg2dp_datain_channel),
    .io_reg2dp_datain_ram_type(NV_NVDLA_CDMA_dc_io_reg2dp_datain_ram_type),
    .io_reg2dp_datain_addr_high_0(NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_high_0),
    .io_reg2dp_datain_addr_low_0(NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_low_0),
    .io_reg2dp_line_stride(NV_NVDLA_CDMA_dc_io_reg2dp_line_stride),
    .io_reg2dp_surf_stride(NV_NVDLA_CDMA_dc_io_reg2dp_surf_stride),
    .io_reg2dp_batch_stride(NV_NVDLA_CDMA_dc_io_reg2dp_batch_stride),
    .io_reg2dp_line_packed(NV_NVDLA_CDMA_dc_io_reg2dp_line_packed),
    .io_reg2dp_surf_packed(NV_NVDLA_CDMA_dc_io_reg2dp_surf_packed),
    .io_reg2dp_batches(NV_NVDLA_CDMA_dc_io_reg2dp_batches),
    .io_reg2dp_entries(NV_NVDLA_CDMA_dc_io_reg2dp_entries),
    .io_reg2dp_grains(NV_NVDLA_CDMA_dc_io_reg2dp_grains),
    .io_reg2dp_data_bank(NV_NVDLA_CDMA_dc_io_reg2dp_data_bank),
    .io_reg2dp_dma_en(NV_NVDLA_CDMA_dc_io_reg2dp_dma_en),
    .io_dp2reg_dc_rd_stall(NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_stall),
    .io_dp2reg_dc_rd_latency(NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_latency),
    .io_dc2status_state(NV_NVDLA_CDMA_dc_io_dc2status_state),
    .io_dc2status_dat_updt_valid(NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_valid),
    .io_dc2status_dat_updt_bits_entries(NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_entries),
    .io_dc2status_dat_updt_bits_slices(NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_slices),
    .io_status2dma_fsm_switch(NV_NVDLA_CDMA_dc_io_status2dma_fsm_switch),
    .io_status2dma_free_entries(NV_NVDLA_CDMA_dc_io_status2dma_free_entries),
    .io_status2dma_wr_idx(NV_NVDLA_CDMA_dc_io_status2dma_wr_idx),
    .io_dc2sbuf_p0_wr_addr_valid(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_valid),
    .io_dc2sbuf_p0_wr_addr_bits(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_bits),
    .io_dc2sbuf_p0_wr_data(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_data),
    .io_dc2sbuf_p0_rd_addr_valid(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_valid),
    .io_dc2sbuf_p0_rd_addr_bits(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_bits),
    .io_dc2sbuf_p0_rd_data(NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_data),
    .io_sc2cdma_dat_pending_req(NV_NVDLA_CDMA_dc_io_sc2cdma_dat_pending_req)
  );
  NV_NVDLA_slcg_1 NV_NVDLA_slcg_1 ( // @[NV_NVDLA_cdma.scala 90:27:@24105.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_1_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_img NV_NVDLA_CDMA_img ( // @[NV_NVDLA_cdma.scala 91:23:@24108.4]
    .reset(NV_NVDLA_CDMA_img_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_img_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CDMA_img_io_nvdla_core_ng_clk),
    .io_img_dat2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_ready),
    .io_img_dat2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_valid),
    .io_img_dat2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_bits),
    .io_mcif2img_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_ready),
    .io_mcif2img_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_valid),
    .io_mcif2img_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_bits),
    .io_img_dat2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_ready),
    .io_img_dat2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_valid),
    .io_img_dat2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_bits),
    .io_cvif2img_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_ready),
    .io_cvif2img_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_valid),
    .io_cvif2img_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_bits),
    .io_img2cvt_dat_wr_sel(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_sel),
    .io_img2cvt_dat_wr_addr_valid(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_valid),
    .io_img2cvt_dat_wr_addr_bits(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_bits),
    .io_img2cvt_dat_wr_data(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_data),
    .io_img2cvt_mn_wr_data(NV_NVDLA_CDMA_img_io_img2cvt_mn_wr_data),
    .io_img2cvt_dat_wr_pad_mask(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_pad_mask),
    .io_img2cvt_dat_wr_info_pd(NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_info_pd),
    .io_img2status_state(NV_NVDLA_CDMA_img_io_img2status_state),
    .io_img2status_dat_updt_valid(NV_NVDLA_CDMA_img_io_img2status_dat_updt_valid),
    .io_img2status_dat_updt_bits_entries(NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_entries),
    .io_img2status_dat_updt_bits_slices(NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_slices),
    .io_status2dma_free_entries(NV_NVDLA_CDMA_img_io_status2dma_free_entries),
    .io_status2dma_wr_idx(NV_NVDLA_CDMA_img_io_status2dma_wr_idx),
    .io_status2dma_fsm_switch(NV_NVDLA_CDMA_img_io_status2dma_fsm_switch),
    .io_img2sbuf_p0_wr_addr_valid(NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_valid),
    .io_img2sbuf_p0_wr_addr_bits(NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_bits),
    .io_img2sbuf_p0_wr_data(NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_data),
    .io_img2sbuf_p0_rd_addr_valid(NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_valid),
    .io_img2sbuf_p0_rd_addr_bits(NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_bits),
    .io_img2sbuf_p0_rd_data(NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_data),
    .io_sc2cdma_dat_pending_req(NV_NVDLA_CDMA_img_io_sc2cdma_dat_pending_req),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_img_io_reg2dp_op_en),
    .io_reg2dp_conv_mode(NV_NVDLA_CDMA_img_io_reg2dp_conv_mode),
    .io_reg2dp_data_reuse(NV_NVDLA_CDMA_img_io_reg2dp_data_reuse),
    .io_reg2dp_skip_data_rls(NV_NVDLA_CDMA_img_io_reg2dp_skip_data_rls),
    .io_reg2dp_datain_format(NV_NVDLA_CDMA_img_io_reg2dp_datain_format),
    .io_reg2dp_pixel_format(NV_NVDLA_CDMA_img_io_reg2dp_pixel_format),
    .io_reg2dp_pixel_sign_override(NV_NVDLA_CDMA_img_io_reg2dp_pixel_sign_override),
    .io_reg2dp_datain_width(NV_NVDLA_CDMA_img_io_reg2dp_datain_width),
    .io_reg2dp_datain_height(NV_NVDLA_CDMA_img_io_reg2dp_datain_height),
    .io_reg2dp_datain_channel(NV_NVDLA_CDMA_img_io_reg2dp_datain_channel),
    .io_reg2dp_pixel_x_offset(NV_NVDLA_CDMA_img_io_reg2dp_pixel_x_offset),
    .io_reg2dp_datain_ram_type(NV_NVDLA_CDMA_img_io_reg2dp_datain_ram_type),
    .io_reg2dp_datain_addr_high_0(NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_0),
    .io_reg2dp_datain_addr_low_0(NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_0),
    .io_reg2dp_datain_addr_low_1(NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_1),
    .io_reg2dp_line_stride(NV_NVDLA_CDMA_img_io_reg2dp_line_stride),
    .io_reg2dp_uv_line_stride(NV_NVDLA_CDMA_img_io_reg2dp_uv_line_stride),
    .io_reg2dp_datain_addr_high_1(NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_1),
    .io_reg2dp_mean_format(NV_NVDLA_CDMA_img_io_reg2dp_mean_format),
    .io_reg2dp_mean_ry(NV_NVDLA_CDMA_img_io_reg2dp_mean_ry),
    .io_reg2dp_mean_gu(NV_NVDLA_CDMA_img_io_reg2dp_mean_gu),
    .io_reg2dp_mean_bv(NV_NVDLA_CDMA_img_io_reg2dp_mean_bv),
    .io_reg2dp_mean_ax(NV_NVDLA_CDMA_img_io_reg2dp_mean_ax),
    .io_reg2dp_entries(NV_NVDLA_CDMA_img_io_reg2dp_entries),
    .io_reg2dp_pad_left(NV_NVDLA_CDMA_img_io_reg2dp_pad_left),
    .io_reg2dp_pad_right(NV_NVDLA_CDMA_img_io_reg2dp_pad_right),
    .io_reg2dp_data_bank(NV_NVDLA_CDMA_img_io_reg2dp_data_bank),
    .io_reg2dp_dma_en(NV_NVDLA_CDMA_img_io_reg2dp_dma_en),
    .io_dp2reg_img_rd_stall(NV_NVDLA_CDMA_img_io_dp2reg_img_rd_stall),
    .io_dp2reg_img_rd_latency(NV_NVDLA_CDMA_img_io_dp2reg_img_rd_latency)
  );
  NV_NVDLA_slcg_1 NV_NVDLA_slcg_2 ( // @[NV_NVDLA_cdma.scala 92:28:@24111.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_2_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_dma_mux NV_NVDLA_CDMA_dma_mux ( // @[NV_NVDLA_cdma.scala 93:27:@24114.4]
    .reset(NV_NVDLA_CDMA_dma_mux_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_dma_mux_io_nvdla_core_clk),
    .io_dc_dat2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_ready),
    .io_dc_dat2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_valid),
    .io_dc_dat2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_bits),
    .io_mcif2dc_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_ready),
    .io_mcif2dc_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_valid),
    .io_mcif2dc_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_bits),
    .io_img_dat2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_ready),
    .io_img_dat2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_valid),
    .io_img_dat2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_bits),
    .io_mcif2img_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_ready),
    .io_mcif2img_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_valid),
    .io_mcif2img_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_bits),
    .io_cdma_dat2mcif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_ready),
    .io_cdma_dat2mcif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_valid),
    .io_cdma_dat2mcif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_bits),
    .io_mcif2cdma_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_ready),
    .io_mcif2cdma_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_valid),
    .io_mcif2cdma_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_bits),
    .io_dc_dat2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_ready),
    .io_dc_dat2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_valid),
    .io_dc_dat2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_bits),
    .io_cvif2dc_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_ready),
    .io_cvif2dc_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_valid),
    .io_cvif2dc_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_bits),
    .io_img_dat2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_ready),
    .io_img_dat2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_valid),
    .io_img_dat2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_bits),
    .io_cvif2img_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_ready),
    .io_cvif2img_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_valid),
    .io_cvif2img_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_bits),
    .io_cdma_dat2cvif_rd_req_pd_ready(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_ready),
    .io_cdma_dat2cvif_rd_req_pd_valid(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_valid),
    .io_cdma_dat2cvif_rd_req_pd_bits(NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_bits),
    .io_cvif2cdma_dat_rd_rsp_pd_ready(NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_ready),
    .io_cvif2cdma_dat_rd_rsp_pd_valid(NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_valid),
    .io_cvif2cdma_dat_rd_rsp_pd_bits(NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_bits)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg_3 ( // @[NV_NVDLA_cdma.scala 94:28:@24117.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_3_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_3_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_cvt NV_NVDLA_CDMA_cvt ( // @[NV_NVDLA_cdma.scala 95:23:@24120.4]
    .reset(NV_NVDLA_CDMA_cvt_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_cvt_io_nvdla_core_clk),
    .io_nvdla_core_ng_clk(NV_NVDLA_CDMA_cvt_io_nvdla_core_ng_clk),
    .io_nvdla_hls_clk(NV_NVDLA_CDMA_cvt_io_nvdla_hls_clk),
    .io_dc2cvt_dat_wr_sel(NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_sel),
    .io_dc2cvt_dat_wr_addr_valid(NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_valid),
    .io_dc2cvt_dat_wr_addr_bits(NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_bits),
    .io_dc2cvt_dat_wr_data(NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_data),
    .io_dc2cvt_dat_wr_info_pd(NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_info_pd),
    .io_img2cvt_dat_wr_sel(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_sel),
    .io_img2cvt_dat_wr_addr_valid(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_valid),
    .io_img2cvt_dat_wr_addr_bits(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_bits),
    .io_img2cvt_dat_wr_data(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_data),
    .io_img2cvt_mn_wr_data(NV_NVDLA_CDMA_cvt_io_img2cvt_mn_wr_data),
    .io_img2cvt_dat_wr_pad_mask(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_pad_mask),
    .io_img2cvt_dat_wr_info_pd(NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_info_pd),
    .io_cdma2buf_dat_wr_sel(NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_sel),
    .io_cdma2buf_dat_wr_addr_valid(NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_valid),
    .io_cdma2buf_dat_wr_addr_bits(NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_bits),
    .io_cdma2buf_dat_wr_data(NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_data),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_cvt_io_reg2dp_op_en),
    .io_reg2dp_proc_precision(NV_NVDLA_CDMA_cvt_io_reg2dp_proc_precision),
    .io_reg2dp_cvt_en(NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_en),
    .io_reg2dp_cvt_truncate(NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_truncate),
    .io_reg2dp_cvt_offset(NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_offset),
    .io_reg2dp_cvt_scale(NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_scale),
    .io_reg2dp_pad_value(NV_NVDLA_CDMA_cvt_io_reg2dp_pad_value),
    .io_dp2reg_done(NV_NVDLA_CDMA_cvt_io_dp2reg_done),
    .io_dp2reg_dat_flush_done(NV_NVDLA_CDMA_cvt_io_dp2reg_dat_flush_done)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg_4 ( // @[NV_NVDLA_cdma.scala 96:28:@24123.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_4_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_4_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_slcg_5 NV_NVDLA_slcg_5 ( // @[NV_NVDLA_cdma.scala 97:28:@24126.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_5_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_5_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_shared_buffer NV_NVDLA_CDMA_shared_buffer ( // @[NV_NVDLA_cdma.scala 98:33:@24129.4]
    .reset(NV_NVDLA_CDMA_shared_buffer_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_shared_buffer_io_nvdla_core_clk),
    .io_dc2sbuf_p_wr_0_addr_valid(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_valid),
    .io_dc2sbuf_p_wr_0_addr_bits(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_bits),
    .io_dc2sbuf_p_wr_0_data(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_data),
    .io_img2sbuf_p_wr_0_addr_valid(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_valid),
    .io_img2sbuf_p_wr_0_addr_bits(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_bits),
    .io_img2sbuf_p_wr_0_data(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_data),
    .io_dc2sbuf_p_rd_0_addr_valid(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_valid),
    .io_dc2sbuf_p_rd_0_addr_bits(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_bits),
    .io_dc2sbuf_p_rd_0_data(NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_data),
    .io_img2sbuf_p_rd_0_addr_valid(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_valid),
    .io_img2sbuf_p_rd_0_addr_bits(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_bits),
    .io_img2sbuf_p_rd_0_data(NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_data)
  );
  NV_NVDLA_slcg NV_NVDLA_slcg_6 ( // @[NV_NVDLA_cdma.scala 99:31:@24132.4]
    .io_nvdla_clock_nvdla_core_clk(NV_NVDLA_slcg_6_io_nvdla_clock_nvdla_core_clk),
    .io_nvdla_core_gated_clk(NV_NVDLA_slcg_6_io_nvdla_core_gated_clk)
  );
  NV_NVDLA_CDMA_status NV_NVDLA_CDMA_status ( // @[NV_NVDLA_cdma.scala 100:26:@24135.4]
    .reset(NV_NVDLA_CDMA_status_reset),
    .io_nvdla_core_clk(NV_NVDLA_CDMA_status_io_nvdla_core_clk),
    .io_dc2status_dat_updt_valid(NV_NVDLA_CDMA_status_io_dc2status_dat_updt_valid),
    .io_dc2status_dat_updt_bits_entries(NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_entries),
    .io_dc2status_dat_updt_bits_slices(NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_slices),
    .io_img2status_dat_updt_valid(NV_NVDLA_CDMA_status_io_img2status_dat_updt_valid),
    .io_img2status_dat_updt_bits_entries(NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_entries),
    .io_img2status_dat_updt_bits_slices(NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_slices),
    .io_sc2cdma_dat_updt_valid(NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_valid),
    .io_sc2cdma_dat_updt_bits_entries(NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_bits_entries),
    .io_cdma2sc_dat_updt_valid(NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_valid),
    .io_cdma2sc_dat_updt_bits_entries(NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_entries),
    .io_cdma2sc_dat_updt_bits_slices(NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_slices),
    .io_status2dma_free_entries(NV_NVDLA_CDMA_status_io_status2dma_free_entries),
    .io_status2dma_wr_idx(NV_NVDLA_CDMA_status_io_status2dma_wr_idx),
    .io_dc2status_state(NV_NVDLA_CDMA_status_io_dc2status_state),
    .io_img2status_state(NV_NVDLA_CDMA_status_io_img2status_state),
    .io_wt2status_state(NV_NVDLA_CDMA_status_io_wt2status_state),
    .io_dp2reg_consumer(NV_NVDLA_CDMA_status_io_dp2reg_consumer),
    .io_dp2reg_done(NV_NVDLA_CDMA_status_io_dp2reg_done),
    .io_reg2dp_op_en(NV_NVDLA_CDMA_status_io_reg2dp_op_en),
    .io_reg2dp_data_bank(NV_NVDLA_CDMA_status_io_reg2dp_data_bank),
    .io_cdma_wt2glb_done_intr_pd(NV_NVDLA_CDMA_status_io_cdma_wt2glb_done_intr_pd),
    .io_cdma_dat2glb_done_intr_pd(NV_NVDLA_CDMA_status_io_cdma_dat2glb_done_intr_pd),
    .io_sc2cdma_dat_pending_req(NV_NVDLA_CDMA_status_io_sc2cdma_dat_pending_req),
    .io_cdma2sc_dat_pending_ack(NV_NVDLA_CDMA_status_io_cdma2sc_dat_pending_ack),
    .io_status2dma_fsm_switch(NV_NVDLA_CDMA_status_io_status2dma_fsm_switch)
  );
  assign io_csb2cdma_req_ready = 1'h1; // @[NV_NVDLA_cdma.scala 106:27:@24143.4]
  assign io_csb2cdma_resp_valid = NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_valid; // @[NV_NVDLA_cdma.scala 106:27:@24140.4]
  assign io_csb2cdma_resp_bits = NV_NVDLA_CDMA_regfile_io_csb2cdma_resp_bits; // @[NV_NVDLA_cdma.scala 106:27:@24139.4]
  assign io_cdma2buf_dat_wr_sel = NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_sel; // @[NV_NVDLA_cdma.scala 373:36:@24388.4]
  assign io_cdma2buf_dat_wr_addr_valid = NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 375:24:@24391.4]
  assign io_cdma2buf_dat_wr_addr_bits = NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 375:24:@24390.4]
  assign io_cdma2buf_dat_wr_data = NV_NVDLA_CDMA_cvt_io_cdma2buf_dat_wr_data; // @[NV_NVDLA_cdma.scala 375:24:@24389.4]
  assign io_cdma2buf_wt_wr_sel = NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_sel; // @[NV_NVDLA_cdma.scala 151:35:@24174.4]
  assign io_cdma2buf_wt_wr_addr_valid = NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_valid; // @[NV_NVDLA_cdma.scala 153:23:@24177.4]
  assign io_cdma2buf_wt_wr_addr_bits = NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_addr_bits; // @[NV_NVDLA_cdma.scala 153:23:@24176.4]
  assign io_cdma2buf_wt_wr_data = NV_NVDLA_CDMA_wt_io_cdma2buf_wt_wr_data; // @[NV_NVDLA_cdma.scala 153:23:@24175.4]
  assign io_cdma_dat2glb_done_intr_pd = NV_NVDLA_CDMA_status_io_cdma_dat2glb_done_intr_pd; // @[NV_NVDLA_cdma.scala 439:34:@24444.4]
  assign io_cdma_wt2glb_done_intr_pd = NV_NVDLA_CDMA_status_io_cdma_wt2glb_done_intr_pd; // @[NV_NVDLA_cdma.scala 438:33:@24443.4]
  assign io_cdma_dat2cvif_rd_req_pd_valid = NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 354:40:@24374.4]
  assign io_cdma_dat2cvif_rd_req_pd_bits = NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 354:40:@24373.4]
  assign io_cvif2cdma_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 355:50:@24378.4]
  assign io_cdma_wt2cvif_rd_req_pd_valid = NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 146:40:@24169.4]
  assign io_cdma_wt2cvif_rd_req_pd_bits = NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 146:40:@24168.4]
  assign io_cvif2cdma_wt_rd_rsp_pd_ready = NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 147:44:@24173.4]
  assign io_cdma_dat2mcif_rd_req_pd_valid = NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 350:32:@24368.4]
  assign io_cdma_dat2mcif_rd_req_pd_bits = NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 350:32:@24367.4]
  assign io_mcif2cdma_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 351:42:@24372.4]
  assign io_cdma_wt2mcif_rd_req_pd_valid = NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 142:31:@24163.4]
  assign io_cdma_wt2mcif_rd_req_pd_bits = NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 142:31:@24162.4]
  assign io_mcif2cdma_wt_rd_rsp_pd_ready = NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 143:36:@24167.4]
  assign io_cdma2sc_dat_pending_ack = NV_NVDLA_CDMA_status_io_cdma2sc_dat_pending_ack[0]; // @[NV_NVDLA_cdma.scala 442:32:@24446.4]
  assign io_cdma2sc_wt_pending_ack = NV_NVDLA_CDMA_wt_io_cdma2sc_wt_pending_ack; // @[NV_NVDLA_cdma.scala 159:31:@24185.4]
  assign io_cdma2sc_dat_updt_valid = NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_valid; // @[NV_NVDLA_cdma.scala 436:25:@24442.4]
  assign io_cdma2sc_dat_updt_bits_entries = NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 436:25:@24441.4]
  assign io_cdma2sc_dat_updt_bits_slices = NV_NVDLA_CDMA_status_io_cdma2sc_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 436:25:@24440.4]
  assign io_cdma2sc_wt_updt_valid = NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_valid; // @[NV_NVDLA_cdma.scala 155:24:@24180.4]
  assign io_cdma2sc_wt_updt_bits_entries = NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_entries; // @[NV_NVDLA_cdma.scala 155:24:@24179.4]
  assign io_cdma2sc_wt_updt_bits_kernels = NV_NVDLA_CDMA_wt_io_cdma2sc_wt_updt_bits_kernels; // @[NV_NVDLA_cdma.scala 155:24:@24178.4]
  assign NV_NVDLA_CDMA_regfile_reset = io_nvdla_core_rstn; // @[:@24095.4]
  assign NV_NVDLA_CDMA_regfile_io_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 104:33:@24138.4]
  assign NV_NVDLA_CDMA_regfile_io_csb2cdma_req_valid = io_csb2cdma_req_valid; // @[NV_NVDLA_cdma.scala 106:27:@24142.4]
  assign NV_NVDLA_CDMA_regfile_io_csb2cdma_req_bits = io_csb2cdma_req_bits; // @[NV_NVDLA_cdma.scala 106:27:@24141.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_done = NV_NVDLA_CDMA_status_io_dp2reg_done; // @[NV_NVDLA_cdma.scala 123:30:@24155.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_latency = NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_latency; // @[NV_NVDLA_cdma.scala 109:39:@24145.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_dc_rd_stall = NV_NVDLA_CDMA_dc_io_dp2reg_dc_rd_stall; // @[NV_NVDLA_cdma.scala 108:37:@24144.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_latency = NV_NVDLA_CDMA_img_io_dp2reg_img_rd_latency; // @[NV_NVDLA_cdma.scala 112:40:@24147.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_img_rd_stall = NV_NVDLA_CDMA_img_io_dp2reg_img_rd_stall; // @[NV_NVDLA_cdma.scala 111:38:@24146.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_dat_flush_done = NV_NVDLA_CDMA_cvt_io_dp2reg_dat_flush_done; // @[NV_NVDLA_cdma.scala 127:40:@24158.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_wt_flush_done = NV_NVDLA_CDMA_wt_io_dp2reg_wt_flush_done; // @[NV_NVDLA_cdma.scala 119:39:@24152.4]
  assign NV_NVDLA_CDMA_regfile_io_dp2reg_wt_rd_stall = NV_NVDLA_CDMA_wt_io_dp2reg_wt_rd_stall; // @[NV_NVDLA_cdma.scala 120:37:@24153.4]
  assign NV_NVDLA_CDMA_wt_reset = io_nvdla_core_rstn; // @[:@24098.4]
  assign NV_NVDLA_CDMA_wt_io_nvdla_core_clk = NV_NVDLA_slcg_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 137:28:@24159.4]
  assign NV_NVDLA_CDMA_wt_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 138:31:@24160.4]
  assign NV_NVDLA_CDMA_wt_io_cdma_wt2mcif_rd_req_pd_ready = io_cdma_wt2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 142:31:@24164.4]
  assign NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_valid = io_mcif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 143:36:@24166.4]
  assign NV_NVDLA_CDMA_wt_io_mcif2cdma_wt_rd_rsp_pd_bits = io_mcif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 143:36:@24165.4]
  assign NV_NVDLA_CDMA_wt_io_cdma_wt2cvif_rd_req_pd_ready = io_cdma_wt2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 146:40:@24170.4]
  assign NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_valid = io_cvif2cdma_wt_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 147:44:@24172.4]
  assign NV_NVDLA_CDMA_wt_io_cvif2cdma_wt_rd_rsp_pd_bits = io_cvif2cdma_wt_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 147:44:@24171.4]
  assign NV_NVDLA_CDMA_wt_io_status2dma_fsm_switch = NV_NVDLA_CDMA_status_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 448:35:@24450.4]
  assign NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_valid = io_sc2cdma_wt_updt_valid; // @[NV_NVDLA_cdma.scala 156:29:@24183.4]
  assign NV_NVDLA_CDMA_wt_io_sc2cdma_wt_updt_bits_entries = io_sc2cdma_wt_updt_bits_entries; // @[NV_NVDLA_cdma.scala 156:29:@24182.4]
  assign NV_NVDLA_CDMA_wt_io_sc2cdma_wt_pending_req = io_sc2cdma_wt_pending_req; // @[NV_NVDLA_cdma.scala 158:36:@24184.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_op_en = NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 164:26:@24188.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_reuse = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_reuse; // @[NV_NVDLA_cdma.scala 166:33:@24190.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_skip_weight_rls = NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_weight_rls; // @[NV_NVDLA_cdma.scala 167:36:@24191.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_byte_per_kernel = NV_NVDLA_CDMA_regfile_io_reg2dp_field_byte_per_kernel; // @[NV_NVDLA_cdma.scala 169:36:@24193.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_kernel = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_kernel; // @[NV_NVDLA_cdma.scala 170:34:@24194.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_ram_type = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_ram_type; // @[NV_NVDLA_cdma.scala 171:36:@24195.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_low = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_low[31:5]; // @[NV_NVDLA_cdma.scala 172:36:@24197.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_addr_high = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_addr_high; // @[NV_NVDLA_cdma.scala 175:37:@24202.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_bytes = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bytes; // @[NV_NVDLA_cdma.scala 176:33:@24203.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_data_bank = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_cdma.scala 180:30:@24207.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_weight_bank = NV_NVDLA_CDMA_regfile_io_reg2dp_field_weight_bank; // @[NV_NVDLA_cdma.scala 181:32:@24208.4]
  assign NV_NVDLA_CDMA_wt_io_reg2dp_dma_en = NV_NVDLA_CDMA_regfile_io_reg2dp_field_dma_en; // @[NV_NVDLA_cdma.scala 183:27:@24210.4]
  assign NV_NVDLA_slcg_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 188:30:@24214.4]
  assign NV_NVDLA_CDMA_dc_reset = io_nvdla_core_rstn; // @[:@24104.4]
  assign NV_NVDLA_CDMA_dc_io_nvdla_core_clk = NV_NVDLA_slcg_1_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 194:28:@24217.4]
  assign NV_NVDLA_CDMA_dc_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 195:31:@24218.4]
  assign NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_ready = NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 198:40:@24222.4]
  assign NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_valid = NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 199:35:@24224.4]
  assign NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_bits = NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 199:35:@24223.4]
  assign NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_ready = NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 201:48:@24228.4]
  assign NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_valid = NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 202:43:@24230.4]
  assign NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_bits = NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 202:43:@24229.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_op_en = NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 223:26:@24252.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_conv_mode = NV_NVDLA_CDMA_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_cdma.scala 224:30:@24253.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_data_reuse = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_reuse; // @[NV_NVDLA_cdma.scala 225:31:@24254.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_skip_data_rls = NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_cdma.scala 226:34:@24255.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_format = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_cdma.scala 227:34:@24256.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_width = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_width; // @[NV_NVDLA_cdma.scala 228:33:@24257.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_height = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_height; // @[NV_NVDLA_cdma.scala 229:34:@24258.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_channel = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_channel; // @[NV_NVDLA_cdma.scala 230:35:@24259.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_ram_type = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_ram_type; // @[NV_NVDLA_cdma.scala 231:36:@24260.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_high_0 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_0; // @[NV_NVDLA_cdma.scala 232:39:@24261.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_datain_addr_low_0 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_0[26:0]; // @[NV_NVDLA_cdma.scala 233:38:@24263.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_line_stride = NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_stride[26:0]; // @[NV_NVDLA_cdma.scala 234:32:@24265.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_surf_stride = NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_stride[26:0]; // @[NV_NVDLA_cdma.scala 235:32:@24267.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_batch_stride = NV_NVDLA_CDMA_regfile_io_reg2dp_field_batch_stride[26:0]; // @[NV_NVDLA_cdma.scala 236:33:@24269.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_line_packed = NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_packed; // @[NV_NVDLA_cdma.scala 237:32:@24270.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_surf_packed = NV_NVDLA_CDMA_regfile_io_reg2dp_field_surf_packed; // @[NV_NVDLA_cdma.scala 238:32:@24271.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_batches = NV_NVDLA_CDMA_regfile_io_reg2dp_field_batches; // @[NV_NVDLA_cdma.scala 239:28:@24272.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_entries = {{3'd0}, NV_NVDLA_CDMA_regfile_io_reg2dp_field_entries}; // @[NV_NVDLA_cdma.scala 240:28:@24273.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_grains = NV_NVDLA_CDMA_regfile_io_reg2dp_field_grains; // @[NV_NVDLA_cdma.scala 241:27:@24274.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_data_bank = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_cdma.scala 242:30:@24275.4]
  assign NV_NVDLA_CDMA_dc_io_reg2dp_dma_en = NV_NVDLA_CDMA_regfile_io_reg2dp_field_dma_en; // @[NV_NVDLA_cdma.scala 243:27:@24276.4]
  assign NV_NVDLA_CDMA_dc_io_status2dma_fsm_switch = NV_NVDLA_CDMA_status_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 215:35:@24242.4]
  assign NV_NVDLA_CDMA_dc_io_status2dma_free_entries = NV_NVDLA_CDMA_status_io_status2dma_free_entries; // @[NV_NVDLA_cdma.scala 217:37:@24244.4]
  assign NV_NVDLA_CDMA_dc_io_status2dma_wr_idx = NV_NVDLA_CDMA_status_io_status2dma_wr_idx; // @[NV_NVDLA_cdma.scala 218:31:@24245.4]
  assign NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_data = NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_data; // @[NV_NVDLA_cdma.scala 221:40:@24249.4]
  assign NV_NVDLA_CDMA_dc_io_sc2cdma_dat_pending_req = io_sc2cdma_dat_pending_req; // @[NV_NVDLA_cdma.scala 205:37:@24232.4]
  assign NV_NVDLA_slcg_1_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 248:30:@24280.4]
  assign NV_NVDLA_CDMA_img_reset = io_nvdla_core_rstn; // @[:@24110.4]
  assign NV_NVDLA_CDMA_img_io_nvdla_core_clk = NV_NVDLA_slcg_2_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 263:29:@24285.4]
  assign NV_NVDLA_CDMA_img_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 264:32:@24286.4]
  assign NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_ready = NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 268:41:@24290.4]
  assign NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_valid = NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 269:37:@24292.4]
  assign NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_bits = NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 269:37:@24291.4]
  assign NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_ready = NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 271:49:@24296.4]
  assign NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_valid = NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 272:45:@24298.4]
  assign NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_bits = NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 272:45:@24297.4]
  assign NV_NVDLA_CDMA_img_io_status2dma_free_entries = NV_NVDLA_CDMA_status_io_status2dma_free_entries; // @[NV_NVDLA_cdma.scala 288:38:@24313.4]
  assign NV_NVDLA_CDMA_img_io_status2dma_wr_idx = NV_NVDLA_CDMA_status_io_status2dma_wr_idx; // @[NV_NVDLA_cdma.scala 289:32:@24314.4]
  assign NV_NVDLA_CDMA_img_io_status2dma_fsm_switch = NV_NVDLA_CDMA_status_io_status2dma_fsm_switch; // @[NV_NVDLA_cdma.scala 290:36:@24315.4]
  assign NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_data = NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_data; // @[NV_NVDLA_cdma.scala 293:41:@24319.4]
  assign NV_NVDLA_CDMA_img_io_sc2cdma_dat_pending_req = io_sc2cdma_dat_pending_req; // @[NV_NVDLA_cdma.scala 275:38:@24300.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_op_en = NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 295:27:@24322.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_conv_mode = NV_NVDLA_CDMA_regfile_io_reg2dp_field_conv_mode; // @[NV_NVDLA_cdma.scala 296:31:@24323.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_data_reuse = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_reuse; // @[NV_NVDLA_cdma.scala 299:32:@24326.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_skip_data_rls = NV_NVDLA_CDMA_regfile_io_reg2dp_field_skip_data_rls; // @[NV_NVDLA_cdma.scala 300:35:@24327.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_format = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_format; // @[NV_NVDLA_cdma.scala 301:35:@24328.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_pixel_format = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_format; // @[NV_NVDLA_cdma.scala 302:34:@24329.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_pixel_sign_override = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_sign_override; // @[NV_NVDLA_cdma.scala 304:41:@24331.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_width = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_width; // @[NV_NVDLA_cdma.scala 305:34:@24332.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_height = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_height; // @[NV_NVDLA_cdma.scala 306:35:@24333.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_channel = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_channel; // @[NV_NVDLA_cdma.scala 307:36:@24334.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_pixel_x_offset = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pixel_x_offset; // @[NV_NVDLA_cdma.scala 308:36:@24335.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_ram_type = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_ram_type; // @[NV_NVDLA_cdma.scala 310:37:@24337.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_0 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_0; // @[NV_NVDLA_cdma.scala 311:40:@24338.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_0 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_0; // @[NV_NVDLA_cdma.scala 312:39:@24339.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_low_1 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_low_1; // @[NV_NVDLA_cdma.scala 313:39:@24340.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_line_stride = NV_NVDLA_CDMA_regfile_io_reg2dp_field_line_stride; // @[NV_NVDLA_cdma.scala 314:33:@24341.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_uv_line_stride = NV_NVDLA_CDMA_regfile_io_reg2dp_field_uv_line_stride; // @[NV_NVDLA_cdma.scala 315:36:@24342.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_datain_addr_high_1 = NV_NVDLA_CDMA_regfile_io_reg2dp_field_datain_addr_high_1; // @[NV_NVDLA_cdma.scala 316:40:@24343.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_mean_format = NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_format; // @[NV_NVDLA_cdma.scala 317:33:@24344.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_mean_ry = NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ry; // @[NV_NVDLA_cdma.scala 318:29:@24345.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_mean_gu = NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_gu; // @[NV_NVDLA_cdma.scala 319:29:@24346.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_mean_bv = NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_bv; // @[NV_NVDLA_cdma.scala 320:29:@24347.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_mean_ax = NV_NVDLA_CDMA_regfile_io_reg2dp_field_mean_ax; // @[NV_NVDLA_cdma.scala 321:29:@24348.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_entries = NV_NVDLA_CDMA_regfile_io_reg2dp_field_entries; // @[NV_NVDLA_cdma.scala 322:29:@24349.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_pad_left = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_left; // @[NV_NVDLA_cdma.scala 323:30:@24350.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_pad_right = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_right; // @[NV_NVDLA_cdma.scala 324:31:@24351.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_data_bank = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_cdma.scala 325:31:@24352.4]
  assign NV_NVDLA_CDMA_img_io_reg2dp_dma_en = NV_NVDLA_CDMA_regfile_io_reg2dp_field_dma_en; // @[NV_NVDLA_cdma.scala 326:28:@24353.4]
  assign NV_NVDLA_slcg_2_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 338:31:@24361.4]
  assign NV_NVDLA_CDMA_dma_mux_reset = io_nvdla_core_rstn; // @[:@24116.4]
  assign NV_NVDLA_CDMA_dma_mux_io_nvdla_core_clk = NV_NVDLA_slcg_3_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 348:33:@24366.4]
  assign NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_valid = NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 198:40:@24221.4]
  assign NV_NVDLA_CDMA_dma_mux_io_dc_dat2mcif_rd_req_pd_bits = NV_NVDLA_CDMA_dc_io_dc_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 198:40:@24220.4]
  assign NV_NVDLA_CDMA_dma_mux_io_mcif2dc_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_dc_io_mcif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 199:35:@24225.4]
  assign NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_valid = NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 268:41:@24289.4]
  assign NV_NVDLA_CDMA_dma_mux_io_img_dat2mcif_rd_req_pd_bits = NV_NVDLA_CDMA_img_io_img_dat2mcif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 268:41:@24288.4]
  assign NV_NVDLA_CDMA_dma_mux_io_mcif2img_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_img_io_mcif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 269:37:@24293.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cdma_dat2mcif_rd_req_pd_ready = io_cdma_dat2mcif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 350:32:@24369.4]
  assign NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_valid = io_mcif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 351:42:@24371.4]
  assign NV_NVDLA_CDMA_dma_mux_io_mcif2cdma_dat_rd_rsp_pd_bits = io_mcif2cdma_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 351:42:@24370.4]
  assign NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_valid = NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 201:48:@24227.4]
  assign NV_NVDLA_CDMA_dma_mux_io_dc_dat2cvif_rd_req_pd_bits = NV_NVDLA_CDMA_dc_io_dc_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 201:48:@24226.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cvif2dc_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_dc_io_cvif2dc_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 202:43:@24231.4]
  assign NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_valid = NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_valid; // @[NV_NVDLA_cdma.scala 271:49:@24295.4]
  assign NV_NVDLA_CDMA_dma_mux_io_img_dat2cvif_rd_req_pd_bits = NV_NVDLA_CDMA_img_io_img_dat2cvif_rd_req_pd_bits; // @[NV_NVDLA_cdma.scala 271:49:@24294.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cvif2img_dat_rd_rsp_pd_ready = NV_NVDLA_CDMA_img_io_cvif2img_dat_rd_rsp_pd_ready; // @[NV_NVDLA_cdma.scala 272:45:@24299.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cdma_dat2cvif_rd_req_pd_ready = io_cdma_dat2cvif_rd_req_pd_ready; // @[NV_NVDLA_cdma.scala 354:40:@24375.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_valid = io_cvif2cdma_dat_rd_rsp_pd_valid; // @[NV_NVDLA_cdma.scala 355:50:@24377.4]
  assign NV_NVDLA_CDMA_dma_mux_io_cvif2cdma_dat_rd_rsp_pd_bits = io_cvif2cdma_dat_rd_rsp_pd_bits; // @[NV_NVDLA_cdma.scala 355:50:@24376.4]
  assign NV_NVDLA_slcg_3_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 361:31:@24382.4]
  assign NV_NVDLA_CDMA_cvt_reset = io_nvdla_core_rstn; // @[:@24122.4]
  assign NV_NVDLA_CDMA_cvt_io_nvdla_core_clk = NV_NVDLA_slcg_4_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 367:29:@24385.4]
  assign NV_NVDLA_CDMA_cvt_io_nvdla_core_ng_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 369:32:@24387.4]
  assign NV_NVDLA_CDMA_cvt_io_nvdla_hls_clk = NV_NVDLA_slcg_5_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 368:28:@24386.4]
  assign NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_sel = NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 208:40:@24233.4]
  assign NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_valid = NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 210:28:@24236.4]
  assign NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_addr_bits = NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 210:28:@24235.4]
  assign NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_data = NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 210:28:@24234.4]
  assign NV_NVDLA_CDMA_cvt_io_dc2cvt_dat_wr_info_pd = NV_NVDLA_CDMA_dc_io_dc2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 211:36:@24237.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_sel = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_sel; // @[NV_NVDLA_cdma.scala 278:41:@24301.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_valid = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_valid; // @[NV_NVDLA_cdma.scala 280:29:@24304.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_addr_bits = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_addr_bits; // @[NV_NVDLA_cdma.scala 280:29:@24303.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_data = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_data; // @[NV_NVDLA_cdma.scala 280:29:@24302.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_mn_wr_data = NV_NVDLA_CDMA_img_io_img2cvt_mn_wr_data; // @[NV_NVDLA_cdma.scala 281:33:@24305.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_pad_mask = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_pad_mask; // @[NV_NVDLA_cdma.scala 282:38:@24306.4]
  assign NV_NVDLA_CDMA_cvt_io_img2cvt_dat_wr_info_pd = NV_NVDLA_CDMA_img_io_img2cvt_dat_wr_info_pd; // @[NV_NVDLA_cdma.scala 283:37:@24307.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_op_en = NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 378:27:@24392.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_proc_precision = NV_NVDLA_CDMA_regfile_io_reg2dp_field_proc_precision; // @[NV_NVDLA_cdma.scala 380:36:@24394.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_en = NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_en; // @[NV_NVDLA_cdma.scala 381:28:@24395.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_truncate = NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_truncate; // @[NV_NVDLA_cdma.scala 382:34:@24396.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_offset = NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_offset; // @[NV_NVDLA_cdma.scala 383:32:@24397.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_cvt_scale = NV_NVDLA_CDMA_regfile_io_reg2dp_field_cvt_scale; // @[NV_NVDLA_cdma.scala 384:31:@24398.4]
  assign NV_NVDLA_CDMA_cvt_io_reg2dp_pad_value = NV_NVDLA_CDMA_regfile_io_reg2dp_field_pad_value; // @[NV_NVDLA_cdma.scala 386:31:@24400.4]
  assign NV_NVDLA_CDMA_cvt_io_dp2reg_done = NV_NVDLA_CDMA_status_io_dp2reg_done; // @[NV_NVDLA_cdma.scala 387:26:@24401.4]
  assign NV_NVDLA_slcg_4_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 392:31:@24405.4]
  assign NV_NVDLA_slcg_5_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 399:31:@24411.4]
  assign NV_NVDLA_CDMA_shared_buffer_reset = io_nvdla_core_rstn; // @[:@24131.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_nvdla_core_clk = NV_NVDLA_slcg_6_io_nvdla_core_gated_clk; // @[NV_NVDLA_cdma.scala 407:39:@24415.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_valid = NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_cdma.scala 220:40:@24248.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_addr_bits = NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_addr_bits; // @[NV_NVDLA_cdma.scala 220:40:@24247.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_wr_0_data = NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_wr_data; // @[NV_NVDLA_cdma.scala 220:40:@24246.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_valid = NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_valid; // @[NV_NVDLA_cdma.scala 292:41:@24318.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_addr_bits = NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_addr_bits; // @[NV_NVDLA_cdma.scala 292:41:@24317.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_wr_0_data = NV_NVDLA_CDMA_img_io_img2sbuf_p0_wr_data; // @[NV_NVDLA_cdma.scala 292:41:@24316.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_valid = NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_cdma.scala 221:40:@24251.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_dc2sbuf_p_rd_0_addr_bits = NV_NVDLA_CDMA_dc_io_dc2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_cdma.scala 221:40:@24250.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_valid = NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_valid; // @[NV_NVDLA_cdma.scala 293:41:@24321.4]
  assign NV_NVDLA_CDMA_shared_buffer_io_img2sbuf_p_rd_0_addr_bits = NV_NVDLA_CDMA_img_io_img2sbuf_p0_rd_addr_bits; // @[NV_NVDLA_cdma.scala 293:41:@24320.4]
  assign NV_NVDLA_slcg_6_io_nvdla_clock_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 425:34:@24430.4]
  assign NV_NVDLA_CDMA_status_reset = io_nvdla_core_rstn; // @[:@24137.4]
  assign NV_NVDLA_CDMA_status_io_nvdla_core_clk = io_nvdla_clock_nvdla_core_clk; // @[NV_NVDLA_cdma.scala 431:32:@24433.4]
  assign NV_NVDLA_CDMA_status_io_dc2status_dat_updt_valid = NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 214:36:@24241.4 NV_NVDLA_cdma.scala 433:36:@24436.4]
  assign NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_entries = NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 214:36:@24240.4 NV_NVDLA_cdma.scala 433:36:@24435.4]
  assign NV_NVDLA_CDMA_status_io_dc2status_dat_updt_bits_slices = NV_NVDLA_CDMA_dc_io_dc2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 214:36:@24239.4 NV_NVDLA_cdma.scala 433:36:@24434.4]
  assign NV_NVDLA_CDMA_status_io_img2status_dat_updt_valid = NV_NVDLA_CDMA_img_io_img2status_dat_updt_valid; // @[NV_NVDLA_cdma.scala 286:37:@24311.4]
  assign NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_entries = NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 286:37:@24310.4]
  assign NV_NVDLA_CDMA_status_io_img2status_dat_updt_bits_slices = NV_NVDLA_CDMA_img_io_img2status_dat_updt_bits_slices; // @[NV_NVDLA_cdma.scala 286:37:@24309.4]
  assign NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_valid = io_sc2cdma_dat_updt_valid; // @[NV_NVDLA_cdma.scala 435:34:@24439.4]
  assign NV_NVDLA_CDMA_status_io_sc2cdma_dat_updt_bits_entries = io_sc2cdma_dat_updt_bits_entries; // @[NV_NVDLA_cdma.scala 435:34:@24438.4]
  assign NV_NVDLA_CDMA_status_io_dc2status_state = NV_NVDLA_CDMA_dc_io_dc2status_state; // @[NV_NVDLA_cdma.scala 213:33:@24238.4]
  assign NV_NVDLA_CDMA_status_io_img2status_state = NV_NVDLA_CDMA_img_io_img2status_state; // @[NV_NVDLA_cdma.scala 285:34:@24308.4]
  assign NV_NVDLA_CDMA_status_io_wt2status_state = NV_NVDLA_CDMA_wt_io_wt2status_state; // @[NV_NVDLA_cdma.scala 449:33:@24451.4]
  assign NV_NVDLA_CDMA_status_io_dp2reg_consumer = NV_NVDLA_CDMA_regfile_io_dp2reg_consumer; // @[NV_NVDLA_cdma.scala 446:33:@24449.4]
  assign NV_NVDLA_CDMA_status_io_reg2dp_op_en = NV_NVDLA_CDMA_regfile_io_reg2dp_op_en; // @[NV_NVDLA_cdma.scala 444:30:@24447.4]
  assign NV_NVDLA_CDMA_status_io_reg2dp_data_bank = NV_NVDLA_CDMA_regfile_io_reg2dp_field_data_bank; // @[NV_NVDLA_cdma.scala 445:34:@24448.4]
  assign NV_NVDLA_CDMA_status_io_sc2cdma_dat_pending_req = {{1'd0}, io_sc2cdma_dat_pending_req}; // @[NV_NVDLA_cdma.scala 441:41:@24445.4]
endmodule
