// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CMAC_CORE_active_gold.v
// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CMAC.h
module NV_NVDLA_CMAC_CORE_active_gold (
   nvdla_core_clk
  ,nvdla_core_rstn
//: for(my $i=0; $i<64; $i++){
//: print qq(
//: ,in_dat_data${i})
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,in_dat_data0
,in_dat_data1
,in_dat_data2
,in_dat_data3
,in_dat_data4
,in_dat_data5
,in_dat_data6
,in_dat_data7
,in_dat_data8
,in_dat_data9
,in_dat_data10
,in_dat_data11
,in_dat_data12
,in_dat_data13
,in_dat_data14
,in_dat_data15
,in_dat_data16
,in_dat_data17
,in_dat_data18
,in_dat_data19
,in_dat_data20
,in_dat_data21
,in_dat_data22
,in_dat_data23
,in_dat_data24
,in_dat_data25
,in_dat_data26
,in_dat_data27
,in_dat_data28
,in_dat_data29
,in_dat_data30
,in_dat_data31
,in_dat_data32
,in_dat_data33
,in_dat_data34
,in_dat_data35
,in_dat_data36
,in_dat_data37
,in_dat_data38
,in_dat_data39
,in_dat_data40
,in_dat_data41
,in_dat_data42
,in_dat_data43
,in_dat_data44
,in_dat_data45
,in_dat_data46
,in_dat_data47
,in_dat_data48
,in_dat_data49
,in_dat_data50
,in_dat_data51
,in_dat_data52
,in_dat_data53
,in_dat_data54
,in_dat_data55
,in_dat_data56
,in_dat_data57
,in_dat_data58
,in_dat_data59
,in_dat_data60
,in_dat_data61
,in_dat_data62
,in_dat_data63
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,in_dat_mask
  ,in_dat_pvld
  ,in_dat_stripe_end
  ,in_dat_stripe_st
//: for(my $i=0; $i<64; $i++){
//: print qq(
//: ,in_wt_data${i})
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,in_wt_data0
,in_wt_data1
,in_wt_data2
,in_wt_data3
,in_wt_data4
,in_wt_data5
,in_wt_data6
,in_wt_data7
,in_wt_data8
,in_wt_data9
,in_wt_data10
,in_wt_data11
,in_wt_data12
,in_wt_data13
,in_wt_data14
,in_wt_data15
,in_wt_data16
,in_wt_data17
,in_wt_data18
,in_wt_data19
,in_wt_data20
,in_wt_data21
,in_wt_data22
,in_wt_data23
,in_wt_data24
,in_wt_data25
,in_wt_data26
,in_wt_data27
,in_wt_data28
,in_wt_data29
,in_wt_data30
,in_wt_data31
,in_wt_data32
,in_wt_data33
,in_wt_data34
,in_wt_data35
,in_wt_data36
,in_wt_data37
,in_wt_data38
,in_wt_data39
,in_wt_data40
,in_wt_data41
,in_wt_data42
,in_wt_data43
,in_wt_data44
,in_wt_data45
,in_wt_data46
,in_wt_data47
,in_wt_data48
,in_wt_data49
,in_wt_data50
,in_wt_data51
,in_wt_data52
,in_wt_data53
,in_wt_data54
,in_wt_data55
,in_wt_data56
,in_wt_data57
,in_wt_data58
,in_wt_data59
,in_wt_data60
,in_wt_data61
,in_wt_data62
,in_wt_data63
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,in_wt_mask
  ,in_wt_pvld
  ,in_wt_sel
//: for(my $i=0; $i<32/2; $i++){
//: print qq(
//: ,dat${i}_actv_data
//: ,dat${i}_actv_nz
//: ,dat${i}_actv_pvld
//: ,dat${i}_pre_mask
//: ,dat${i}_pre_pvld
//: ,dat${i}_pre_stripe_end
//: ,dat${i}_pre_stripe_st
//: )
//: }
//: for(my $i=0; $i<32/2; $i++){
//: print qq(
//: ,wt${i}_actv_data
//: ,wt${i}_actv_nz
//: ,wt${i}_actv_pvld
//: ,wt${i}_sd_mask
//: ,wt${i}_sd_pvld
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,dat0_actv_data
,dat0_actv_nz
,dat0_actv_pvld
,dat0_pre_mask
,dat0_pre_pvld
,dat0_pre_stripe_end
,dat0_pre_stripe_st

,dat1_actv_data
,dat1_actv_nz
,dat1_actv_pvld
,dat1_pre_mask
,dat1_pre_pvld
,dat1_pre_stripe_end
,dat1_pre_stripe_st

,dat2_actv_data
,dat2_actv_nz
,dat2_actv_pvld
,dat2_pre_mask
,dat2_pre_pvld
,dat2_pre_stripe_end
,dat2_pre_stripe_st

,dat3_actv_data
,dat3_actv_nz
,dat3_actv_pvld
,dat3_pre_mask
,dat3_pre_pvld
,dat3_pre_stripe_end
,dat3_pre_stripe_st

,dat4_actv_data
,dat4_actv_nz
,dat4_actv_pvld
,dat4_pre_mask
,dat4_pre_pvld
,dat4_pre_stripe_end
,dat4_pre_stripe_st

,dat5_actv_data
,dat5_actv_nz
,dat5_actv_pvld
,dat5_pre_mask
,dat5_pre_pvld
,dat5_pre_stripe_end
,dat5_pre_stripe_st

,dat6_actv_data
,dat6_actv_nz
,dat6_actv_pvld
,dat6_pre_mask
,dat6_pre_pvld
,dat6_pre_stripe_end
,dat6_pre_stripe_st

,dat7_actv_data
,dat7_actv_nz
,dat7_actv_pvld
,dat7_pre_mask
,dat7_pre_pvld
,dat7_pre_stripe_end
,dat7_pre_stripe_st

,dat8_actv_data
,dat8_actv_nz
,dat8_actv_pvld
,dat8_pre_mask
,dat8_pre_pvld
,dat8_pre_stripe_end
,dat8_pre_stripe_st

,dat9_actv_data
,dat9_actv_nz
,dat9_actv_pvld
,dat9_pre_mask
,dat9_pre_pvld
,dat9_pre_stripe_end
,dat9_pre_stripe_st

,dat10_actv_data
,dat10_actv_nz
,dat10_actv_pvld
,dat10_pre_mask
,dat10_pre_pvld
,dat10_pre_stripe_end
,dat10_pre_stripe_st

,dat11_actv_data
,dat11_actv_nz
,dat11_actv_pvld
,dat11_pre_mask
,dat11_pre_pvld
,dat11_pre_stripe_end
,dat11_pre_stripe_st

,dat12_actv_data
,dat12_actv_nz
,dat12_actv_pvld
,dat12_pre_mask
,dat12_pre_pvld
,dat12_pre_stripe_end
,dat12_pre_stripe_st

,dat13_actv_data
,dat13_actv_nz
,dat13_actv_pvld
,dat13_pre_mask
,dat13_pre_pvld
,dat13_pre_stripe_end
,dat13_pre_stripe_st

,dat14_actv_data
,dat14_actv_nz
,dat14_actv_pvld
,dat14_pre_mask
,dat14_pre_pvld
,dat14_pre_stripe_end
,dat14_pre_stripe_st

,dat15_actv_data
,dat15_actv_nz
,dat15_actv_pvld
,dat15_pre_mask
,dat15_pre_pvld
,dat15_pre_stripe_end
,dat15_pre_stripe_st

,wt0_actv_data
,wt0_actv_nz
,wt0_actv_pvld
,wt0_sd_mask
,wt0_sd_pvld

,wt1_actv_data
,wt1_actv_nz
,wt1_actv_pvld
,wt1_sd_mask
,wt1_sd_pvld

,wt2_actv_data
,wt2_actv_nz
,wt2_actv_pvld
,wt2_sd_mask
,wt2_sd_pvld

,wt3_actv_data
,wt3_actv_nz
,wt3_actv_pvld
,wt3_sd_mask
,wt3_sd_pvld

,wt4_actv_data
,wt4_actv_nz
,wt4_actv_pvld
,wt4_sd_mask
,wt4_sd_pvld

,wt5_actv_data
,wt5_actv_nz
,wt5_actv_pvld
,wt5_sd_mask
,wt5_sd_pvld

,wt6_actv_data
,wt6_actv_nz
,wt6_actv_pvld
,wt6_sd_mask
,wt6_sd_pvld

,wt7_actv_data
,wt7_actv_nz
,wt7_actv_pvld
,wt7_sd_mask
,wt7_sd_pvld

,wt8_actv_data
,wt8_actv_nz
,wt8_actv_pvld
,wt8_sd_mask
,wt8_sd_pvld

,wt9_actv_data
,wt9_actv_nz
,wt9_actv_pvld
,wt9_sd_mask
,wt9_sd_pvld

,wt10_actv_data
,wt10_actv_nz
,wt10_actv_pvld
,wt10_sd_mask
,wt10_sd_pvld

,wt11_actv_data
,wt11_actv_nz
,wt11_actv_pvld
,wt11_sd_mask
,wt11_sd_pvld

,wt12_actv_data
,wt12_actv_nz
,wt12_actv_pvld
,wt12_sd_mask
,wt12_sd_pvld

,wt13_actv_data
,wt13_actv_nz
,wt13_actv_pvld
,wt13_sd_mask
,wt13_sd_pvld

,wt14_actv_data
,wt14_actv_nz
,wt14_actv_pvld
,wt14_sd_mask
,wt14_sd_pvld

,wt15_actv_data
,wt15_actv_nz
,wt15_actv_pvld
,wt15_sd_mask
,wt15_sd_pvld

//| eperl: generated_end (DO NOT EDIT ABOVE)
  );
input nvdla_core_clk;
input nvdla_core_rstn;
//: for(my $i=0; $i<64; $i++){
//: print qq(
//: input [8 -1:0] in_dat_data${i};)
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

input [8 -1:0] in_dat_data0;
input [8 -1:0] in_dat_data1;
input [8 -1:0] in_dat_data2;
input [8 -1:0] in_dat_data3;
input [8 -1:0] in_dat_data4;
input [8 -1:0] in_dat_data5;
input [8 -1:0] in_dat_data6;
input [8 -1:0] in_dat_data7;
input [8 -1:0] in_dat_data8;
input [8 -1:0] in_dat_data9;
input [8 -1:0] in_dat_data10;
input [8 -1:0] in_dat_data11;
input [8 -1:0] in_dat_data12;
input [8 -1:0] in_dat_data13;
input [8 -1:0] in_dat_data14;
input [8 -1:0] in_dat_data15;
input [8 -1:0] in_dat_data16;
input [8 -1:0] in_dat_data17;
input [8 -1:0] in_dat_data18;
input [8 -1:0] in_dat_data19;
input [8 -1:0] in_dat_data20;
input [8 -1:0] in_dat_data21;
input [8 -1:0] in_dat_data22;
input [8 -1:0] in_dat_data23;
input [8 -1:0] in_dat_data24;
input [8 -1:0] in_dat_data25;
input [8 -1:0] in_dat_data26;
input [8 -1:0] in_dat_data27;
input [8 -1:0] in_dat_data28;
input [8 -1:0] in_dat_data29;
input [8 -1:0] in_dat_data30;
input [8 -1:0] in_dat_data31;
input [8 -1:0] in_dat_data32;
input [8 -1:0] in_dat_data33;
input [8 -1:0] in_dat_data34;
input [8 -1:0] in_dat_data35;
input [8 -1:0] in_dat_data36;
input [8 -1:0] in_dat_data37;
input [8 -1:0] in_dat_data38;
input [8 -1:0] in_dat_data39;
input [8 -1:0] in_dat_data40;
input [8 -1:0] in_dat_data41;
input [8 -1:0] in_dat_data42;
input [8 -1:0] in_dat_data43;
input [8 -1:0] in_dat_data44;
input [8 -1:0] in_dat_data45;
input [8 -1:0] in_dat_data46;
input [8 -1:0] in_dat_data47;
input [8 -1:0] in_dat_data48;
input [8 -1:0] in_dat_data49;
input [8 -1:0] in_dat_data50;
input [8 -1:0] in_dat_data51;
input [8 -1:0] in_dat_data52;
input [8 -1:0] in_dat_data53;
input [8 -1:0] in_dat_data54;
input [8 -1:0] in_dat_data55;
input [8 -1:0] in_dat_data56;
input [8 -1:0] in_dat_data57;
input [8 -1:0] in_dat_data58;
input [8 -1:0] in_dat_data59;
input [8 -1:0] in_dat_data60;
input [8 -1:0] in_dat_data61;
input [8 -1:0] in_dat_data62;
input [8 -1:0] in_dat_data63;
//| eperl: generated_end (DO NOT EDIT ABOVE)
input [64 -1:0] in_dat_mask;
input in_dat_pvld;
input in_dat_stripe_end;
input in_dat_stripe_st;
//: for(my $i=0; $i<64; $i++){
//: print qq(
//: input [8 -1:0] in_wt_data${i};)
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

input [8 -1:0] in_wt_data0;
input [8 -1:0] in_wt_data1;
input [8 -1:0] in_wt_data2;
input [8 -1:0] in_wt_data3;
input [8 -1:0] in_wt_data4;
input [8 -1:0] in_wt_data5;
input [8 -1:0] in_wt_data6;
input [8 -1:0] in_wt_data7;
input [8 -1:0] in_wt_data8;
input [8 -1:0] in_wt_data9;
input [8 -1:0] in_wt_data10;
input [8 -1:0] in_wt_data11;
input [8 -1:0] in_wt_data12;
input [8 -1:0] in_wt_data13;
input [8 -1:0] in_wt_data14;
input [8 -1:0] in_wt_data15;
input [8 -1:0] in_wt_data16;
input [8 -1:0] in_wt_data17;
input [8 -1:0] in_wt_data18;
input [8 -1:0] in_wt_data19;
input [8 -1:0] in_wt_data20;
input [8 -1:0] in_wt_data21;
input [8 -1:0] in_wt_data22;
input [8 -1:0] in_wt_data23;
input [8 -1:0] in_wt_data24;
input [8 -1:0] in_wt_data25;
input [8 -1:0] in_wt_data26;
input [8 -1:0] in_wt_data27;
input [8 -1:0] in_wt_data28;
input [8 -1:0] in_wt_data29;
input [8 -1:0] in_wt_data30;
input [8 -1:0] in_wt_data31;
input [8 -1:0] in_wt_data32;
input [8 -1:0] in_wt_data33;
input [8 -1:0] in_wt_data34;
input [8 -1:0] in_wt_data35;
input [8 -1:0] in_wt_data36;
input [8 -1:0] in_wt_data37;
input [8 -1:0] in_wt_data38;
input [8 -1:0] in_wt_data39;
input [8 -1:0] in_wt_data40;
input [8 -1:0] in_wt_data41;
input [8 -1:0] in_wt_data42;
input [8 -1:0] in_wt_data43;
input [8 -1:0] in_wt_data44;
input [8 -1:0] in_wt_data45;
input [8 -1:0] in_wt_data46;
input [8 -1:0] in_wt_data47;
input [8 -1:0] in_wt_data48;
input [8 -1:0] in_wt_data49;
input [8 -1:0] in_wt_data50;
input [8 -1:0] in_wt_data51;
input [8 -1:0] in_wt_data52;
input [8 -1:0] in_wt_data53;
input [8 -1:0] in_wt_data54;
input [8 -1:0] in_wt_data55;
input [8 -1:0] in_wt_data56;
input [8 -1:0] in_wt_data57;
input [8 -1:0] in_wt_data58;
input [8 -1:0] in_wt_data59;
input [8 -1:0] in_wt_data60;
input [8 -1:0] in_wt_data61;
input [8 -1:0] in_wt_data62;
input [8 -1:0] in_wt_data63;
//| eperl: generated_end (DO NOT EDIT ABOVE)
input [64 -1:0] in_wt_mask;
input in_wt_pvld;
input [32/2 -1:0] in_wt_sel;
//: for(my $i=0; $i<32/2; $i++){
//: print qq(
//: output [8*64 -1:0] dat${i}_actv_data;
//: output [64 -1:0] dat${i}_actv_nz;
//: output [64 -1:0] dat${i}_actv_pvld;
//: output [64 -1:0] dat${i}_pre_mask;
//: output dat${i}_pre_pvld;
//: output dat${i}_pre_stripe_end;
//: output dat${i}_pre_stripe_st;
//: )
//: }
//: for(my $i=0; $i<32/2; $i++){
//: print qq(
//: output [8*64 -1:0] wt${i}_actv_data;
//: output [64 -1:0] wt${i}_actv_nz;
//: output [64 -1:0] wt${i}_actv_pvld;
//: output [64 -1:0] wt${i}_sd_mask;
//: output wt${i}_sd_pvld;
//: )
//: }
//: for(my $i=0; $i<32/2; $i++){
//: print qq(
//: reg [8*64 -1:0] dat_actv_data_reg${i};
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

output [8*64 -1:0] dat0_actv_data;
output [64 -1:0] dat0_actv_nz;
output [64 -1:0] dat0_actv_pvld;
output [64 -1:0] dat0_pre_mask;
output dat0_pre_pvld;
output dat0_pre_stripe_end;
output dat0_pre_stripe_st;

output [8*64 -1:0] dat1_actv_data;
output [64 -1:0] dat1_actv_nz;
output [64 -1:0] dat1_actv_pvld;
output [64 -1:0] dat1_pre_mask;
output dat1_pre_pvld;
output dat1_pre_stripe_end;
output dat1_pre_stripe_st;

output [8*64 -1:0] dat2_actv_data;
output [64 -1:0] dat2_actv_nz;
output [64 -1:0] dat2_actv_pvld;
output [64 -1:0] dat2_pre_mask;
output dat2_pre_pvld;
output dat2_pre_stripe_end;
output dat2_pre_stripe_st;

output [8*64 -1:0] dat3_actv_data;
output [64 -1:0] dat3_actv_nz;
output [64 -1:0] dat3_actv_pvld;
output [64 -1:0] dat3_pre_mask;
output dat3_pre_pvld;
output dat3_pre_stripe_end;
output dat3_pre_stripe_st;

output [8*64 -1:0] dat4_actv_data;
output [64 -1:0] dat4_actv_nz;
output [64 -1:0] dat4_actv_pvld;
output [64 -1:0] dat4_pre_mask;
output dat4_pre_pvld;
output dat4_pre_stripe_end;
output dat4_pre_stripe_st;

output [8*64 -1:0] dat5_actv_data;
output [64 -1:0] dat5_actv_nz;
output [64 -1:0] dat5_actv_pvld;
output [64 -1:0] dat5_pre_mask;
output dat5_pre_pvld;
output dat5_pre_stripe_end;
output dat5_pre_stripe_st;

output [8*64 -1:0] dat6_actv_data;
output [64 -1:0] dat6_actv_nz;
output [64 -1:0] dat6_actv_pvld;
output [64 -1:0] dat6_pre_mask;
output dat6_pre_pvld;
output dat6_pre_stripe_end;
output dat6_pre_stripe_st;

output [8*64 -1:0] dat7_actv_data;
output [64 -1:0] dat7_actv_nz;
output [64 -1:0] dat7_actv_pvld;
output [64 -1:0] dat7_pre_mask;
output dat7_pre_pvld;
output dat7_pre_stripe_end;
output dat7_pre_stripe_st;

output [8*64 -1:0] dat8_actv_data;
output [64 -1:0] dat8_actv_nz;
output [64 -1:0] dat8_actv_pvld;
output [64 -1:0] dat8_pre_mask;
output dat8_pre_pvld;
output dat8_pre_stripe_end;
output dat8_pre_stripe_st;

output [8*64 -1:0] dat9_actv_data;
output [64 -1:0] dat9_actv_nz;
output [64 -1:0] dat9_actv_pvld;
output [64 -1:0] dat9_pre_mask;
output dat9_pre_pvld;
output dat9_pre_stripe_end;
output dat9_pre_stripe_st;

output [8*64 -1:0] dat10_actv_data;
output [64 -1:0] dat10_actv_nz;
output [64 -1:0] dat10_actv_pvld;
output [64 -1:0] dat10_pre_mask;
output dat10_pre_pvld;
output dat10_pre_stripe_end;
output dat10_pre_stripe_st;

output [8*64 -1:0] dat11_actv_data;
output [64 -1:0] dat11_actv_nz;
output [64 -1:0] dat11_actv_pvld;
output [64 -1:0] dat11_pre_mask;
output dat11_pre_pvld;
output dat11_pre_stripe_end;
output dat11_pre_stripe_st;

output [8*64 -1:0] dat12_actv_data;
output [64 -1:0] dat12_actv_nz;
output [64 -1:0] dat12_actv_pvld;
output [64 -1:0] dat12_pre_mask;
output dat12_pre_pvld;
output dat12_pre_stripe_end;
output dat12_pre_stripe_st;

output [8*64 -1:0] dat13_actv_data;
output [64 -1:0] dat13_actv_nz;
output [64 -1:0] dat13_actv_pvld;
output [64 -1:0] dat13_pre_mask;
output dat13_pre_pvld;
output dat13_pre_stripe_end;
output dat13_pre_stripe_st;

output [8*64 -1:0] dat14_actv_data;
output [64 -1:0] dat14_actv_nz;
output [64 -1:0] dat14_actv_pvld;
output [64 -1:0] dat14_pre_mask;
output dat14_pre_pvld;
output dat14_pre_stripe_end;
output dat14_pre_stripe_st;

output [8*64 -1:0] dat15_actv_data;
output [64 -1:0] dat15_actv_nz;
output [64 -1:0] dat15_actv_pvld;
output [64 -1:0] dat15_pre_mask;
output dat15_pre_pvld;
output dat15_pre_stripe_end;
output dat15_pre_stripe_st;

output [8*64 -1:0] wt0_actv_data;
output [64 -1:0] wt0_actv_nz;
output [64 -1:0] wt0_actv_pvld;
output [64 -1:0] wt0_sd_mask;
output wt0_sd_pvld;

output [8*64 -1:0] wt1_actv_data;
output [64 -1:0] wt1_actv_nz;
output [64 -1:0] wt1_actv_pvld;
output [64 -1:0] wt1_sd_mask;
output wt1_sd_pvld;

output [8*64 -1:0] wt2_actv_data;
output [64 -1:0] wt2_actv_nz;
output [64 -1:0] wt2_actv_pvld;
output [64 -1:0] wt2_sd_mask;
output wt2_sd_pvld;

output [8*64 -1:0] wt3_actv_data;
output [64 -1:0] wt3_actv_nz;
output [64 -1:0] wt3_actv_pvld;
output [64 -1:0] wt3_sd_mask;
output wt3_sd_pvld;

output [8*64 -1:0] wt4_actv_data;
output [64 -1:0] wt4_actv_nz;
output [64 -1:0] wt4_actv_pvld;
output [64 -1:0] wt4_sd_mask;
output wt4_sd_pvld;

output [8*64 -1:0] wt5_actv_data;
output [64 -1:0] wt5_actv_nz;
output [64 -1:0] wt5_actv_pvld;
output [64 -1:0] wt5_sd_mask;
output wt5_sd_pvld;

output [8*64 -1:0] wt6_actv_data;
output [64 -1:0] wt6_actv_nz;
output [64 -1:0] wt6_actv_pvld;
output [64 -1:0] wt6_sd_mask;
output wt6_sd_pvld;

output [8*64 -1:0] wt7_actv_data;
output [64 -1:0] wt7_actv_nz;
output [64 -1:0] wt7_actv_pvld;
output [64 -1:0] wt7_sd_mask;
output wt7_sd_pvld;

output [8*64 -1:0] wt8_actv_data;
output [64 -1:0] wt8_actv_nz;
output [64 -1:0] wt8_actv_pvld;
output [64 -1:0] wt8_sd_mask;
output wt8_sd_pvld;

output [8*64 -1:0] wt9_actv_data;
output [64 -1:0] wt9_actv_nz;
output [64 -1:0] wt9_actv_pvld;
output [64 -1:0] wt9_sd_mask;
output wt9_sd_pvld;

output [8*64 -1:0] wt10_actv_data;
output [64 -1:0] wt10_actv_nz;
output [64 -1:0] wt10_actv_pvld;
output [64 -1:0] wt10_sd_mask;
output wt10_sd_pvld;

output [8*64 -1:0] wt11_actv_data;
output [64 -1:0] wt11_actv_nz;
output [64 -1:0] wt11_actv_pvld;
output [64 -1:0] wt11_sd_mask;
output wt11_sd_pvld;

output [8*64 -1:0] wt12_actv_data;
output [64 -1:0] wt12_actv_nz;
output [64 -1:0] wt12_actv_pvld;
output [64 -1:0] wt12_sd_mask;
output wt12_sd_pvld;

output [8*64 -1:0] wt13_actv_data;
output [64 -1:0] wt13_actv_nz;
output [64 -1:0] wt13_actv_pvld;
output [64 -1:0] wt13_sd_mask;
output wt13_sd_pvld;

output [8*64 -1:0] wt14_actv_data;
output [64 -1:0] wt14_actv_nz;
output [64 -1:0] wt14_actv_pvld;
output [64 -1:0] wt14_sd_mask;
output wt14_sd_pvld;

output [8*64 -1:0] wt15_actv_data;
output [64 -1:0] wt15_actv_nz;
output [64 -1:0] wt15_actv_pvld;
output [64 -1:0] wt15_sd_mask;
output wt15_sd_pvld;

NV_NVDLA_CMAC_CORE_active_gate sodla_active(
    .io_nvdla_core_clk(nvdla_core_clk),
    .io_nvdla_core_rstn(nvdla_core_rstn),
    .io_in_dat_valid(in_dat_pvld),
    .io_in_dat_bits_mask_0(in_dat_mask[0]),
    .io_in_dat_bits_mask_1(in_dat_mask[1]),
    .io_in_dat_bits_mask_2(in_dat_mask[2]),
    .io_in_dat_bits_mask_3(in_dat_mask[3]),
    .io_in_dat_bits_mask_4(in_dat_mask[4]),
    .io_in_dat_bits_mask_5(in_dat_mask[5]),
    .io_in_dat_bits_mask_6(in_dat_mask[6]),
    .io_in_dat_bits_mask_7(in_dat_mask[7]),
    .io_in_dat_bits_mask_8(in_dat_mask[8]),
    .io_in_dat_bits_mask_9(in_dat_mask[9]),
    .io_in_dat_bits_mask_10(in_dat_mask[10]),
    .io_in_dat_bits_mask_11(in_dat_mask[11]),
    .io_in_dat_bits_mask_12(in_dat_mask[12]),
    .io_in_dat_bits_mask_13(in_dat_mask[13]),
    .io_in_dat_bits_mask_14(in_dat_mask[14]),
    .io_in_dat_bits_mask_15(in_dat_mask[15]),
    .io_in_dat_bits_mask_16(in_dat_mask[16]),
    .io_in_dat_bits_mask_17(in_dat_mask[17]),
    .io_in_dat_bits_mask_18(in_dat_mask[18]),
    .io_in_dat_bits_mask_19(in_dat_mask[19]),
    .io_in_dat_bits_mask_20(in_dat_mask[20]),
    .io_in_dat_bits_mask_21(in_dat_mask[21]),
    .io_in_dat_bits_mask_22(in_dat_mask[22]),
    .io_in_dat_bits_mask_23(in_dat_mask[23]),
    .io_in_dat_bits_mask_24(in_dat_mask[24]),
    .io_in_dat_bits_mask_25(in_dat_mask[25]),
    .io_in_dat_bits_mask_26(in_dat_mask[26]),
    .io_in_dat_bits_mask_27(in_dat_mask[27]),
    .io_in_dat_bits_mask_28(in_dat_mask[28]),
    .io_in_dat_bits_mask_29(in_dat_mask[29]),
    .io_in_dat_bits_mask_30(in_dat_mask[30]),
    .io_in_dat_bits_mask_31(in_dat_mask[31]),
    .io_in_dat_bits_mask_32(in_dat_mask[32]),
    .io_in_dat_bits_mask_33(in_dat_mask[33]),
    .io_in_dat_bits_mask_34(in_dat_mask[34]),
    .io_in_dat_bits_mask_35(in_dat_mask[35]),
    .io_in_dat_bits_mask_36(in_dat_mask[36]),
    .io_in_dat_bits_mask_37(in_dat_mask[37]),
    .io_in_dat_bits_mask_38(in_dat_mask[38]),
    .io_in_dat_bits_mask_39(in_dat_mask[39]),
    .io_in_dat_bits_mask_40(in_dat_mask[40]),
    .io_in_dat_bits_mask_41(in_dat_mask[41]),
    .io_in_dat_bits_mask_42(in_dat_mask[42]),
    .io_in_dat_bits_mask_43(in_dat_mask[43]),
    .io_in_dat_bits_mask_44(in_dat_mask[44]),
    .io_in_dat_bits_mask_45(in_dat_mask[45]),
    .io_in_dat_bits_mask_46(in_dat_mask[46]),
    .io_in_dat_bits_mask_47(in_dat_mask[47]),
    .io_in_dat_bits_mask_48(in_dat_mask[48]),
    .io_in_dat_bits_mask_49(in_dat_mask[49]),
    .io_in_dat_bits_mask_50(in_dat_mask[50]),
    .io_in_dat_bits_mask_51(in_dat_mask[51]),
    .io_in_dat_bits_mask_52(in_dat_mask[52]),
    .io_in_dat_bits_mask_53(in_dat_mask[53]),
    .io_in_dat_bits_mask_54(in_dat_mask[54]),
    .io_in_dat_bits_mask_55(in_dat_mask[55]),
    .io_in_dat_bits_mask_56(in_dat_mask[56]),
    .io_in_dat_bits_mask_57(in_dat_mask[57]),
    .io_in_dat_bits_mask_58(in_dat_mask[58]),
    .io_in_dat_bits_mask_59(in_dat_mask[59]),
    .io_in_dat_bits_mask_60(in_dat_mask[60]),
    .io_in_dat_bits_mask_61(in_dat_mask[61]),
    .io_in_dat_bits_mask_62(in_dat_mask[62]),
    .io_in_dat_bits_mask_63(in_dat_mask[63]),
    .io_in_dat_bits_data_0(in_dat_data0),
    .io_in_dat_bits_data_1(in_dat_data1),
    .io_in_dat_bits_data_2(in_dat_data2),
    .io_in_dat_bits_data_3(in_dat_data3),
    .io_in_dat_bits_data_4(in_dat_data4),
    .io_in_dat_bits_data_5(in_dat_data5),
    .io_in_dat_bits_data_6(in_dat_data6),
    .io_in_dat_bits_data_7(in_dat_data7),
    .io_in_dat_bits_data_8(in_dat_data8),
    .io_in_dat_bits_data_9(in_dat_data9),
    .io_in_dat_bits_data_10(in_dat_data10),
    .io_in_dat_bits_data_11(in_dat_data11),
    .io_in_dat_bits_data_12(in_dat_data12),
    .io_in_dat_bits_data_13(in_dat_data13),
    .io_in_dat_bits_data_14(in_dat_data14),
    .io_in_dat_bits_data_15(in_dat_data15),
    .io_in_dat_bits_data_16(in_dat_data16),
    .io_in_dat_bits_data_17(in_dat_data17),
    .io_in_dat_bits_data_18(in_dat_data18),
    .io_in_dat_bits_data_19(in_dat_data19),
    .io_in_dat_bits_data_20(in_dat_data20),
    .io_in_dat_bits_data_21(in_dat_data21),
    .io_in_dat_bits_data_22(in_dat_data22),
    .io_in_dat_bits_data_23(in_dat_data23),
    .io_in_dat_bits_data_24(in_dat_data24),
    .io_in_dat_bits_data_25(in_dat_data25),
    .io_in_dat_bits_data_26(in_dat_data26),
    .io_in_dat_bits_data_27(in_dat_data27),
    .io_in_dat_bits_data_28(in_dat_data28),
    .io_in_dat_bits_data_29(in_dat_data29),
    .io_in_dat_bits_data_30(in_dat_data30),
    .io_in_dat_bits_data_31(in_dat_data31),
    .io_in_dat_bits_data_32(in_dat_data32),
    .io_in_dat_bits_data_33(in_dat_data33),
    .io_in_dat_bits_data_34(in_dat_data34),
    .io_in_dat_bits_data_35(in_dat_data35),
    .io_in_dat_bits_data_36(in_dat_data36),
    .io_in_dat_bits_data_37(in_dat_data37),
    .io_in_dat_bits_data_38(in_dat_data38),
    .io_in_dat_bits_data_39(in_dat_data39),
    .io_in_dat_bits_data_40(in_dat_data40),
    .io_in_dat_bits_data_41(in_dat_data41),
    .io_in_dat_bits_data_42(in_dat_data42),
    .io_in_dat_bits_data_43(in_dat_data43),
    .io_in_dat_bits_data_44(in_dat_data44),
    .io_in_dat_bits_data_45(in_dat_data45),
    .io_in_dat_bits_data_46(in_dat_data46),
    .io_in_dat_bits_data_47(in_dat_data47),
    .io_in_dat_bits_data_48(in_dat_data48),
    .io_in_dat_bits_data_49(in_dat_data49),
    .io_in_dat_bits_data_50(in_dat_data50),
    .io_in_dat_bits_data_51(in_dat_data51),
    .io_in_dat_bits_data_52(in_dat_data52),
    .io_in_dat_bits_data_53(in_dat_data53),
    .io_in_dat_bits_data_54(in_dat_data54),
    .io_in_dat_bits_data_55(in_dat_data55),
    .io_in_dat_bits_data_56(in_dat_data56),
    .io_in_dat_bits_data_57(in_dat_data57),
    .io_in_dat_bits_data_58(in_dat_data58),
    .io_in_dat_bits_data_59(in_dat_data59),
    .io_in_dat_bits_data_60(in_dat_data60),
    .io_in_dat_bits_data_61(in_dat_data61),
    .io_in_dat_bits_data_62(in_dat_data62),
    .io_in_dat_bits_data_63(in_dat_data63),
//    .io_in_dat_bits_pd(xxx),
    .io_in_dat_stripe_st(in_dat_stripe_st),
    .io_in_dat_stripe_end(in_dat_stripe_end),
    .io_in_wt_valid(in_wt_pvld),
    .io_in_wt_bits_sel_0(in_wt_sel[0]),
    .io_in_wt_bits_sel_1(in_wt_sel[1]),
    .io_in_wt_bits_sel_2(in_wt_sel[2]),
    .io_in_wt_bits_sel_3(in_wt_sel[3]),
    .io_in_wt_bits_sel_4(in_wt_sel[4]),
    .io_in_wt_bits_sel_5(in_wt_sel[5]),
    .io_in_wt_bits_sel_6(in_wt_sel[6]),
    .io_in_wt_bits_sel_7(in_wt_sel[7]),
    .io_in_wt_bits_sel_8(in_wt_sel[8]),
    .io_in_wt_bits_sel_9(in_wt_sel[9]),
    .io_in_wt_bits_sel_10(in_wt_sel[10]),
    .io_in_wt_bits_sel_11(in_wt_sel[11]),
    .io_in_wt_bits_sel_12(in_wt_sel[12]),
    .io_in_wt_bits_sel_13(in_wt_sel[13]),
    .io_in_wt_bits_sel_14(in_wt_sel[14]),
    .io_in_wt_bits_sel_15(in_wt_sel[15]),
    .io_in_wt_bits_mask_0(in_wt_mask[0]),
    .io_in_wt_bits_mask_1(in_wt_mask[1]),
    .io_in_wt_bits_mask_2(in_wt_mask[2]),
    .io_in_wt_bits_mask_3(in_wt_mask[3]),
    .io_in_wt_bits_mask_4(in_wt_mask[4]),
    .io_in_wt_bits_mask_5(in_wt_mask[5]),
    .io_in_wt_bits_mask_6(in_wt_mask[6]),
    .io_in_wt_bits_mask_7(in_wt_mask[7]),
    .io_in_wt_bits_mask_8(in_wt_mask[8]),
    .io_in_wt_bits_mask_9(in_wt_mask[9]),
    .io_in_wt_bits_mask_10(in_wt_mask[10]),
    .io_in_wt_bits_mask_11(in_wt_mask[11]),
    .io_in_wt_bits_mask_12(in_wt_mask[12]),
    .io_in_wt_bits_mask_13(in_wt_mask[13]),
    .io_in_wt_bits_mask_14(in_wt_mask[14]),
    .io_in_wt_bits_mask_15(in_wt_mask[15]),
    .io_in_wt_bits_mask_16(in_wt_mask[16]),
    .io_in_wt_bits_mask_17(in_wt_mask[17]),
    .io_in_wt_bits_mask_18(in_wt_mask[18]),
    .io_in_wt_bits_mask_19(in_wt_mask[19]),
    .io_in_wt_bits_mask_20(in_wt_mask[20]),
    .io_in_wt_bits_mask_21(in_wt_mask[21]),
    .io_in_wt_bits_mask_22(in_wt_mask[22]),
    .io_in_wt_bits_mask_23(in_wt_mask[23]),
    .io_in_wt_bits_mask_24(in_wt_mask[24]),
    .io_in_wt_bits_mask_25(in_wt_mask[25]),
    .io_in_wt_bits_mask_26(in_wt_mask[26]),
    .io_in_wt_bits_mask_27(in_wt_mask[27]),
    .io_in_wt_bits_mask_28(in_wt_mask[28]),
    .io_in_wt_bits_mask_29(in_wt_mask[29]),
    .io_in_wt_bits_mask_30(in_wt_mask[30]),
    .io_in_wt_bits_mask_31(in_wt_mask[31]),
    .io_in_wt_bits_mask_32(in_wt_mask[32]),
    .io_in_wt_bits_mask_33(in_wt_mask[33]),
    .io_in_wt_bits_mask_34(in_wt_mask[34]),
    .io_in_wt_bits_mask_35(in_wt_mask[35]),
    .io_in_wt_bits_mask_36(in_wt_mask[36]),
    .io_in_wt_bits_mask_37(in_wt_mask[37]),
    .io_in_wt_bits_mask_38(in_wt_mask[38]),
    .io_in_wt_bits_mask_39(in_wt_mask[39]),
    .io_in_wt_bits_mask_40(in_wt_mask[40]),
    .io_in_wt_bits_mask_41(in_wt_mask[41]),
    .io_in_wt_bits_mask_42(in_wt_mask[42]),
    .io_in_wt_bits_mask_43(in_wt_mask[43]),
    .io_in_wt_bits_mask_44(in_wt_mask[44]),
    .io_in_wt_bits_mask_45(in_wt_mask[45]),
    .io_in_wt_bits_mask_46(in_wt_mask[46]),
    .io_in_wt_bits_mask_47(in_wt_mask[47]),
    .io_in_wt_bits_mask_48(in_wt_mask[48]),
    .io_in_wt_bits_mask_49(in_wt_mask[49]),
    .io_in_wt_bits_mask_50(in_wt_mask[50]),
    .io_in_wt_bits_mask_51(in_wt_mask[51]),
    .io_in_wt_bits_mask_52(in_wt_mask[52]),
    .io_in_wt_bits_mask_53(in_wt_mask[53]),
    .io_in_wt_bits_mask_54(in_wt_mask[54]),
    .io_in_wt_bits_mask_55(in_wt_mask[55]),
    .io_in_wt_bits_mask_56(in_wt_mask[56]),
    .io_in_wt_bits_mask_57(in_wt_mask[57]),
    .io_in_wt_bits_mask_58(in_wt_mask[58]),
    .io_in_wt_bits_mask_59(in_wt_mask[59]),
    .io_in_wt_bits_mask_60(in_wt_mask[60]),
    .io_in_wt_bits_mask_61(in_wt_mask[61]),
    .io_in_wt_bits_mask_62(in_wt_mask[62]),
    .io_in_wt_bits_mask_63(in_wt_mask[63]),
    .io_in_wt_bits_data_0(in_wt_data0),
    .io_in_wt_bits_data_1(in_wt_data1),
    .io_in_wt_bits_data_2(in_wt_data2),
    .io_in_wt_bits_data_3(in_wt_data3),
    .io_in_wt_bits_data_4(in_wt_data4),
    .io_in_wt_bits_data_5(in_wt_data5),
    .io_in_wt_bits_data_6(in_wt_data6),
    .io_in_wt_bits_data_7(in_wt_data7),
    .io_in_wt_bits_data_8(in_wt_data8),
    .io_in_wt_bits_data_9(in_wt_data9),
    .io_in_wt_bits_data_10(in_wt_data10),
    .io_in_wt_bits_data_11(in_wt_data11),
    .io_in_wt_bits_data_12(in_wt_data12),
    .io_in_wt_bits_data_13(in_wt_data13),
    .io_in_wt_bits_data_14(in_wt_data14),
    .io_in_wt_bits_data_15(in_wt_data15),
    .io_in_wt_bits_data_16(in_wt_data16),
    .io_in_wt_bits_data_17(in_wt_data17),
    .io_in_wt_bits_data_18(in_wt_data18),
    .io_in_wt_bits_data_19(in_wt_data19),
    .io_in_wt_bits_data_20(in_wt_data20),
    .io_in_wt_bits_data_21(in_wt_data21),
    .io_in_wt_bits_data_22(in_wt_data22),
    .io_in_wt_bits_data_23(in_wt_data23),
    .io_in_wt_bits_data_24(in_wt_data24),
    .io_in_wt_bits_data_25(in_wt_data25),
    .io_in_wt_bits_data_26(in_wt_data26),
    .io_in_wt_bits_data_27(in_wt_data27),
    .io_in_wt_bits_data_28(in_wt_data28),
    .io_in_wt_bits_data_29(in_wt_data29),
    .io_in_wt_bits_data_30(in_wt_data30),
    .io_in_wt_bits_data_31(in_wt_data31),
    .io_in_wt_bits_data_32(in_wt_data32),
    .io_in_wt_bits_data_33(in_wt_data33),
    .io_in_wt_bits_data_34(in_wt_data34),
    .io_in_wt_bits_data_35(in_wt_data35),
    .io_in_wt_bits_data_36(in_wt_data36),
    .io_in_wt_bits_data_37(in_wt_data37),
    .io_in_wt_bits_data_38(in_wt_data38),
    .io_in_wt_bits_data_39(in_wt_data39),
    .io_in_wt_bits_data_40(in_wt_data40),
    .io_in_wt_bits_data_41(in_wt_data41),
    .io_in_wt_bits_data_42(in_wt_data42),
    .io_in_wt_bits_data_43(in_wt_data43),
    .io_in_wt_bits_data_44(in_wt_data44),
    .io_in_wt_bits_data_45(in_wt_data45),
    .io_in_wt_bits_data_46(in_wt_data46),
    .io_in_wt_bits_data_47(in_wt_data47),
    .io_in_wt_bits_data_48(in_wt_data48),
    .io_in_wt_bits_data_49(in_wt_data49),
    .io_in_wt_bits_data_50(in_wt_data50),
    .io_in_wt_bits_data_51(in_wt_data51),
    .io_in_wt_bits_data_52(in_wt_data52),
    .io_in_wt_bits_data_53(in_wt_data53),
    .io_in_wt_bits_data_54(in_wt_data54),
    .io_in_wt_bits_data_55(in_wt_data55),
    .io_in_wt_bits_data_56(in_wt_data56),
    .io_in_wt_bits_data_57(in_wt_data57),
    .io_in_wt_bits_data_58(in_wt_data58),
    .io_in_wt_bits_data_59(in_wt_data59),
    .io_in_wt_bits_data_60(in_wt_data60),
    .io_in_wt_bits_data_61(in_wt_data61),
    .io_in_wt_bits_data_62(in_wt_data62),
    .io_in_wt_bits_data_63(in_wt_data63),
    .io_dat_actv_0_0_valid(dat0_actv_pvld[0]),
.io_dat_actv_0_0_bits_nz(dat0_actv_nz[0]),
.io_dat_actv_0_0_bits_data(dat0_actv_data[7:0]),

.io_dat_actv_0_1_valid(dat0_actv_pvld[1]),
.io_dat_actv_0_1_bits_nz(dat0_actv_nz[1]),
.io_dat_actv_0_1_bits_data(dat0_actv_data[15:8]),

.io_dat_actv_0_2_valid(dat0_actv_pvld[2]),
.io_dat_actv_0_2_bits_nz(dat0_actv_nz[2]),
.io_dat_actv_0_2_bits_data(dat0_actv_data[23:16]),

.io_dat_actv_0_3_valid(dat0_actv_pvld[3]),
.io_dat_actv_0_3_bits_nz(dat0_actv_nz[3]),
.io_dat_actv_0_3_bits_data(dat0_actv_data[31:24]),

.io_dat_actv_0_4_valid(dat0_actv_pvld[4]),
.io_dat_actv_0_4_bits_nz(dat0_actv_nz[4]),
.io_dat_actv_0_4_bits_data(dat0_actv_data[39:32]),

.io_dat_actv_0_5_valid(dat0_actv_pvld[5]),
.io_dat_actv_0_5_bits_nz(dat0_actv_nz[5]),
.io_dat_actv_0_5_bits_data(dat0_actv_data[47:40]),

.io_dat_actv_0_6_valid(dat0_actv_pvld[6]),
.io_dat_actv_0_6_bits_nz(dat0_actv_nz[6]),
.io_dat_actv_0_6_bits_data(dat0_actv_data[55:48]),

.io_dat_actv_0_7_valid(dat0_actv_pvld[7]),
.io_dat_actv_0_7_bits_nz(dat0_actv_nz[7]),
.io_dat_actv_0_7_bits_data(dat0_actv_data[63:56]),

.io_dat_actv_0_8_valid(dat0_actv_pvld[8]),
.io_dat_actv_0_8_bits_nz(dat0_actv_nz[8]),
.io_dat_actv_0_8_bits_data(dat0_actv_data[71:64]),

.io_dat_actv_0_9_valid(dat0_actv_pvld[9]),
.io_dat_actv_0_9_bits_nz(dat0_actv_nz[9]),
.io_dat_actv_0_9_bits_data(dat0_actv_data[79:72]),

.io_dat_actv_0_10_valid(dat0_actv_pvld[10]),
.io_dat_actv_0_10_bits_nz(dat0_actv_nz[10]),
.io_dat_actv_0_10_bits_data(dat0_actv_data[87:80]),

.io_dat_actv_0_11_valid(dat0_actv_pvld[11]),
.io_dat_actv_0_11_bits_nz(dat0_actv_nz[11]),
.io_dat_actv_0_11_bits_data(dat0_actv_data[95:88]),

.io_dat_actv_0_12_valid(dat0_actv_pvld[12]),
.io_dat_actv_0_12_bits_nz(dat0_actv_nz[12]),
.io_dat_actv_0_12_bits_data(dat0_actv_data[103:96]),

.io_dat_actv_0_13_valid(dat0_actv_pvld[13]),
.io_dat_actv_0_13_bits_nz(dat0_actv_nz[13]),
.io_dat_actv_0_13_bits_data(dat0_actv_data[111:104]),

.io_dat_actv_0_14_valid(dat0_actv_pvld[14]),
.io_dat_actv_0_14_bits_nz(dat0_actv_nz[14]),
.io_dat_actv_0_14_bits_data(dat0_actv_data[119:112]),

.io_dat_actv_0_15_valid(dat0_actv_pvld[15]),
.io_dat_actv_0_15_bits_nz(dat0_actv_nz[15]),
.io_dat_actv_0_15_bits_data(dat0_actv_data[127:120]),

.io_dat_actv_0_16_valid(dat0_actv_pvld[16]),
.io_dat_actv_0_16_bits_nz(dat0_actv_nz[16]),
.io_dat_actv_0_16_bits_data(dat0_actv_data[135:128]),

.io_dat_actv_0_17_valid(dat0_actv_pvld[17]),
.io_dat_actv_0_17_bits_nz(dat0_actv_nz[17]),
.io_dat_actv_0_17_bits_data(dat0_actv_data[143:136]),

.io_dat_actv_0_18_valid(dat0_actv_pvld[18]),
.io_dat_actv_0_18_bits_nz(dat0_actv_nz[18]),
.io_dat_actv_0_18_bits_data(dat0_actv_data[151:144]),

.io_dat_actv_0_19_valid(dat0_actv_pvld[19]),
.io_dat_actv_0_19_bits_nz(dat0_actv_nz[19]),
.io_dat_actv_0_19_bits_data(dat0_actv_data[159:152]),

.io_dat_actv_0_20_valid(dat0_actv_pvld[20]),
.io_dat_actv_0_20_bits_nz(dat0_actv_nz[20]),
.io_dat_actv_0_20_bits_data(dat0_actv_data[167:160]),

.io_dat_actv_0_21_valid(dat0_actv_pvld[21]),
.io_dat_actv_0_21_bits_nz(dat0_actv_nz[21]),
.io_dat_actv_0_21_bits_data(dat0_actv_data[175:168]),

.io_dat_actv_0_22_valid(dat0_actv_pvld[22]),
.io_dat_actv_0_22_bits_nz(dat0_actv_nz[22]),
.io_dat_actv_0_22_bits_data(dat0_actv_data[183:176]),

.io_dat_actv_0_23_valid(dat0_actv_pvld[23]),
.io_dat_actv_0_23_bits_nz(dat0_actv_nz[23]),
.io_dat_actv_0_23_bits_data(dat0_actv_data[191:184]),

.io_dat_actv_0_24_valid(dat0_actv_pvld[24]),
.io_dat_actv_0_24_bits_nz(dat0_actv_nz[24]),
.io_dat_actv_0_24_bits_data(dat0_actv_data[199:192]),

.io_dat_actv_0_25_valid(dat0_actv_pvld[25]),
.io_dat_actv_0_25_bits_nz(dat0_actv_nz[25]),
.io_dat_actv_0_25_bits_data(dat0_actv_data[207:200]),

.io_dat_actv_0_26_valid(dat0_actv_pvld[26]),
.io_dat_actv_0_26_bits_nz(dat0_actv_nz[26]),
.io_dat_actv_0_26_bits_data(dat0_actv_data[215:208]),

.io_dat_actv_0_27_valid(dat0_actv_pvld[27]),
.io_dat_actv_0_27_bits_nz(dat0_actv_nz[27]),
.io_dat_actv_0_27_bits_data(dat0_actv_data[223:216]),

.io_dat_actv_0_28_valid(dat0_actv_pvld[28]),
.io_dat_actv_0_28_bits_nz(dat0_actv_nz[28]),
.io_dat_actv_0_28_bits_data(dat0_actv_data[231:224]),

.io_dat_actv_0_29_valid(dat0_actv_pvld[29]),
.io_dat_actv_0_29_bits_nz(dat0_actv_nz[29]),
.io_dat_actv_0_29_bits_data(dat0_actv_data[239:232]),

.io_dat_actv_0_30_valid(dat0_actv_pvld[30]),
.io_dat_actv_0_30_bits_nz(dat0_actv_nz[30]),
.io_dat_actv_0_30_bits_data(dat0_actv_data[247:240]),

.io_dat_actv_0_31_valid(dat0_actv_pvld[31]),
.io_dat_actv_0_31_bits_nz(dat0_actv_nz[31]),
.io_dat_actv_0_31_bits_data(dat0_actv_data[255:248]),

.io_dat_actv_0_32_valid(dat0_actv_pvld[32]),
.io_dat_actv_0_32_bits_nz(dat0_actv_nz[32]),
.io_dat_actv_0_32_bits_data(dat0_actv_data[263:256]),

.io_dat_actv_0_33_valid(dat0_actv_pvld[33]),
.io_dat_actv_0_33_bits_nz(dat0_actv_nz[33]),
.io_dat_actv_0_33_bits_data(dat0_actv_data[271:264]),

.io_dat_actv_0_34_valid(dat0_actv_pvld[34]),
.io_dat_actv_0_34_bits_nz(dat0_actv_nz[34]),
.io_dat_actv_0_34_bits_data(dat0_actv_data[279:272]),

.io_dat_actv_0_35_valid(dat0_actv_pvld[35]),
.io_dat_actv_0_35_bits_nz(dat0_actv_nz[35]),
.io_dat_actv_0_35_bits_data(dat0_actv_data[287:280]),

.io_dat_actv_0_36_valid(dat0_actv_pvld[36]),
.io_dat_actv_0_36_bits_nz(dat0_actv_nz[36]),
.io_dat_actv_0_36_bits_data(dat0_actv_data[295:288]),

.io_dat_actv_0_37_valid(dat0_actv_pvld[37]),
.io_dat_actv_0_37_bits_nz(dat0_actv_nz[37]),
.io_dat_actv_0_37_bits_data(dat0_actv_data[303:296]),

.io_dat_actv_0_38_valid(dat0_actv_pvld[38]),
.io_dat_actv_0_38_bits_nz(dat0_actv_nz[38]),
.io_dat_actv_0_38_bits_data(dat0_actv_data[311:304]),

.io_dat_actv_0_39_valid(dat0_actv_pvld[39]),
.io_dat_actv_0_39_bits_nz(dat0_actv_nz[39]),
.io_dat_actv_0_39_bits_data(dat0_actv_data[319:312]),

.io_dat_actv_0_40_valid(dat0_actv_pvld[40]),
.io_dat_actv_0_40_bits_nz(dat0_actv_nz[40]),
.io_dat_actv_0_40_bits_data(dat0_actv_data[327:320]),

.io_dat_actv_0_41_valid(dat0_actv_pvld[41]),
.io_dat_actv_0_41_bits_nz(dat0_actv_nz[41]),
.io_dat_actv_0_41_bits_data(dat0_actv_data[335:328]),

.io_dat_actv_0_42_valid(dat0_actv_pvld[42]),
.io_dat_actv_0_42_bits_nz(dat0_actv_nz[42]),
.io_dat_actv_0_42_bits_data(dat0_actv_data[343:336]),

.io_dat_actv_0_43_valid(dat0_actv_pvld[43]),
.io_dat_actv_0_43_bits_nz(dat0_actv_nz[43]),
.io_dat_actv_0_43_bits_data(dat0_actv_data[351:344]),

.io_dat_actv_0_44_valid(dat0_actv_pvld[44]),
.io_dat_actv_0_44_bits_nz(dat0_actv_nz[44]),
.io_dat_actv_0_44_bits_data(dat0_actv_data[359:352]),

.io_dat_actv_0_45_valid(dat0_actv_pvld[45]),
.io_dat_actv_0_45_bits_nz(dat0_actv_nz[45]),
.io_dat_actv_0_45_bits_data(dat0_actv_data[367:360]),

.io_dat_actv_0_46_valid(dat0_actv_pvld[46]),
.io_dat_actv_0_46_bits_nz(dat0_actv_nz[46]),
.io_dat_actv_0_46_bits_data(dat0_actv_data[375:368]),

.io_dat_actv_0_47_valid(dat0_actv_pvld[47]),
.io_dat_actv_0_47_bits_nz(dat0_actv_nz[47]),
.io_dat_actv_0_47_bits_data(dat0_actv_data[383:376]),

.io_dat_actv_0_48_valid(dat0_actv_pvld[48]),
.io_dat_actv_0_48_bits_nz(dat0_actv_nz[48]),
.io_dat_actv_0_48_bits_data(dat0_actv_data[391:384]),

.io_dat_actv_0_49_valid(dat0_actv_pvld[49]),
.io_dat_actv_0_49_bits_nz(dat0_actv_nz[49]),
.io_dat_actv_0_49_bits_data(dat0_actv_data[399:392]),

.io_dat_actv_0_50_valid(dat0_actv_pvld[50]),
.io_dat_actv_0_50_bits_nz(dat0_actv_nz[50]),
.io_dat_actv_0_50_bits_data(dat0_actv_data[407:400]),

.io_dat_actv_0_51_valid(dat0_actv_pvld[51]),
.io_dat_actv_0_51_bits_nz(dat0_actv_nz[51]),
.io_dat_actv_0_51_bits_data(dat0_actv_data[415:408]),

.io_dat_actv_0_52_valid(dat0_actv_pvld[52]),
.io_dat_actv_0_52_bits_nz(dat0_actv_nz[52]),
.io_dat_actv_0_52_bits_data(dat0_actv_data[423:416]),

.io_dat_actv_0_53_valid(dat0_actv_pvld[53]),
.io_dat_actv_0_53_bits_nz(dat0_actv_nz[53]),
.io_dat_actv_0_53_bits_data(dat0_actv_data[431:424]),

.io_dat_actv_0_54_valid(dat0_actv_pvld[54]),
.io_dat_actv_0_54_bits_nz(dat0_actv_nz[54]),
.io_dat_actv_0_54_bits_data(dat0_actv_data[439:432]),

.io_dat_actv_0_55_valid(dat0_actv_pvld[55]),
.io_dat_actv_0_55_bits_nz(dat0_actv_nz[55]),
.io_dat_actv_0_55_bits_data(dat0_actv_data[447:440]),

.io_dat_actv_0_56_valid(dat0_actv_pvld[56]),
.io_dat_actv_0_56_bits_nz(dat0_actv_nz[56]),
.io_dat_actv_0_56_bits_data(dat0_actv_data[455:448]),

.io_dat_actv_0_57_valid(dat0_actv_pvld[57]),
.io_dat_actv_0_57_bits_nz(dat0_actv_nz[57]),
.io_dat_actv_0_57_bits_data(dat0_actv_data[463:456]),

.io_dat_actv_0_58_valid(dat0_actv_pvld[58]),
.io_dat_actv_0_58_bits_nz(dat0_actv_nz[58]),
.io_dat_actv_0_58_bits_data(dat0_actv_data[471:464]),

.io_dat_actv_0_59_valid(dat0_actv_pvld[59]),
.io_dat_actv_0_59_bits_nz(dat0_actv_nz[59]),
.io_dat_actv_0_59_bits_data(dat0_actv_data[479:472]),

.io_dat_actv_0_60_valid(dat0_actv_pvld[60]),
.io_dat_actv_0_60_bits_nz(dat0_actv_nz[60]),
.io_dat_actv_0_60_bits_data(dat0_actv_data[487:480]),

.io_dat_actv_0_61_valid(dat0_actv_pvld[61]),
.io_dat_actv_0_61_bits_nz(dat0_actv_nz[61]),
.io_dat_actv_0_61_bits_data(dat0_actv_data[495:488]),

.io_dat_actv_0_62_valid(dat0_actv_pvld[62]),
.io_dat_actv_0_62_bits_nz(dat0_actv_nz[62]),
.io_dat_actv_0_62_bits_data(dat0_actv_data[503:496]),

.io_dat_actv_0_63_valid(dat0_actv_pvld[63]),
.io_dat_actv_0_63_bits_nz(dat0_actv_nz[63]),
.io_dat_actv_0_63_bits_data(dat0_actv_data[511:504]),

.io_dat_actv_1_0_valid(dat1_actv_pvld[0]),
.io_dat_actv_1_0_bits_nz(dat1_actv_nz[0]),
.io_dat_actv_1_0_bits_data(dat1_actv_data[7:0]),

.io_dat_actv_1_1_valid(dat1_actv_pvld[1]),
.io_dat_actv_1_1_bits_nz(dat1_actv_nz[1]),
.io_dat_actv_1_1_bits_data(dat1_actv_data[15:8]),

.io_dat_actv_1_2_valid(dat1_actv_pvld[2]),
.io_dat_actv_1_2_bits_nz(dat1_actv_nz[2]),
.io_dat_actv_1_2_bits_data(dat1_actv_data[23:16]),

.io_dat_actv_1_3_valid(dat1_actv_pvld[3]),
.io_dat_actv_1_3_bits_nz(dat1_actv_nz[3]),
.io_dat_actv_1_3_bits_data(dat1_actv_data[31:24]),

.io_dat_actv_1_4_valid(dat1_actv_pvld[4]),
.io_dat_actv_1_4_bits_nz(dat1_actv_nz[4]),
.io_dat_actv_1_4_bits_data(dat1_actv_data[39:32]),

.io_dat_actv_1_5_valid(dat1_actv_pvld[5]),
.io_dat_actv_1_5_bits_nz(dat1_actv_nz[5]),
.io_dat_actv_1_5_bits_data(dat1_actv_data[47:40]),

.io_dat_actv_1_6_valid(dat1_actv_pvld[6]),
.io_dat_actv_1_6_bits_nz(dat1_actv_nz[6]),
.io_dat_actv_1_6_bits_data(dat1_actv_data[55:48]),

.io_dat_actv_1_7_valid(dat1_actv_pvld[7]),
.io_dat_actv_1_7_bits_nz(dat1_actv_nz[7]),
.io_dat_actv_1_7_bits_data(dat1_actv_data[63:56]),

.io_dat_actv_1_8_valid(dat1_actv_pvld[8]),
.io_dat_actv_1_8_bits_nz(dat1_actv_nz[8]),
.io_dat_actv_1_8_bits_data(dat1_actv_data[71:64]),

.io_dat_actv_1_9_valid(dat1_actv_pvld[9]),
.io_dat_actv_1_9_bits_nz(dat1_actv_nz[9]),
.io_dat_actv_1_9_bits_data(dat1_actv_data[79:72]),

.io_dat_actv_1_10_valid(dat1_actv_pvld[10]),
.io_dat_actv_1_10_bits_nz(dat1_actv_nz[10]),
.io_dat_actv_1_10_bits_data(dat1_actv_data[87:80]),

.io_dat_actv_1_11_valid(dat1_actv_pvld[11]),
.io_dat_actv_1_11_bits_nz(dat1_actv_nz[11]),
.io_dat_actv_1_11_bits_data(dat1_actv_data[95:88]),

.io_dat_actv_1_12_valid(dat1_actv_pvld[12]),
.io_dat_actv_1_12_bits_nz(dat1_actv_nz[12]),
.io_dat_actv_1_12_bits_data(dat1_actv_data[103:96]),

.io_dat_actv_1_13_valid(dat1_actv_pvld[13]),
.io_dat_actv_1_13_bits_nz(dat1_actv_nz[13]),
.io_dat_actv_1_13_bits_data(dat1_actv_data[111:104]),

.io_dat_actv_1_14_valid(dat1_actv_pvld[14]),
.io_dat_actv_1_14_bits_nz(dat1_actv_nz[14]),
.io_dat_actv_1_14_bits_data(dat1_actv_data[119:112]),

.io_dat_actv_1_15_valid(dat1_actv_pvld[15]),
.io_dat_actv_1_15_bits_nz(dat1_actv_nz[15]),
.io_dat_actv_1_15_bits_data(dat1_actv_data[127:120]),

.io_dat_actv_1_16_valid(dat1_actv_pvld[16]),
.io_dat_actv_1_16_bits_nz(dat1_actv_nz[16]),
.io_dat_actv_1_16_bits_data(dat1_actv_data[135:128]),

.io_dat_actv_1_17_valid(dat1_actv_pvld[17]),
.io_dat_actv_1_17_bits_nz(dat1_actv_nz[17]),
.io_dat_actv_1_17_bits_data(dat1_actv_data[143:136]),

.io_dat_actv_1_18_valid(dat1_actv_pvld[18]),
.io_dat_actv_1_18_bits_nz(dat1_actv_nz[18]),
.io_dat_actv_1_18_bits_data(dat1_actv_data[151:144]),

.io_dat_actv_1_19_valid(dat1_actv_pvld[19]),
.io_dat_actv_1_19_bits_nz(dat1_actv_nz[19]),
.io_dat_actv_1_19_bits_data(dat1_actv_data[159:152]),

.io_dat_actv_1_20_valid(dat1_actv_pvld[20]),
.io_dat_actv_1_20_bits_nz(dat1_actv_nz[20]),
.io_dat_actv_1_20_bits_data(dat1_actv_data[167:160]),

.io_dat_actv_1_21_valid(dat1_actv_pvld[21]),
.io_dat_actv_1_21_bits_nz(dat1_actv_nz[21]),
.io_dat_actv_1_21_bits_data(dat1_actv_data[175:168]),

.io_dat_actv_1_22_valid(dat1_actv_pvld[22]),
.io_dat_actv_1_22_bits_nz(dat1_actv_nz[22]),
.io_dat_actv_1_22_bits_data(dat1_actv_data[183:176]),

.io_dat_actv_1_23_valid(dat1_actv_pvld[23]),
.io_dat_actv_1_23_bits_nz(dat1_actv_nz[23]),
.io_dat_actv_1_23_bits_data(dat1_actv_data[191:184]),

.io_dat_actv_1_24_valid(dat1_actv_pvld[24]),
.io_dat_actv_1_24_bits_nz(dat1_actv_nz[24]),
.io_dat_actv_1_24_bits_data(dat1_actv_data[199:192]),

.io_dat_actv_1_25_valid(dat1_actv_pvld[25]),
.io_dat_actv_1_25_bits_nz(dat1_actv_nz[25]),
.io_dat_actv_1_25_bits_data(dat1_actv_data[207:200]),

.io_dat_actv_1_26_valid(dat1_actv_pvld[26]),
.io_dat_actv_1_26_bits_nz(dat1_actv_nz[26]),
.io_dat_actv_1_26_bits_data(dat1_actv_data[215:208]),

.io_dat_actv_1_27_valid(dat1_actv_pvld[27]),
.io_dat_actv_1_27_bits_nz(dat1_actv_nz[27]),
.io_dat_actv_1_27_bits_data(dat1_actv_data[223:216]),

.io_dat_actv_1_28_valid(dat1_actv_pvld[28]),
.io_dat_actv_1_28_bits_nz(dat1_actv_nz[28]),
.io_dat_actv_1_28_bits_data(dat1_actv_data[231:224]),

.io_dat_actv_1_29_valid(dat1_actv_pvld[29]),
.io_dat_actv_1_29_bits_nz(dat1_actv_nz[29]),
.io_dat_actv_1_29_bits_data(dat1_actv_data[239:232]),

.io_dat_actv_1_30_valid(dat1_actv_pvld[30]),
.io_dat_actv_1_30_bits_nz(dat1_actv_nz[30]),
.io_dat_actv_1_30_bits_data(dat1_actv_data[247:240]),

.io_dat_actv_1_31_valid(dat1_actv_pvld[31]),
.io_dat_actv_1_31_bits_nz(dat1_actv_nz[31]),
.io_dat_actv_1_31_bits_data(dat1_actv_data[255:248]),

.io_dat_actv_1_32_valid(dat1_actv_pvld[32]),
.io_dat_actv_1_32_bits_nz(dat1_actv_nz[32]),
.io_dat_actv_1_32_bits_data(dat1_actv_data[263:256]),

.io_dat_actv_1_33_valid(dat1_actv_pvld[33]),
.io_dat_actv_1_33_bits_nz(dat1_actv_nz[33]),
.io_dat_actv_1_33_bits_data(dat1_actv_data[271:264]),

.io_dat_actv_1_34_valid(dat1_actv_pvld[34]),
.io_dat_actv_1_34_bits_nz(dat1_actv_nz[34]),
.io_dat_actv_1_34_bits_data(dat1_actv_data[279:272]),

.io_dat_actv_1_35_valid(dat1_actv_pvld[35]),
.io_dat_actv_1_35_bits_nz(dat1_actv_nz[35]),
.io_dat_actv_1_35_bits_data(dat1_actv_data[287:280]),

.io_dat_actv_1_36_valid(dat1_actv_pvld[36]),
.io_dat_actv_1_36_bits_nz(dat1_actv_nz[36]),
.io_dat_actv_1_36_bits_data(dat1_actv_data[295:288]),

.io_dat_actv_1_37_valid(dat1_actv_pvld[37]),
.io_dat_actv_1_37_bits_nz(dat1_actv_nz[37]),
.io_dat_actv_1_37_bits_data(dat1_actv_data[303:296]),

.io_dat_actv_1_38_valid(dat1_actv_pvld[38]),
.io_dat_actv_1_38_bits_nz(dat1_actv_nz[38]),
.io_dat_actv_1_38_bits_data(dat1_actv_data[311:304]),

.io_dat_actv_1_39_valid(dat1_actv_pvld[39]),
.io_dat_actv_1_39_bits_nz(dat1_actv_nz[39]),
.io_dat_actv_1_39_bits_data(dat1_actv_data[319:312]),

.io_dat_actv_1_40_valid(dat1_actv_pvld[40]),
.io_dat_actv_1_40_bits_nz(dat1_actv_nz[40]),
.io_dat_actv_1_40_bits_data(dat1_actv_data[327:320]),

.io_dat_actv_1_41_valid(dat1_actv_pvld[41]),
.io_dat_actv_1_41_bits_nz(dat1_actv_nz[41]),
.io_dat_actv_1_41_bits_data(dat1_actv_data[335:328]),

.io_dat_actv_1_42_valid(dat1_actv_pvld[42]),
.io_dat_actv_1_42_bits_nz(dat1_actv_nz[42]),
.io_dat_actv_1_42_bits_data(dat1_actv_data[343:336]),

.io_dat_actv_1_43_valid(dat1_actv_pvld[43]),
.io_dat_actv_1_43_bits_nz(dat1_actv_nz[43]),
.io_dat_actv_1_43_bits_data(dat1_actv_data[351:344]),

.io_dat_actv_1_44_valid(dat1_actv_pvld[44]),
.io_dat_actv_1_44_bits_nz(dat1_actv_nz[44]),
.io_dat_actv_1_44_bits_data(dat1_actv_data[359:352]),

.io_dat_actv_1_45_valid(dat1_actv_pvld[45]),
.io_dat_actv_1_45_bits_nz(dat1_actv_nz[45]),
.io_dat_actv_1_45_bits_data(dat1_actv_data[367:360]),

.io_dat_actv_1_46_valid(dat1_actv_pvld[46]),
.io_dat_actv_1_46_bits_nz(dat1_actv_nz[46]),
.io_dat_actv_1_46_bits_data(dat1_actv_data[375:368]),

.io_dat_actv_1_47_valid(dat1_actv_pvld[47]),
.io_dat_actv_1_47_bits_nz(dat1_actv_nz[47]),
.io_dat_actv_1_47_bits_data(dat1_actv_data[383:376]),

.io_dat_actv_1_48_valid(dat1_actv_pvld[48]),
.io_dat_actv_1_48_bits_nz(dat1_actv_nz[48]),
.io_dat_actv_1_48_bits_data(dat1_actv_data[391:384]),

.io_dat_actv_1_49_valid(dat1_actv_pvld[49]),
.io_dat_actv_1_49_bits_nz(dat1_actv_nz[49]),
.io_dat_actv_1_49_bits_data(dat1_actv_data[399:392]),

.io_dat_actv_1_50_valid(dat1_actv_pvld[50]),
.io_dat_actv_1_50_bits_nz(dat1_actv_nz[50]),
.io_dat_actv_1_50_bits_data(dat1_actv_data[407:400]),

.io_dat_actv_1_51_valid(dat1_actv_pvld[51]),
.io_dat_actv_1_51_bits_nz(dat1_actv_nz[51]),
.io_dat_actv_1_51_bits_data(dat1_actv_data[415:408]),

.io_dat_actv_1_52_valid(dat1_actv_pvld[52]),
.io_dat_actv_1_52_bits_nz(dat1_actv_nz[52]),
.io_dat_actv_1_52_bits_data(dat1_actv_data[423:416]),

.io_dat_actv_1_53_valid(dat1_actv_pvld[53]),
.io_dat_actv_1_53_bits_nz(dat1_actv_nz[53]),
.io_dat_actv_1_53_bits_data(dat1_actv_data[431:424]),

.io_dat_actv_1_54_valid(dat1_actv_pvld[54]),
.io_dat_actv_1_54_bits_nz(dat1_actv_nz[54]),
.io_dat_actv_1_54_bits_data(dat1_actv_data[439:432]),

.io_dat_actv_1_55_valid(dat1_actv_pvld[55]),
.io_dat_actv_1_55_bits_nz(dat1_actv_nz[55]),
.io_dat_actv_1_55_bits_data(dat1_actv_data[447:440]),

.io_dat_actv_1_56_valid(dat1_actv_pvld[56]),
.io_dat_actv_1_56_bits_nz(dat1_actv_nz[56]),
.io_dat_actv_1_56_bits_data(dat1_actv_data[455:448]),

.io_dat_actv_1_57_valid(dat1_actv_pvld[57]),
.io_dat_actv_1_57_bits_nz(dat1_actv_nz[57]),
.io_dat_actv_1_57_bits_data(dat1_actv_data[463:456]),

.io_dat_actv_1_58_valid(dat1_actv_pvld[58]),
.io_dat_actv_1_58_bits_nz(dat1_actv_nz[58]),
.io_dat_actv_1_58_bits_data(dat1_actv_data[471:464]),

.io_dat_actv_1_59_valid(dat1_actv_pvld[59]),
.io_dat_actv_1_59_bits_nz(dat1_actv_nz[59]),
.io_dat_actv_1_59_bits_data(dat1_actv_data[479:472]),

.io_dat_actv_1_60_valid(dat1_actv_pvld[60]),
.io_dat_actv_1_60_bits_nz(dat1_actv_nz[60]),
.io_dat_actv_1_60_bits_data(dat1_actv_data[487:480]),

.io_dat_actv_1_61_valid(dat1_actv_pvld[61]),
.io_dat_actv_1_61_bits_nz(dat1_actv_nz[61]),
.io_dat_actv_1_61_bits_data(dat1_actv_data[495:488]),

.io_dat_actv_1_62_valid(dat1_actv_pvld[62]),
.io_dat_actv_1_62_bits_nz(dat1_actv_nz[62]),
.io_dat_actv_1_62_bits_data(dat1_actv_data[503:496]),

.io_dat_actv_1_63_valid(dat1_actv_pvld[63]),
.io_dat_actv_1_63_bits_nz(dat1_actv_nz[63]),
.io_dat_actv_1_63_bits_data(dat1_actv_data[511:504]),

.io_dat_actv_2_0_valid(dat2_actv_pvld[0]),
.io_dat_actv_2_0_bits_nz(dat2_actv_nz[0]),
.io_dat_actv_2_0_bits_data(dat2_actv_data[7:0]),

.io_dat_actv_2_1_valid(dat2_actv_pvld[1]),
.io_dat_actv_2_1_bits_nz(dat2_actv_nz[1]),
.io_dat_actv_2_1_bits_data(dat2_actv_data[15:8]),

.io_dat_actv_2_2_valid(dat2_actv_pvld[2]),
.io_dat_actv_2_2_bits_nz(dat2_actv_nz[2]),
.io_dat_actv_2_2_bits_data(dat2_actv_data[23:16]),

.io_dat_actv_2_3_valid(dat2_actv_pvld[3]),
.io_dat_actv_2_3_bits_nz(dat2_actv_nz[3]),
.io_dat_actv_2_3_bits_data(dat2_actv_data[31:24]),

.io_dat_actv_2_4_valid(dat2_actv_pvld[4]),
.io_dat_actv_2_4_bits_nz(dat2_actv_nz[4]),
.io_dat_actv_2_4_bits_data(dat2_actv_data[39:32]),

.io_dat_actv_2_5_valid(dat2_actv_pvld[5]),
.io_dat_actv_2_5_bits_nz(dat2_actv_nz[5]),
.io_dat_actv_2_5_bits_data(dat2_actv_data[47:40]),

.io_dat_actv_2_6_valid(dat2_actv_pvld[6]),
.io_dat_actv_2_6_bits_nz(dat2_actv_nz[6]),
.io_dat_actv_2_6_bits_data(dat2_actv_data[55:48]),

.io_dat_actv_2_7_valid(dat2_actv_pvld[7]),
.io_dat_actv_2_7_bits_nz(dat2_actv_nz[7]),
.io_dat_actv_2_7_bits_data(dat2_actv_data[63:56]),

.io_dat_actv_2_8_valid(dat2_actv_pvld[8]),
.io_dat_actv_2_8_bits_nz(dat2_actv_nz[8]),
.io_dat_actv_2_8_bits_data(dat2_actv_data[71:64]),

.io_dat_actv_2_9_valid(dat2_actv_pvld[9]),
.io_dat_actv_2_9_bits_nz(dat2_actv_nz[9]),
.io_dat_actv_2_9_bits_data(dat2_actv_data[79:72]),

.io_dat_actv_2_10_valid(dat2_actv_pvld[10]),
.io_dat_actv_2_10_bits_nz(dat2_actv_nz[10]),
.io_dat_actv_2_10_bits_data(dat2_actv_data[87:80]),

.io_dat_actv_2_11_valid(dat2_actv_pvld[11]),
.io_dat_actv_2_11_bits_nz(dat2_actv_nz[11]),
.io_dat_actv_2_11_bits_data(dat2_actv_data[95:88]),

.io_dat_actv_2_12_valid(dat2_actv_pvld[12]),
.io_dat_actv_2_12_bits_nz(dat2_actv_nz[12]),
.io_dat_actv_2_12_bits_data(dat2_actv_data[103:96]),

.io_dat_actv_2_13_valid(dat2_actv_pvld[13]),
.io_dat_actv_2_13_bits_nz(dat2_actv_nz[13]),
.io_dat_actv_2_13_bits_data(dat2_actv_data[111:104]),

.io_dat_actv_2_14_valid(dat2_actv_pvld[14]),
.io_dat_actv_2_14_bits_nz(dat2_actv_nz[14]),
.io_dat_actv_2_14_bits_data(dat2_actv_data[119:112]),

.io_dat_actv_2_15_valid(dat2_actv_pvld[15]),
.io_dat_actv_2_15_bits_nz(dat2_actv_nz[15]),
.io_dat_actv_2_15_bits_data(dat2_actv_data[127:120]),

.io_dat_actv_2_16_valid(dat2_actv_pvld[16]),
.io_dat_actv_2_16_bits_nz(dat2_actv_nz[16]),
.io_dat_actv_2_16_bits_data(dat2_actv_data[135:128]),

.io_dat_actv_2_17_valid(dat2_actv_pvld[17]),
.io_dat_actv_2_17_bits_nz(dat2_actv_nz[17]),
.io_dat_actv_2_17_bits_data(dat2_actv_data[143:136]),

.io_dat_actv_2_18_valid(dat2_actv_pvld[18]),
.io_dat_actv_2_18_bits_nz(dat2_actv_nz[18]),
.io_dat_actv_2_18_bits_data(dat2_actv_data[151:144]),

.io_dat_actv_2_19_valid(dat2_actv_pvld[19]),
.io_dat_actv_2_19_bits_nz(dat2_actv_nz[19]),
.io_dat_actv_2_19_bits_data(dat2_actv_data[159:152]),

.io_dat_actv_2_20_valid(dat2_actv_pvld[20]),
.io_dat_actv_2_20_bits_nz(dat2_actv_nz[20]),
.io_dat_actv_2_20_bits_data(dat2_actv_data[167:160]),

.io_dat_actv_2_21_valid(dat2_actv_pvld[21]),
.io_dat_actv_2_21_bits_nz(dat2_actv_nz[21]),
.io_dat_actv_2_21_bits_data(dat2_actv_data[175:168]),

.io_dat_actv_2_22_valid(dat2_actv_pvld[22]),
.io_dat_actv_2_22_bits_nz(dat2_actv_nz[22]),
.io_dat_actv_2_22_bits_data(dat2_actv_data[183:176]),

.io_dat_actv_2_23_valid(dat2_actv_pvld[23]),
.io_dat_actv_2_23_bits_nz(dat2_actv_nz[23]),
.io_dat_actv_2_23_bits_data(dat2_actv_data[191:184]),

.io_dat_actv_2_24_valid(dat2_actv_pvld[24]),
.io_dat_actv_2_24_bits_nz(dat2_actv_nz[24]),
.io_dat_actv_2_24_bits_data(dat2_actv_data[199:192]),

.io_dat_actv_2_25_valid(dat2_actv_pvld[25]),
.io_dat_actv_2_25_bits_nz(dat2_actv_nz[25]),
.io_dat_actv_2_25_bits_data(dat2_actv_data[207:200]),

.io_dat_actv_2_26_valid(dat2_actv_pvld[26]),
.io_dat_actv_2_26_bits_nz(dat2_actv_nz[26]),
.io_dat_actv_2_26_bits_data(dat2_actv_data[215:208]),

.io_dat_actv_2_27_valid(dat2_actv_pvld[27]),
.io_dat_actv_2_27_bits_nz(dat2_actv_nz[27]),
.io_dat_actv_2_27_bits_data(dat2_actv_data[223:216]),

.io_dat_actv_2_28_valid(dat2_actv_pvld[28]),
.io_dat_actv_2_28_bits_nz(dat2_actv_nz[28]),
.io_dat_actv_2_28_bits_data(dat2_actv_data[231:224]),

.io_dat_actv_2_29_valid(dat2_actv_pvld[29]),
.io_dat_actv_2_29_bits_nz(dat2_actv_nz[29]),
.io_dat_actv_2_29_bits_data(dat2_actv_data[239:232]),

.io_dat_actv_2_30_valid(dat2_actv_pvld[30]),
.io_dat_actv_2_30_bits_nz(dat2_actv_nz[30]),
.io_dat_actv_2_30_bits_data(dat2_actv_data[247:240]),

.io_dat_actv_2_31_valid(dat2_actv_pvld[31]),
.io_dat_actv_2_31_bits_nz(dat2_actv_nz[31]),
.io_dat_actv_2_31_bits_data(dat2_actv_data[255:248]),

.io_dat_actv_2_32_valid(dat2_actv_pvld[32]),
.io_dat_actv_2_32_bits_nz(dat2_actv_nz[32]),
.io_dat_actv_2_32_bits_data(dat2_actv_data[263:256]),

.io_dat_actv_2_33_valid(dat2_actv_pvld[33]),
.io_dat_actv_2_33_bits_nz(dat2_actv_nz[33]),
.io_dat_actv_2_33_bits_data(dat2_actv_data[271:264]),

.io_dat_actv_2_34_valid(dat2_actv_pvld[34]),
.io_dat_actv_2_34_bits_nz(dat2_actv_nz[34]),
.io_dat_actv_2_34_bits_data(dat2_actv_data[279:272]),

.io_dat_actv_2_35_valid(dat2_actv_pvld[35]),
.io_dat_actv_2_35_bits_nz(dat2_actv_nz[35]),
.io_dat_actv_2_35_bits_data(dat2_actv_data[287:280]),

.io_dat_actv_2_36_valid(dat2_actv_pvld[36]),
.io_dat_actv_2_36_bits_nz(dat2_actv_nz[36]),
.io_dat_actv_2_36_bits_data(dat2_actv_data[295:288]),

.io_dat_actv_2_37_valid(dat2_actv_pvld[37]),
.io_dat_actv_2_37_bits_nz(dat2_actv_nz[37]),
.io_dat_actv_2_37_bits_data(dat2_actv_data[303:296]),

.io_dat_actv_2_38_valid(dat2_actv_pvld[38]),
.io_dat_actv_2_38_bits_nz(dat2_actv_nz[38]),
.io_dat_actv_2_38_bits_data(dat2_actv_data[311:304]),

.io_dat_actv_2_39_valid(dat2_actv_pvld[39]),
.io_dat_actv_2_39_bits_nz(dat2_actv_nz[39]),
.io_dat_actv_2_39_bits_data(dat2_actv_data[319:312]),

.io_dat_actv_2_40_valid(dat2_actv_pvld[40]),
.io_dat_actv_2_40_bits_nz(dat2_actv_nz[40]),
.io_dat_actv_2_40_bits_data(dat2_actv_data[327:320]),

.io_dat_actv_2_41_valid(dat2_actv_pvld[41]),
.io_dat_actv_2_41_bits_nz(dat2_actv_nz[41]),
.io_dat_actv_2_41_bits_data(dat2_actv_data[335:328]),

.io_dat_actv_2_42_valid(dat2_actv_pvld[42]),
.io_dat_actv_2_42_bits_nz(dat2_actv_nz[42]),
.io_dat_actv_2_42_bits_data(dat2_actv_data[343:336]),

.io_dat_actv_2_43_valid(dat2_actv_pvld[43]),
.io_dat_actv_2_43_bits_nz(dat2_actv_nz[43]),
.io_dat_actv_2_43_bits_data(dat2_actv_data[351:344]),

.io_dat_actv_2_44_valid(dat2_actv_pvld[44]),
.io_dat_actv_2_44_bits_nz(dat2_actv_nz[44]),
.io_dat_actv_2_44_bits_data(dat2_actv_data[359:352]),

.io_dat_actv_2_45_valid(dat2_actv_pvld[45]),
.io_dat_actv_2_45_bits_nz(dat2_actv_nz[45]),
.io_dat_actv_2_45_bits_data(dat2_actv_data[367:360]),

.io_dat_actv_2_46_valid(dat2_actv_pvld[46]),
.io_dat_actv_2_46_bits_nz(dat2_actv_nz[46]),
.io_dat_actv_2_46_bits_data(dat2_actv_data[375:368]),

.io_dat_actv_2_47_valid(dat2_actv_pvld[47]),
.io_dat_actv_2_47_bits_nz(dat2_actv_nz[47]),
.io_dat_actv_2_47_bits_data(dat2_actv_data[383:376]),

.io_dat_actv_2_48_valid(dat2_actv_pvld[48]),
.io_dat_actv_2_48_bits_nz(dat2_actv_nz[48]),
.io_dat_actv_2_48_bits_data(dat2_actv_data[391:384]),

.io_dat_actv_2_49_valid(dat2_actv_pvld[49]),
.io_dat_actv_2_49_bits_nz(dat2_actv_nz[49]),
.io_dat_actv_2_49_bits_data(dat2_actv_data[399:392]),

.io_dat_actv_2_50_valid(dat2_actv_pvld[50]),
.io_dat_actv_2_50_bits_nz(dat2_actv_nz[50]),
.io_dat_actv_2_50_bits_data(dat2_actv_data[407:400]),

.io_dat_actv_2_51_valid(dat2_actv_pvld[51]),
.io_dat_actv_2_51_bits_nz(dat2_actv_nz[51]),
.io_dat_actv_2_51_bits_data(dat2_actv_data[415:408]),

.io_dat_actv_2_52_valid(dat2_actv_pvld[52]),
.io_dat_actv_2_52_bits_nz(dat2_actv_nz[52]),
.io_dat_actv_2_52_bits_data(dat2_actv_data[423:416]),

.io_dat_actv_2_53_valid(dat2_actv_pvld[53]),
.io_dat_actv_2_53_bits_nz(dat2_actv_nz[53]),
.io_dat_actv_2_53_bits_data(dat2_actv_data[431:424]),

.io_dat_actv_2_54_valid(dat2_actv_pvld[54]),
.io_dat_actv_2_54_bits_nz(dat2_actv_nz[54]),
.io_dat_actv_2_54_bits_data(dat2_actv_data[439:432]),

.io_dat_actv_2_55_valid(dat2_actv_pvld[55]),
.io_dat_actv_2_55_bits_nz(dat2_actv_nz[55]),
.io_dat_actv_2_55_bits_data(dat2_actv_data[447:440]),

.io_dat_actv_2_56_valid(dat2_actv_pvld[56]),
.io_dat_actv_2_56_bits_nz(dat2_actv_nz[56]),
.io_dat_actv_2_56_bits_data(dat2_actv_data[455:448]),

.io_dat_actv_2_57_valid(dat2_actv_pvld[57]),
.io_dat_actv_2_57_bits_nz(dat2_actv_nz[57]),
.io_dat_actv_2_57_bits_data(dat2_actv_data[463:456]),

.io_dat_actv_2_58_valid(dat2_actv_pvld[58]),
.io_dat_actv_2_58_bits_nz(dat2_actv_nz[58]),
.io_dat_actv_2_58_bits_data(dat2_actv_data[471:464]),

.io_dat_actv_2_59_valid(dat2_actv_pvld[59]),
.io_dat_actv_2_59_bits_nz(dat2_actv_nz[59]),
.io_dat_actv_2_59_bits_data(dat2_actv_data[479:472]),

.io_dat_actv_2_60_valid(dat2_actv_pvld[60]),
.io_dat_actv_2_60_bits_nz(dat2_actv_nz[60]),
.io_dat_actv_2_60_bits_data(dat2_actv_data[487:480]),

.io_dat_actv_2_61_valid(dat2_actv_pvld[61]),
.io_dat_actv_2_61_bits_nz(dat2_actv_nz[61]),
.io_dat_actv_2_61_bits_data(dat2_actv_data[495:488]),

.io_dat_actv_2_62_valid(dat2_actv_pvld[62]),
.io_dat_actv_2_62_bits_nz(dat2_actv_nz[62]),
.io_dat_actv_2_62_bits_data(dat2_actv_data[503:496]),

.io_dat_actv_2_63_valid(dat2_actv_pvld[63]),
.io_dat_actv_2_63_bits_nz(dat2_actv_nz[63]),
.io_dat_actv_2_63_bits_data(dat2_actv_data[511:504]),

.io_dat_actv_3_0_valid(dat3_actv_pvld[0]),
.io_dat_actv_3_0_bits_nz(dat3_actv_nz[0]),
.io_dat_actv_3_0_bits_data(dat3_actv_data[7:0]),

.io_dat_actv_3_1_valid(dat3_actv_pvld[1]),
.io_dat_actv_3_1_bits_nz(dat3_actv_nz[1]),
.io_dat_actv_3_1_bits_data(dat3_actv_data[15:8]),

.io_dat_actv_3_2_valid(dat3_actv_pvld[2]),
.io_dat_actv_3_2_bits_nz(dat3_actv_nz[2]),
.io_dat_actv_3_2_bits_data(dat3_actv_data[23:16]),

.io_dat_actv_3_3_valid(dat3_actv_pvld[3]),
.io_dat_actv_3_3_bits_nz(dat3_actv_nz[3]),
.io_dat_actv_3_3_bits_data(dat3_actv_data[31:24]),

.io_dat_actv_3_4_valid(dat3_actv_pvld[4]),
.io_dat_actv_3_4_bits_nz(dat3_actv_nz[4]),
.io_dat_actv_3_4_bits_data(dat3_actv_data[39:32]),

.io_dat_actv_3_5_valid(dat3_actv_pvld[5]),
.io_dat_actv_3_5_bits_nz(dat3_actv_nz[5]),
.io_dat_actv_3_5_bits_data(dat3_actv_data[47:40]),

.io_dat_actv_3_6_valid(dat3_actv_pvld[6]),
.io_dat_actv_3_6_bits_nz(dat3_actv_nz[6]),
.io_dat_actv_3_6_bits_data(dat3_actv_data[55:48]),

.io_dat_actv_3_7_valid(dat3_actv_pvld[7]),
.io_dat_actv_3_7_bits_nz(dat3_actv_nz[7]),
.io_dat_actv_3_7_bits_data(dat3_actv_data[63:56]),

.io_dat_actv_3_8_valid(dat3_actv_pvld[8]),
.io_dat_actv_3_8_bits_nz(dat3_actv_nz[8]),
.io_dat_actv_3_8_bits_data(dat3_actv_data[71:64]),

.io_dat_actv_3_9_valid(dat3_actv_pvld[9]),
.io_dat_actv_3_9_bits_nz(dat3_actv_nz[9]),
.io_dat_actv_3_9_bits_data(dat3_actv_data[79:72]),

.io_dat_actv_3_10_valid(dat3_actv_pvld[10]),
.io_dat_actv_3_10_bits_nz(dat3_actv_nz[10]),
.io_dat_actv_3_10_bits_data(dat3_actv_data[87:80]),

.io_dat_actv_3_11_valid(dat3_actv_pvld[11]),
.io_dat_actv_3_11_bits_nz(dat3_actv_nz[11]),
.io_dat_actv_3_11_bits_data(dat3_actv_data[95:88]),

.io_dat_actv_3_12_valid(dat3_actv_pvld[12]),
.io_dat_actv_3_12_bits_nz(dat3_actv_nz[12]),
.io_dat_actv_3_12_bits_data(dat3_actv_data[103:96]),

.io_dat_actv_3_13_valid(dat3_actv_pvld[13]),
.io_dat_actv_3_13_bits_nz(dat3_actv_nz[13]),
.io_dat_actv_3_13_bits_data(dat3_actv_data[111:104]),

.io_dat_actv_3_14_valid(dat3_actv_pvld[14]),
.io_dat_actv_3_14_bits_nz(dat3_actv_nz[14]),
.io_dat_actv_3_14_bits_data(dat3_actv_data[119:112]),

.io_dat_actv_3_15_valid(dat3_actv_pvld[15]),
.io_dat_actv_3_15_bits_nz(dat3_actv_nz[15]),
.io_dat_actv_3_15_bits_data(dat3_actv_data[127:120]),

.io_dat_actv_3_16_valid(dat3_actv_pvld[16]),
.io_dat_actv_3_16_bits_nz(dat3_actv_nz[16]),
.io_dat_actv_3_16_bits_data(dat3_actv_data[135:128]),

.io_dat_actv_3_17_valid(dat3_actv_pvld[17]),
.io_dat_actv_3_17_bits_nz(dat3_actv_nz[17]),
.io_dat_actv_3_17_bits_data(dat3_actv_data[143:136]),

.io_dat_actv_3_18_valid(dat3_actv_pvld[18]),
.io_dat_actv_3_18_bits_nz(dat3_actv_nz[18]),
.io_dat_actv_3_18_bits_data(dat3_actv_data[151:144]),

.io_dat_actv_3_19_valid(dat3_actv_pvld[19]),
.io_dat_actv_3_19_bits_nz(dat3_actv_nz[19]),
.io_dat_actv_3_19_bits_data(dat3_actv_data[159:152]),

.io_dat_actv_3_20_valid(dat3_actv_pvld[20]),
.io_dat_actv_3_20_bits_nz(dat3_actv_nz[20]),
.io_dat_actv_3_20_bits_data(dat3_actv_data[167:160]),

.io_dat_actv_3_21_valid(dat3_actv_pvld[21]),
.io_dat_actv_3_21_bits_nz(dat3_actv_nz[21]),
.io_dat_actv_3_21_bits_data(dat3_actv_data[175:168]),

.io_dat_actv_3_22_valid(dat3_actv_pvld[22]),
.io_dat_actv_3_22_bits_nz(dat3_actv_nz[22]),
.io_dat_actv_3_22_bits_data(dat3_actv_data[183:176]),

.io_dat_actv_3_23_valid(dat3_actv_pvld[23]),
.io_dat_actv_3_23_bits_nz(dat3_actv_nz[23]),
.io_dat_actv_3_23_bits_data(dat3_actv_data[191:184]),

.io_dat_actv_3_24_valid(dat3_actv_pvld[24]),
.io_dat_actv_3_24_bits_nz(dat3_actv_nz[24]),
.io_dat_actv_3_24_bits_data(dat3_actv_data[199:192]),

.io_dat_actv_3_25_valid(dat3_actv_pvld[25]),
.io_dat_actv_3_25_bits_nz(dat3_actv_nz[25]),
.io_dat_actv_3_25_bits_data(dat3_actv_data[207:200]),

.io_dat_actv_3_26_valid(dat3_actv_pvld[26]),
.io_dat_actv_3_26_bits_nz(dat3_actv_nz[26]),
.io_dat_actv_3_26_bits_data(dat3_actv_data[215:208]),

.io_dat_actv_3_27_valid(dat3_actv_pvld[27]),
.io_dat_actv_3_27_bits_nz(dat3_actv_nz[27]),
.io_dat_actv_3_27_bits_data(dat3_actv_data[223:216]),

.io_dat_actv_3_28_valid(dat3_actv_pvld[28]),
.io_dat_actv_3_28_bits_nz(dat3_actv_nz[28]),
.io_dat_actv_3_28_bits_data(dat3_actv_data[231:224]),

.io_dat_actv_3_29_valid(dat3_actv_pvld[29]),
.io_dat_actv_3_29_bits_nz(dat3_actv_nz[29]),
.io_dat_actv_3_29_bits_data(dat3_actv_data[239:232]),

.io_dat_actv_3_30_valid(dat3_actv_pvld[30]),
.io_dat_actv_3_30_bits_nz(dat3_actv_nz[30]),
.io_dat_actv_3_30_bits_data(dat3_actv_data[247:240]),

.io_dat_actv_3_31_valid(dat3_actv_pvld[31]),
.io_dat_actv_3_31_bits_nz(dat3_actv_nz[31]),
.io_dat_actv_3_31_bits_data(dat3_actv_data[255:248]),

.io_dat_actv_3_32_valid(dat3_actv_pvld[32]),
.io_dat_actv_3_32_bits_nz(dat3_actv_nz[32]),
.io_dat_actv_3_32_bits_data(dat3_actv_data[263:256]),

.io_dat_actv_3_33_valid(dat3_actv_pvld[33]),
.io_dat_actv_3_33_bits_nz(dat3_actv_nz[33]),
.io_dat_actv_3_33_bits_data(dat3_actv_data[271:264]),

.io_dat_actv_3_34_valid(dat3_actv_pvld[34]),
.io_dat_actv_3_34_bits_nz(dat3_actv_nz[34]),
.io_dat_actv_3_34_bits_data(dat3_actv_data[279:272]),

.io_dat_actv_3_35_valid(dat3_actv_pvld[35]),
.io_dat_actv_3_35_bits_nz(dat3_actv_nz[35]),
.io_dat_actv_3_35_bits_data(dat3_actv_data[287:280]),

.io_dat_actv_3_36_valid(dat3_actv_pvld[36]),
.io_dat_actv_3_36_bits_nz(dat3_actv_nz[36]),
.io_dat_actv_3_36_bits_data(dat3_actv_data[295:288]),

.io_dat_actv_3_37_valid(dat3_actv_pvld[37]),
.io_dat_actv_3_37_bits_nz(dat3_actv_nz[37]),
.io_dat_actv_3_37_bits_data(dat3_actv_data[303:296]),

.io_dat_actv_3_38_valid(dat3_actv_pvld[38]),
.io_dat_actv_3_38_bits_nz(dat3_actv_nz[38]),
.io_dat_actv_3_38_bits_data(dat3_actv_data[311:304]),

.io_dat_actv_3_39_valid(dat3_actv_pvld[39]),
.io_dat_actv_3_39_bits_nz(dat3_actv_nz[39]),
.io_dat_actv_3_39_bits_data(dat3_actv_data[319:312]),

.io_dat_actv_3_40_valid(dat3_actv_pvld[40]),
.io_dat_actv_3_40_bits_nz(dat3_actv_nz[40]),
.io_dat_actv_3_40_bits_data(dat3_actv_data[327:320]),

.io_dat_actv_3_41_valid(dat3_actv_pvld[41]),
.io_dat_actv_3_41_bits_nz(dat3_actv_nz[41]),
.io_dat_actv_3_41_bits_data(dat3_actv_data[335:328]),

.io_dat_actv_3_42_valid(dat3_actv_pvld[42]),
.io_dat_actv_3_42_bits_nz(dat3_actv_nz[42]),
.io_dat_actv_3_42_bits_data(dat3_actv_data[343:336]),

.io_dat_actv_3_43_valid(dat3_actv_pvld[43]),
.io_dat_actv_3_43_bits_nz(dat3_actv_nz[43]),
.io_dat_actv_3_43_bits_data(dat3_actv_data[351:344]),

.io_dat_actv_3_44_valid(dat3_actv_pvld[44]),
.io_dat_actv_3_44_bits_nz(dat3_actv_nz[44]),
.io_dat_actv_3_44_bits_data(dat3_actv_data[359:352]),

.io_dat_actv_3_45_valid(dat3_actv_pvld[45]),
.io_dat_actv_3_45_bits_nz(dat3_actv_nz[45]),
.io_dat_actv_3_45_bits_data(dat3_actv_data[367:360]),

.io_dat_actv_3_46_valid(dat3_actv_pvld[46]),
.io_dat_actv_3_46_bits_nz(dat3_actv_nz[46]),
.io_dat_actv_3_46_bits_data(dat3_actv_data[375:368]),

.io_dat_actv_3_47_valid(dat3_actv_pvld[47]),
.io_dat_actv_3_47_bits_nz(dat3_actv_nz[47]),
.io_dat_actv_3_47_bits_data(dat3_actv_data[383:376]),

.io_dat_actv_3_48_valid(dat3_actv_pvld[48]),
.io_dat_actv_3_48_bits_nz(dat3_actv_nz[48]),
.io_dat_actv_3_48_bits_data(dat3_actv_data[391:384]),

.io_dat_actv_3_49_valid(dat3_actv_pvld[49]),
.io_dat_actv_3_49_bits_nz(dat3_actv_nz[49]),
.io_dat_actv_3_49_bits_data(dat3_actv_data[399:392]),

.io_dat_actv_3_50_valid(dat3_actv_pvld[50]),
.io_dat_actv_3_50_bits_nz(dat3_actv_nz[50]),
.io_dat_actv_3_50_bits_data(dat3_actv_data[407:400]),

.io_dat_actv_3_51_valid(dat3_actv_pvld[51]),
.io_dat_actv_3_51_bits_nz(dat3_actv_nz[51]),
.io_dat_actv_3_51_bits_data(dat3_actv_data[415:408]),

.io_dat_actv_3_52_valid(dat3_actv_pvld[52]),
.io_dat_actv_3_52_bits_nz(dat3_actv_nz[52]),
.io_dat_actv_3_52_bits_data(dat3_actv_data[423:416]),

.io_dat_actv_3_53_valid(dat3_actv_pvld[53]),
.io_dat_actv_3_53_bits_nz(dat3_actv_nz[53]),
.io_dat_actv_3_53_bits_data(dat3_actv_data[431:424]),

.io_dat_actv_3_54_valid(dat3_actv_pvld[54]),
.io_dat_actv_3_54_bits_nz(dat3_actv_nz[54]),
.io_dat_actv_3_54_bits_data(dat3_actv_data[439:432]),

.io_dat_actv_3_55_valid(dat3_actv_pvld[55]),
.io_dat_actv_3_55_bits_nz(dat3_actv_nz[55]),
.io_dat_actv_3_55_bits_data(dat3_actv_data[447:440]),

.io_dat_actv_3_56_valid(dat3_actv_pvld[56]),
.io_dat_actv_3_56_bits_nz(dat3_actv_nz[56]),
.io_dat_actv_3_56_bits_data(dat3_actv_data[455:448]),

.io_dat_actv_3_57_valid(dat3_actv_pvld[57]),
.io_dat_actv_3_57_bits_nz(dat3_actv_nz[57]),
.io_dat_actv_3_57_bits_data(dat3_actv_data[463:456]),

.io_dat_actv_3_58_valid(dat3_actv_pvld[58]),
.io_dat_actv_3_58_bits_nz(dat3_actv_nz[58]),
.io_dat_actv_3_58_bits_data(dat3_actv_data[471:464]),

.io_dat_actv_3_59_valid(dat3_actv_pvld[59]),
.io_dat_actv_3_59_bits_nz(dat3_actv_nz[59]),
.io_dat_actv_3_59_bits_data(dat3_actv_data[479:472]),

.io_dat_actv_3_60_valid(dat3_actv_pvld[60]),
.io_dat_actv_3_60_bits_nz(dat3_actv_nz[60]),
.io_dat_actv_3_60_bits_data(dat3_actv_data[487:480]),

.io_dat_actv_3_61_valid(dat3_actv_pvld[61]),
.io_dat_actv_3_61_bits_nz(dat3_actv_nz[61]),
.io_dat_actv_3_61_bits_data(dat3_actv_data[495:488]),

.io_dat_actv_3_62_valid(dat3_actv_pvld[62]),
.io_dat_actv_3_62_bits_nz(dat3_actv_nz[62]),
.io_dat_actv_3_62_bits_data(dat3_actv_data[503:496]),

.io_dat_actv_3_63_valid(dat3_actv_pvld[63]),
.io_dat_actv_3_63_bits_nz(dat3_actv_nz[63]),
.io_dat_actv_3_63_bits_data(dat3_actv_data[511:504]),

.io_dat_actv_4_0_valid(dat4_actv_pvld[0]),
.io_dat_actv_4_0_bits_nz(dat4_actv_nz[0]),
.io_dat_actv_4_0_bits_data(dat4_actv_data[7:0]),

.io_dat_actv_4_1_valid(dat4_actv_pvld[1]),
.io_dat_actv_4_1_bits_nz(dat4_actv_nz[1]),
.io_dat_actv_4_1_bits_data(dat4_actv_data[15:8]),

.io_dat_actv_4_2_valid(dat4_actv_pvld[2]),
.io_dat_actv_4_2_bits_nz(dat4_actv_nz[2]),
.io_dat_actv_4_2_bits_data(dat4_actv_data[23:16]),

.io_dat_actv_4_3_valid(dat4_actv_pvld[3]),
.io_dat_actv_4_3_bits_nz(dat4_actv_nz[3]),
.io_dat_actv_4_3_bits_data(dat4_actv_data[31:24]),

.io_dat_actv_4_4_valid(dat4_actv_pvld[4]),
.io_dat_actv_4_4_bits_nz(dat4_actv_nz[4]),
.io_dat_actv_4_4_bits_data(dat4_actv_data[39:32]),

.io_dat_actv_4_5_valid(dat4_actv_pvld[5]),
.io_dat_actv_4_5_bits_nz(dat4_actv_nz[5]),
.io_dat_actv_4_5_bits_data(dat4_actv_data[47:40]),

.io_dat_actv_4_6_valid(dat4_actv_pvld[6]),
.io_dat_actv_4_6_bits_nz(dat4_actv_nz[6]),
.io_dat_actv_4_6_bits_data(dat4_actv_data[55:48]),

.io_dat_actv_4_7_valid(dat4_actv_pvld[7]),
.io_dat_actv_4_7_bits_nz(dat4_actv_nz[7]),
.io_dat_actv_4_7_bits_data(dat4_actv_data[63:56]),

.io_dat_actv_4_8_valid(dat4_actv_pvld[8]),
.io_dat_actv_4_8_bits_nz(dat4_actv_nz[8]),
.io_dat_actv_4_8_bits_data(dat4_actv_data[71:64]),

.io_dat_actv_4_9_valid(dat4_actv_pvld[9]),
.io_dat_actv_4_9_bits_nz(dat4_actv_nz[9]),
.io_dat_actv_4_9_bits_data(dat4_actv_data[79:72]),

.io_dat_actv_4_10_valid(dat4_actv_pvld[10]),
.io_dat_actv_4_10_bits_nz(dat4_actv_nz[10]),
.io_dat_actv_4_10_bits_data(dat4_actv_data[87:80]),

.io_dat_actv_4_11_valid(dat4_actv_pvld[11]),
.io_dat_actv_4_11_bits_nz(dat4_actv_nz[11]),
.io_dat_actv_4_11_bits_data(dat4_actv_data[95:88]),

.io_dat_actv_4_12_valid(dat4_actv_pvld[12]),
.io_dat_actv_4_12_bits_nz(dat4_actv_nz[12]),
.io_dat_actv_4_12_bits_data(dat4_actv_data[103:96]),

.io_dat_actv_4_13_valid(dat4_actv_pvld[13]),
.io_dat_actv_4_13_bits_nz(dat4_actv_nz[13]),
.io_dat_actv_4_13_bits_data(dat4_actv_data[111:104]),

.io_dat_actv_4_14_valid(dat4_actv_pvld[14]),
.io_dat_actv_4_14_bits_nz(dat4_actv_nz[14]),
.io_dat_actv_4_14_bits_data(dat4_actv_data[119:112]),

.io_dat_actv_4_15_valid(dat4_actv_pvld[15]),
.io_dat_actv_4_15_bits_nz(dat4_actv_nz[15]),
.io_dat_actv_4_15_bits_data(dat4_actv_data[127:120]),

.io_dat_actv_4_16_valid(dat4_actv_pvld[16]),
.io_dat_actv_4_16_bits_nz(dat4_actv_nz[16]),
.io_dat_actv_4_16_bits_data(dat4_actv_data[135:128]),

.io_dat_actv_4_17_valid(dat4_actv_pvld[17]),
.io_dat_actv_4_17_bits_nz(dat4_actv_nz[17]),
.io_dat_actv_4_17_bits_data(dat4_actv_data[143:136]),

.io_dat_actv_4_18_valid(dat4_actv_pvld[18]),
.io_dat_actv_4_18_bits_nz(dat4_actv_nz[18]),
.io_dat_actv_4_18_bits_data(dat4_actv_data[151:144]),

.io_dat_actv_4_19_valid(dat4_actv_pvld[19]),
.io_dat_actv_4_19_bits_nz(dat4_actv_nz[19]),
.io_dat_actv_4_19_bits_data(dat4_actv_data[159:152]),

.io_dat_actv_4_20_valid(dat4_actv_pvld[20]),
.io_dat_actv_4_20_bits_nz(dat4_actv_nz[20]),
.io_dat_actv_4_20_bits_data(dat4_actv_data[167:160]),

.io_dat_actv_4_21_valid(dat4_actv_pvld[21]),
.io_dat_actv_4_21_bits_nz(dat4_actv_nz[21]),
.io_dat_actv_4_21_bits_data(dat4_actv_data[175:168]),

.io_dat_actv_4_22_valid(dat4_actv_pvld[22]),
.io_dat_actv_4_22_bits_nz(dat4_actv_nz[22]),
.io_dat_actv_4_22_bits_data(dat4_actv_data[183:176]),

.io_dat_actv_4_23_valid(dat4_actv_pvld[23]),
.io_dat_actv_4_23_bits_nz(dat4_actv_nz[23]),
.io_dat_actv_4_23_bits_data(dat4_actv_data[191:184]),

.io_dat_actv_4_24_valid(dat4_actv_pvld[24]),
.io_dat_actv_4_24_bits_nz(dat4_actv_nz[24]),
.io_dat_actv_4_24_bits_data(dat4_actv_data[199:192]),

.io_dat_actv_4_25_valid(dat4_actv_pvld[25]),
.io_dat_actv_4_25_bits_nz(dat4_actv_nz[25]),
.io_dat_actv_4_25_bits_data(dat4_actv_data[207:200]),

.io_dat_actv_4_26_valid(dat4_actv_pvld[26]),
.io_dat_actv_4_26_bits_nz(dat4_actv_nz[26]),
.io_dat_actv_4_26_bits_data(dat4_actv_data[215:208]),

.io_dat_actv_4_27_valid(dat4_actv_pvld[27]),
.io_dat_actv_4_27_bits_nz(dat4_actv_nz[27]),
.io_dat_actv_4_27_bits_data(dat4_actv_data[223:216]),

.io_dat_actv_4_28_valid(dat4_actv_pvld[28]),
.io_dat_actv_4_28_bits_nz(dat4_actv_nz[28]),
.io_dat_actv_4_28_bits_data(dat4_actv_data[231:224]),

.io_dat_actv_4_29_valid(dat4_actv_pvld[29]),
.io_dat_actv_4_29_bits_nz(dat4_actv_nz[29]),
.io_dat_actv_4_29_bits_data(dat4_actv_data[239:232]),

.io_dat_actv_4_30_valid(dat4_actv_pvld[30]),
.io_dat_actv_4_30_bits_nz(dat4_actv_nz[30]),
.io_dat_actv_4_30_bits_data(dat4_actv_data[247:240]),

.io_dat_actv_4_31_valid(dat4_actv_pvld[31]),
.io_dat_actv_4_31_bits_nz(dat4_actv_nz[31]),
.io_dat_actv_4_31_bits_data(dat4_actv_data[255:248]),

.io_dat_actv_4_32_valid(dat4_actv_pvld[32]),
.io_dat_actv_4_32_bits_nz(dat4_actv_nz[32]),
.io_dat_actv_4_32_bits_data(dat4_actv_data[263:256]),

.io_dat_actv_4_33_valid(dat4_actv_pvld[33]),
.io_dat_actv_4_33_bits_nz(dat4_actv_nz[33]),
.io_dat_actv_4_33_bits_data(dat4_actv_data[271:264]),

.io_dat_actv_4_34_valid(dat4_actv_pvld[34]),
.io_dat_actv_4_34_bits_nz(dat4_actv_nz[34]),
.io_dat_actv_4_34_bits_data(dat4_actv_data[279:272]),

.io_dat_actv_4_35_valid(dat4_actv_pvld[35]),
.io_dat_actv_4_35_bits_nz(dat4_actv_nz[35]),
.io_dat_actv_4_35_bits_data(dat4_actv_data[287:280]),

.io_dat_actv_4_36_valid(dat4_actv_pvld[36]),
.io_dat_actv_4_36_bits_nz(dat4_actv_nz[36]),
.io_dat_actv_4_36_bits_data(dat4_actv_data[295:288]),

.io_dat_actv_4_37_valid(dat4_actv_pvld[37]),
.io_dat_actv_4_37_bits_nz(dat4_actv_nz[37]),
.io_dat_actv_4_37_bits_data(dat4_actv_data[303:296]),

.io_dat_actv_4_38_valid(dat4_actv_pvld[38]),
.io_dat_actv_4_38_bits_nz(dat4_actv_nz[38]),
.io_dat_actv_4_38_bits_data(dat4_actv_data[311:304]),

.io_dat_actv_4_39_valid(dat4_actv_pvld[39]),
.io_dat_actv_4_39_bits_nz(dat4_actv_nz[39]),
.io_dat_actv_4_39_bits_data(dat4_actv_data[319:312]),

.io_dat_actv_4_40_valid(dat4_actv_pvld[40]),
.io_dat_actv_4_40_bits_nz(dat4_actv_nz[40]),
.io_dat_actv_4_40_bits_data(dat4_actv_data[327:320]),

.io_dat_actv_4_41_valid(dat4_actv_pvld[41]),
.io_dat_actv_4_41_bits_nz(dat4_actv_nz[41]),
.io_dat_actv_4_41_bits_data(dat4_actv_data[335:328]),

.io_dat_actv_4_42_valid(dat4_actv_pvld[42]),
.io_dat_actv_4_42_bits_nz(dat4_actv_nz[42]),
.io_dat_actv_4_42_bits_data(dat4_actv_data[343:336]),

.io_dat_actv_4_43_valid(dat4_actv_pvld[43]),
.io_dat_actv_4_43_bits_nz(dat4_actv_nz[43]),
.io_dat_actv_4_43_bits_data(dat4_actv_data[351:344]),

.io_dat_actv_4_44_valid(dat4_actv_pvld[44]),
.io_dat_actv_4_44_bits_nz(dat4_actv_nz[44]),
.io_dat_actv_4_44_bits_data(dat4_actv_data[359:352]),

.io_dat_actv_4_45_valid(dat4_actv_pvld[45]),
.io_dat_actv_4_45_bits_nz(dat4_actv_nz[45]),
.io_dat_actv_4_45_bits_data(dat4_actv_data[367:360]),

.io_dat_actv_4_46_valid(dat4_actv_pvld[46]),
.io_dat_actv_4_46_bits_nz(dat4_actv_nz[46]),
.io_dat_actv_4_46_bits_data(dat4_actv_data[375:368]),

.io_dat_actv_4_47_valid(dat4_actv_pvld[47]),
.io_dat_actv_4_47_bits_nz(dat4_actv_nz[47]),
.io_dat_actv_4_47_bits_data(dat4_actv_data[383:376]),

.io_dat_actv_4_48_valid(dat4_actv_pvld[48]),
.io_dat_actv_4_48_bits_nz(dat4_actv_nz[48]),
.io_dat_actv_4_48_bits_data(dat4_actv_data[391:384]),

.io_dat_actv_4_49_valid(dat4_actv_pvld[49]),
.io_dat_actv_4_49_bits_nz(dat4_actv_nz[49]),
.io_dat_actv_4_49_bits_data(dat4_actv_data[399:392]),

.io_dat_actv_4_50_valid(dat4_actv_pvld[50]),
.io_dat_actv_4_50_bits_nz(dat4_actv_nz[50]),
.io_dat_actv_4_50_bits_data(dat4_actv_data[407:400]),

.io_dat_actv_4_51_valid(dat4_actv_pvld[51]),
.io_dat_actv_4_51_bits_nz(dat4_actv_nz[51]),
.io_dat_actv_4_51_bits_data(dat4_actv_data[415:408]),

.io_dat_actv_4_52_valid(dat4_actv_pvld[52]),
.io_dat_actv_4_52_bits_nz(dat4_actv_nz[52]),
.io_dat_actv_4_52_bits_data(dat4_actv_data[423:416]),

.io_dat_actv_4_53_valid(dat4_actv_pvld[53]),
.io_dat_actv_4_53_bits_nz(dat4_actv_nz[53]),
.io_dat_actv_4_53_bits_data(dat4_actv_data[431:424]),

.io_dat_actv_4_54_valid(dat4_actv_pvld[54]),
.io_dat_actv_4_54_bits_nz(dat4_actv_nz[54]),
.io_dat_actv_4_54_bits_data(dat4_actv_data[439:432]),

.io_dat_actv_4_55_valid(dat4_actv_pvld[55]),
.io_dat_actv_4_55_bits_nz(dat4_actv_nz[55]),
.io_dat_actv_4_55_bits_data(dat4_actv_data[447:440]),

.io_dat_actv_4_56_valid(dat4_actv_pvld[56]),
.io_dat_actv_4_56_bits_nz(dat4_actv_nz[56]),
.io_dat_actv_4_56_bits_data(dat4_actv_data[455:448]),

.io_dat_actv_4_57_valid(dat4_actv_pvld[57]),
.io_dat_actv_4_57_bits_nz(dat4_actv_nz[57]),
.io_dat_actv_4_57_bits_data(dat4_actv_data[463:456]),

.io_dat_actv_4_58_valid(dat4_actv_pvld[58]),
.io_dat_actv_4_58_bits_nz(dat4_actv_nz[58]),
.io_dat_actv_4_58_bits_data(dat4_actv_data[471:464]),

.io_dat_actv_4_59_valid(dat4_actv_pvld[59]),
.io_dat_actv_4_59_bits_nz(dat4_actv_nz[59]),
.io_dat_actv_4_59_bits_data(dat4_actv_data[479:472]),

.io_dat_actv_4_60_valid(dat4_actv_pvld[60]),
.io_dat_actv_4_60_bits_nz(dat4_actv_nz[60]),
.io_dat_actv_4_60_bits_data(dat4_actv_data[487:480]),

.io_dat_actv_4_61_valid(dat4_actv_pvld[61]),
.io_dat_actv_4_61_bits_nz(dat4_actv_nz[61]),
.io_dat_actv_4_61_bits_data(dat4_actv_data[495:488]),

.io_dat_actv_4_62_valid(dat4_actv_pvld[62]),
.io_dat_actv_4_62_bits_nz(dat4_actv_nz[62]),
.io_dat_actv_4_62_bits_data(dat4_actv_data[503:496]),

.io_dat_actv_4_63_valid(dat4_actv_pvld[63]),
.io_dat_actv_4_63_bits_nz(dat4_actv_nz[63]),
.io_dat_actv_4_63_bits_data(dat4_actv_data[511:504]),

.io_dat_actv_5_0_valid(dat5_actv_pvld[0]),
.io_dat_actv_5_0_bits_nz(dat5_actv_nz[0]),
.io_dat_actv_5_0_bits_data(dat5_actv_data[7:0]),

.io_dat_actv_5_1_valid(dat5_actv_pvld[1]),
.io_dat_actv_5_1_bits_nz(dat5_actv_nz[1]),
.io_dat_actv_5_1_bits_data(dat5_actv_data[15:8]),

.io_dat_actv_5_2_valid(dat5_actv_pvld[2]),
.io_dat_actv_5_2_bits_nz(dat5_actv_nz[2]),
.io_dat_actv_5_2_bits_data(dat5_actv_data[23:16]),

.io_dat_actv_5_3_valid(dat5_actv_pvld[3]),
.io_dat_actv_5_3_bits_nz(dat5_actv_nz[3]),
.io_dat_actv_5_3_bits_data(dat5_actv_data[31:24]),

.io_dat_actv_5_4_valid(dat5_actv_pvld[4]),
.io_dat_actv_5_4_bits_nz(dat5_actv_nz[4]),
.io_dat_actv_5_4_bits_data(dat5_actv_data[39:32]),

.io_dat_actv_5_5_valid(dat5_actv_pvld[5]),
.io_dat_actv_5_5_bits_nz(dat5_actv_nz[5]),
.io_dat_actv_5_5_bits_data(dat5_actv_data[47:40]),

.io_dat_actv_5_6_valid(dat5_actv_pvld[6]),
.io_dat_actv_5_6_bits_nz(dat5_actv_nz[6]),
.io_dat_actv_5_6_bits_data(dat5_actv_data[55:48]),

.io_dat_actv_5_7_valid(dat5_actv_pvld[7]),
.io_dat_actv_5_7_bits_nz(dat5_actv_nz[7]),
.io_dat_actv_5_7_bits_data(dat5_actv_data[63:56]),

.io_dat_actv_5_8_valid(dat5_actv_pvld[8]),
.io_dat_actv_5_8_bits_nz(dat5_actv_nz[8]),
.io_dat_actv_5_8_bits_data(dat5_actv_data[71:64]),

.io_dat_actv_5_9_valid(dat5_actv_pvld[9]),
.io_dat_actv_5_9_bits_nz(dat5_actv_nz[9]),
.io_dat_actv_5_9_bits_data(dat5_actv_data[79:72]),

.io_dat_actv_5_10_valid(dat5_actv_pvld[10]),
.io_dat_actv_5_10_bits_nz(dat5_actv_nz[10]),
.io_dat_actv_5_10_bits_data(dat5_actv_data[87:80]),

.io_dat_actv_5_11_valid(dat5_actv_pvld[11]),
.io_dat_actv_5_11_bits_nz(dat5_actv_nz[11]),
.io_dat_actv_5_11_bits_data(dat5_actv_data[95:88]),

.io_dat_actv_5_12_valid(dat5_actv_pvld[12]),
.io_dat_actv_5_12_bits_nz(dat5_actv_nz[12]),
.io_dat_actv_5_12_bits_data(dat5_actv_data[103:96]),

.io_dat_actv_5_13_valid(dat5_actv_pvld[13]),
.io_dat_actv_5_13_bits_nz(dat5_actv_nz[13]),
.io_dat_actv_5_13_bits_data(dat5_actv_data[111:104]),

.io_dat_actv_5_14_valid(dat5_actv_pvld[14]),
.io_dat_actv_5_14_bits_nz(dat5_actv_nz[14]),
.io_dat_actv_5_14_bits_data(dat5_actv_data[119:112]),

.io_dat_actv_5_15_valid(dat5_actv_pvld[15]),
.io_dat_actv_5_15_bits_nz(dat5_actv_nz[15]),
.io_dat_actv_5_15_bits_data(dat5_actv_data[127:120]),

.io_dat_actv_5_16_valid(dat5_actv_pvld[16]),
.io_dat_actv_5_16_bits_nz(dat5_actv_nz[16]),
.io_dat_actv_5_16_bits_data(dat5_actv_data[135:128]),

.io_dat_actv_5_17_valid(dat5_actv_pvld[17]),
.io_dat_actv_5_17_bits_nz(dat5_actv_nz[17]),
.io_dat_actv_5_17_bits_data(dat5_actv_data[143:136]),

.io_dat_actv_5_18_valid(dat5_actv_pvld[18]),
.io_dat_actv_5_18_bits_nz(dat5_actv_nz[18]),
.io_dat_actv_5_18_bits_data(dat5_actv_data[151:144]),

.io_dat_actv_5_19_valid(dat5_actv_pvld[19]),
.io_dat_actv_5_19_bits_nz(dat5_actv_nz[19]),
.io_dat_actv_5_19_bits_data(dat5_actv_data[159:152]),

.io_dat_actv_5_20_valid(dat5_actv_pvld[20]),
.io_dat_actv_5_20_bits_nz(dat5_actv_nz[20]),
.io_dat_actv_5_20_bits_data(dat5_actv_data[167:160]),

.io_dat_actv_5_21_valid(dat5_actv_pvld[21]),
.io_dat_actv_5_21_bits_nz(dat5_actv_nz[21]),
.io_dat_actv_5_21_bits_data(dat5_actv_data[175:168]),

.io_dat_actv_5_22_valid(dat5_actv_pvld[22]),
.io_dat_actv_5_22_bits_nz(dat5_actv_nz[22]),
.io_dat_actv_5_22_bits_data(dat5_actv_data[183:176]),

.io_dat_actv_5_23_valid(dat5_actv_pvld[23]),
.io_dat_actv_5_23_bits_nz(dat5_actv_nz[23]),
.io_dat_actv_5_23_bits_data(dat5_actv_data[191:184]),

.io_dat_actv_5_24_valid(dat5_actv_pvld[24]),
.io_dat_actv_5_24_bits_nz(dat5_actv_nz[24]),
.io_dat_actv_5_24_bits_data(dat5_actv_data[199:192]),

.io_dat_actv_5_25_valid(dat5_actv_pvld[25]),
.io_dat_actv_5_25_bits_nz(dat5_actv_nz[25]),
.io_dat_actv_5_25_bits_data(dat5_actv_data[207:200]),

.io_dat_actv_5_26_valid(dat5_actv_pvld[26]),
.io_dat_actv_5_26_bits_nz(dat5_actv_nz[26]),
.io_dat_actv_5_26_bits_data(dat5_actv_data[215:208]),

.io_dat_actv_5_27_valid(dat5_actv_pvld[27]),
.io_dat_actv_5_27_bits_nz(dat5_actv_nz[27]),
.io_dat_actv_5_27_bits_data(dat5_actv_data[223:216]),

.io_dat_actv_5_28_valid(dat5_actv_pvld[28]),
.io_dat_actv_5_28_bits_nz(dat5_actv_nz[28]),
.io_dat_actv_5_28_bits_data(dat5_actv_data[231:224]),

.io_dat_actv_5_29_valid(dat5_actv_pvld[29]),
.io_dat_actv_5_29_bits_nz(dat5_actv_nz[29]),
.io_dat_actv_5_29_bits_data(dat5_actv_data[239:232]),

.io_dat_actv_5_30_valid(dat5_actv_pvld[30]),
.io_dat_actv_5_30_bits_nz(dat5_actv_nz[30]),
.io_dat_actv_5_30_bits_data(dat5_actv_data[247:240]),

.io_dat_actv_5_31_valid(dat5_actv_pvld[31]),
.io_dat_actv_5_31_bits_nz(dat5_actv_nz[31]),
.io_dat_actv_5_31_bits_data(dat5_actv_data[255:248]),

.io_dat_actv_5_32_valid(dat5_actv_pvld[32]),
.io_dat_actv_5_32_bits_nz(dat5_actv_nz[32]),
.io_dat_actv_5_32_bits_data(dat5_actv_data[263:256]),

.io_dat_actv_5_33_valid(dat5_actv_pvld[33]),
.io_dat_actv_5_33_bits_nz(dat5_actv_nz[33]),
.io_dat_actv_5_33_bits_data(dat5_actv_data[271:264]),

.io_dat_actv_5_34_valid(dat5_actv_pvld[34]),
.io_dat_actv_5_34_bits_nz(dat5_actv_nz[34]),
.io_dat_actv_5_34_bits_data(dat5_actv_data[279:272]),

.io_dat_actv_5_35_valid(dat5_actv_pvld[35]),
.io_dat_actv_5_35_bits_nz(dat5_actv_nz[35]),
.io_dat_actv_5_35_bits_data(dat5_actv_data[287:280]),

.io_dat_actv_5_36_valid(dat5_actv_pvld[36]),
.io_dat_actv_5_36_bits_nz(dat5_actv_nz[36]),
.io_dat_actv_5_36_bits_data(dat5_actv_data[295:288]),

.io_dat_actv_5_37_valid(dat5_actv_pvld[37]),
.io_dat_actv_5_37_bits_nz(dat5_actv_nz[37]),
.io_dat_actv_5_37_bits_data(dat5_actv_data[303:296]),

.io_dat_actv_5_38_valid(dat5_actv_pvld[38]),
.io_dat_actv_5_38_bits_nz(dat5_actv_nz[38]),
.io_dat_actv_5_38_bits_data(dat5_actv_data[311:304]),

.io_dat_actv_5_39_valid(dat5_actv_pvld[39]),
.io_dat_actv_5_39_bits_nz(dat5_actv_nz[39]),
.io_dat_actv_5_39_bits_data(dat5_actv_data[319:312]),

.io_dat_actv_5_40_valid(dat5_actv_pvld[40]),
.io_dat_actv_5_40_bits_nz(dat5_actv_nz[40]),
.io_dat_actv_5_40_bits_data(dat5_actv_data[327:320]),

.io_dat_actv_5_41_valid(dat5_actv_pvld[41]),
.io_dat_actv_5_41_bits_nz(dat5_actv_nz[41]),
.io_dat_actv_5_41_bits_data(dat5_actv_data[335:328]),

.io_dat_actv_5_42_valid(dat5_actv_pvld[42]),
.io_dat_actv_5_42_bits_nz(dat5_actv_nz[42]),
.io_dat_actv_5_42_bits_data(dat5_actv_data[343:336]),

.io_dat_actv_5_43_valid(dat5_actv_pvld[43]),
.io_dat_actv_5_43_bits_nz(dat5_actv_nz[43]),
.io_dat_actv_5_43_bits_data(dat5_actv_data[351:344]),

.io_dat_actv_5_44_valid(dat5_actv_pvld[44]),
.io_dat_actv_5_44_bits_nz(dat5_actv_nz[44]),
.io_dat_actv_5_44_bits_data(dat5_actv_data[359:352]),

.io_dat_actv_5_45_valid(dat5_actv_pvld[45]),
.io_dat_actv_5_45_bits_nz(dat5_actv_nz[45]),
.io_dat_actv_5_45_bits_data(dat5_actv_data[367:360]),

.io_dat_actv_5_46_valid(dat5_actv_pvld[46]),
.io_dat_actv_5_46_bits_nz(dat5_actv_nz[46]),
.io_dat_actv_5_46_bits_data(dat5_actv_data[375:368]),

.io_dat_actv_5_47_valid(dat5_actv_pvld[47]),
.io_dat_actv_5_47_bits_nz(dat5_actv_nz[47]),
.io_dat_actv_5_47_bits_data(dat5_actv_data[383:376]),

.io_dat_actv_5_48_valid(dat5_actv_pvld[48]),
.io_dat_actv_5_48_bits_nz(dat5_actv_nz[48]),
.io_dat_actv_5_48_bits_data(dat5_actv_data[391:384]),

.io_dat_actv_5_49_valid(dat5_actv_pvld[49]),
.io_dat_actv_5_49_bits_nz(dat5_actv_nz[49]),
.io_dat_actv_5_49_bits_data(dat5_actv_data[399:392]),

.io_dat_actv_5_50_valid(dat5_actv_pvld[50]),
.io_dat_actv_5_50_bits_nz(dat5_actv_nz[50]),
.io_dat_actv_5_50_bits_data(dat5_actv_data[407:400]),

.io_dat_actv_5_51_valid(dat5_actv_pvld[51]),
.io_dat_actv_5_51_bits_nz(dat5_actv_nz[51]),
.io_dat_actv_5_51_bits_data(dat5_actv_data[415:408]),

.io_dat_actv_5_52_valid(dat5_actv_pvld[52]),
.io_dat_actv_5_52_bits_nz(dat5_actv_nz[52]),
.io_dat_actv_5_52_bits_data(dat5_actv_data[423:416]),

.io_dat_actv_5_53_valid(dat5_actv_pvld[53]),
.io_dat_actv_5_53_bits_nz(dat5_actv_nz[53]),
.io_dat_actv_5_53_bits_data(dat5_actv_data[431:424]),

.io_dat_actv_5_54_valid(dat5_actv_pvld[54]),
.io_dat_actv_5_54_bits_nz(dat5_actv_nz[54]),
.io_dat_actv_5_54_bits_data(dat5_actv_data[439:432]),

.io_dat_actv_5_55_valid(dat5_actv_pvld[55]),
.io_dat_actv_5_55_bits_nz(dat5_actv_nz[55]),
.io_dat_actv_5_55_bits_data(dat5_actv_data[447:440]),

.io_dat_actv_5_56_valid(dat5_actv_pvld[56]),
.io_dat_actv_5_56_bits_nz(dat5_actv_nz[56]),
.io_dat_actv_5_56_bits_data(dat5_actv_data[455:448]),

.io_dat_actv_5_57_valid(dat5_actv_pvld[57]),
.io_dat_actv_5_57_bits_nz(dat5_actv_nz[57]),
.io_dat_actv_5_57_bits_data(dat5_actv_data[463:456]),

.io_dat_actv_5_58_valid(dat5_actv_pvld[58]),
.io_dat_actv_5_58_bits_nz(dat5_actv_nz[58]),
.io_dat_actv_5_58_bits_data(dat5_actv_data[471:464]),

.io_dat_actv_5_59_valid(dat5_actv_pvld[59]),
.io_dat_actv_5_59_bits_nz(dat5_actv_nz[59]),
.io_dat_actv_5_59_bits_data(dat5_actv_data[479:472]),

.io_dat_actv_5_60_valid(dat5_actv_pvld[60]),
.io_dat_actv_5_60_bits_nz(dat5_actv_nz[60]),
.io_dat_actv_5_60_bits_data(dat5_actv_data[487:480]),

.io_dat_actv_5_61_valid(dat5_actv_pvld[61]),
.io_dat_actv_5_61_bits_nz(dat5_actv_nz[61]),
.io_dat_actv_5_61_bits_data(dat5_actv_data[495:488]),

.io_dat_actv_5_62_valid(dat5_actv_pvld[62]),
.io_dat_actv_5_62_bits_nz(dat5_actv_nz[62]),
.io_dat_actv_5_62_bits_data(dat5_actv_data[503:496]),

.io_dat_actv_5_63_valid(dat5_actv_pvld[63]),
.io_dat_actv_5_63_bits_nz(dat5_actv_nz[63]),
.io_dat_actv_5_63_bits_data(dat5_actv_data[511:504]),

.io_dat_actv_6_0_valid(dat6_actv_pvld[0]),
.io_dat_actv_6_0_bits_nz(dat6_actv_nz[0]),
.io_dat_actv_6_0_bits_data(dat6_actv_data[7:0]),

.io_dat_actv_6_1_valid(dat6_actv_pvld[1]),
.io_dat_actv_6_1_bits_nz(dat6_actv_nz[1]),
.io_dat_actv_6_1_bits_data(dat6_actv_data[15:8]),

.io_dat_actv_6_2_valid(dat6_actv_pvld[2]),
.io_dat_actv_6_2_bits_nz(dat6_actv_nz[2]),
.io_dat_actv_6_2_bits_data(dat6_actv_data[23:16]),

.io_dat_actv_6_3_valid(dat6_actv_pvld[3]),
.io_dat_actv_6_3_bits_nz(dat6_actv_nz[3]),
.io_dat_actv_6_3_bits_data(dat6_actv_data[31:24]),

.io_dat_actv_6_4_valid(dat6_actv_pvld[4]),
.io_dat_actv_6_4_bits_nz(dat6_actv_nz[4]),
.io_dat_actv_6_4_bits_data(dat6_actv_data[39:32]),

.io_dat_actv_6_5_valid(dat6_actv_pvld[5]),
.io_dat_actv_6_5_bits_nz(dat6_actv_nz[5]),
.io_dat_actv_6_5_bits_data(dat6_actv_data[47:40]),

.io_dat_actv_6_6_valid(dat6_actv_pvld[6]),
.io_dat_actv_6_6_bits_nz(dat6_actv_nz[6]),
.io_dat_actv_6_6_bits_data(dat6_actv_data[55:48]),

.io_dat_actv_6_7_valid(dat6_actv_pvld[7]),
.io_dat_actv_6_7_bits_nz(dat6_actv_nz[7]),
.io_dat_actv_6_7_bits_data(dat6_actv_data[63:56]),

.io_dat_actv_6_8_valid(dat6_actv_pvld[8]),
.io_dat_actv_6_8_bits_nz(dat6_actv_nz[8]),
.io_dat_actv_6_8_bits_data(dat6_actv_data[71:64]),

.io_dat_actv_6_9_valid(dat6_actv_pvld[9]),
.io_dat_actv_6_9_bits_nz(dat6_actv_nz[9]),
.io_dat_actv_6_9_bits_data(dat6_actv_data[79:72]),

.io_dat_actv_6_10_valid(dat6_actv_pvld[10]),
.io_dat_actv_6_10_bits_nz(dat6_actv_nz[10]),
.io_dat_actv_6_10_bits_data(dat6_actv_data[87:80]),

.io_dat_actv_6_11_valid(dat6_actv_pvld[11]),
.io_dat_actv_6_11_bits_nz(dat6_actv_nz[11]),
.io_dat_actv_6_11_bits_data(dat6_actv_data[95:88]),

.io_dat_actv_6_12_valid(dat6_actv_pvld[12]),
.io_dat_actv_6_12_bits_nz(dat6_actv_nz[12]),
.io_dat_actv_6_12_bits_data(dat6_actv_data[103:96]),

.io_dat_actv_6_13_valid(dat6_actv_pvld[13]),
.io_dat_actv_6_13_bits_nz(dat6_actv_nz[13]),
.io_dat_actv_6_13_bits_data(dat6_actv_data[111:104]),

.io_dat_actv_6_14_valid(dat6_actv_pvld[14]),
.io_dat_actv_6_14_bits_nz(dat6_actv_nz[14]),
.io_dat_actv_6_14_bits_data(dat6_actv_data[119:112]),

.io_dat_actv_6_15_valid(dat6_actv_pvld[15]),
.io_dat_actv_6_15_bits_nz(dat6_actv_nz[15]),
.io_dat_actv_6_15_bits_data(dat6_actv_data[127:120]),

.io_dat_actv_6_16_valid(dat6_actv_pvld[16]),
.io_dat_actv_6_16_bits_nz(dat6_actv_nz[16]),
.io_dat_actv_6_16_bits_data(dat6_actv_data[135:128]),

.io_dat_actv_6_17_valid(dat6_actv_pvld[17]),
.io_dat_actv_6_17_bits_nz(dat6_actv_nz[17]),
.io_dat_actv_6_17_bits_data(dat6_actv_data[143:136]),

.io_dat_actv_6_18_valid(dat6_actv_pvld[18]),
.io_dat_actv_6_18_bits_nz(dat6_actv_nz[18]),
.io_dat_actv_6_18_bits_data(dat6_actv_data[151:144]),

.io_dat_actv_6_19_valid(dat6_actv_pvld[19]),
.io_dat_actv_6_19_bits_nz(dat6_actv_nz[19]),
.io_dat_actv_6_19_bits_data(dat6_actv_data[159:152]),

.io_dat_actv_6_20_valid(dat6_actv_pvld[20]),
.io_dat_actv_6_20_bits_nz(dat6_actv_nz[20]),
.io_dat_actv_6_20_bits_data(dat6_actv_data[167:160]),

.io_dat_actv_6_21_valid(dat6_actv_pvld[21]),
.io_dat_actv_6_21_bits_nz(dat6_actv_nz[21]),
.io_dat_actv_6_21_bits_data(dat6_actv_data[175:168]),

.io_dat_actv_6_22_valid(dat6_actv_pvld[22]),
.io_dat_actv_6_22_bits_nz(dat6_actv_nz[22]),
.io_dat_actv_6_22_bits_data(dat6_actv_data[183:176]),

.io_dat_actv_6_23_valid(dat6_actv_pvld[23]),
.io_dat_actv_6_23_bits_nz(dat6_actv_nz[23]),
.io_dat_actv_6_23_bits_data(dat6_actv_data[191:184]),

.io_dat_actv_6_24_valid(dat6_actv_pvld[24]),
.io_dat_actv_6_24_bits_nz(dat6_actv_nz[24]),
.io_dat_actv_6_24_bits_data(dat6_actv_data[199:192]),

.io_dat_actv_6_25_valid(dat6_actv_pvld[25]),
.io_dat_actv_6_25_bits_nz(dat6_actv_nz[25]),
.io_dat_actv_6_25_bits_data(dat6_actv_data[207:200]),

.io_dat_actv_6_26_valid(dat6_actv_pvld[26]),
.io_dat_actv_6_26_bits_nz(dat6_actv_nz[26]),
.io_dat_actv_6_26_bits_data(dat6_actv_data[215:208]),

.io_dat_actv_6_27_valid(dat6_actv_pvld[27]),
.io_dat_actv_6_27_bits_nz(dat6_actv_nz[27]),
.io_dat_actv_6_27_bits_data(dat6_actv_data[223:216]),

.io_dat_actv_6_28_valid(dat6_actv_pvld[28]),
.io_dat_actv_6_28_bits_nz(dat6_actv_nz[28]),
.io_dat_actv_6_28_bits_data(dat6_actv_data[231:224]),

.io_dat_actv_6_29_valid(dat6_actv_pvld[29]),
.io_dat_actv_6_29_bits_nz(dat6_actv_nz[29]),
.io_dat_actv_6_29_bits_data(dat6_actv_data[239:232]),

.io_dat_actv_6_30_valid(dat6_actv_pvld[30]),
.io_dat_actv_6_30_bits_nz(dat6_actv_nz[30]),
.io_dat_actv_6_30_bits_data(dat6_actv_data[247:240]),

.io_dat_actv_6_31_valid(dat6_actv_pvld[31]),
.io_dat_actv_6_31_bits_nz(dat6_actv_nz[31]),
.io_dat_actv_6_31_bits_data(dat6_actv_data[255:248]),

.io_dat_actv_6_32_valid(dat6_actv_pvld[32]),
.io_dat_actv_6_32_bits_nz(dat6_actv_nz[32]),
.io_dat_actv_6_32_bits_data(dat6_actv_data[263:256]),

.io_dat_actv_6_33_valid(dat6_actv_pvld[33]),
.io_dat_actv_6_33_bits_nz(dat6_actv_nz[33]),
.io_dat_actv_6_33_bits_data(dat6_actv_data[271:264]),

.io_dat_actv_6_34_valid(dat6_actv_pvld[34]),
.io_dat_actv_6_34_bits_nz(dat6_actv_nz[34]),
.io_dat_actv_6_34_bits_data(dat6_actv_data[279:272]),

.io_dat_actv_6_35_valid(dat6_actv_pvld[35]),
.io_dat_actv_6_35_bits_nz(dat6_actv_nz[35]),
.io_dat_actv_6_35_bits_data(dat6_actv_data[287:280]),

.io_dat_actv_6_36_valid(dat6_actv_pvld[36]),
.io_dat_actv_6_36_bits_nz(dat6_actv_nz[36]),
.io_dat_actv_6_36_bits_data(dat6_actv_data[295:288]),

.io_dat_actv_6_37_valid(dat6_actv_pvld[37]),
.io_dat_actv_6_37_bits_nz(dat6_actv_nz[37]),
.io_dat_actv_6_37_bits_data(dat6_actv_data[303:296]),

.io_dat_actv_6_38_valid(dat6_actv_pvld[38]),
.io_dat_actv_6_38_bits_nz(dat6_actv_nz[38]),
.io_dat_actv_6_38_bits_data(dat6_actv_data[311:304]),

.io_dat_actv_6_39_valid(dat6_actv_pvld[39]),
.io_dat_actv_6_39_bits_nz(dat6_actv_nz[39]),
.io_dat_actv_6_39_bits_data(dat6_actv_data[319:312]),

.io_dat_actv_6_40_valid(dat6_actv_pvld[40]),
.io_dat_actv_6_40_bits_nz(dat6_actv_nz[40]),
.io_dat_actv_6_40_bits_data(dat6_actv_data[327:320]),

.io_dat_actv_6_41_valid(dat6_actv_pvld[41]),
.io_dat_actv_6_41_bits_nz(dat6_actv_nz[41]),
.io_dat_actv_6_41_bits_data(dat6_actv_data[335:328]),

.io_dat_actv_6_42_valid(dat6_actv_pvld[42]),
.io_dat_actv_6_42_bits_nz(dat6_actv_nz[42]),
.io_dat_actv_6_42_bits_data(dat6_actv_data[343:336]),

.io_dat_actv_6_43_valid(dat6_actv_pvld[43]),
.io_dat_actv_6_43_bits_nz(dat6_actv_nz[43]),
.io_dat_actv_6_43_bits_data(dat6_actv_data[351:344]),

.io_dat_actv_6_44_valid(dat6_actv_pvld[44]),
.io_dat_actv_6_44_bits_nz(dat6_actv_nz[44]),
.io_dat_actv_6_44_bits_data(dat6_actv_data[359:352]),

.io_dat_actv_6_45_valid(dat6_actv_pvld[45]),
.io_dat_actv_6_45_bits_nz(dat6_actv_nz[45]),
.io_dat_actv_6_45_bits_data(dat6_actv_data[367:360]),

.io_dat_actv_6_46_valid(dat6_actv_pvld[46]),
.io_dat_actv_6_46_bits_nz(dat6_actv_nz[46]),
.io_dat_actv_6_46_bits_data(dat6_actv_data[375:368]),

.io_dat_actv_6_47_valid(dat6_actv_pvld[47]),
.io_dat_actv_6_47_bits_nz(dat6_actv_nz[47]),
.io_dat_actv_6_47_bits_data(dat6_actv_data[383:376]),

.io_dat_actv_6_48_valid(dat6_actv_pvld[48]),
.io_dat_actv_6_48_bits_nz(dat6_actv_nz[48]),
.io_dat_actv_6_48_bits_data(dat6_actv_data[391:384]),

.io_dat_actv_6_49_valid(dat6_actv_pvld[49]),
.io_dat_actv_6_49_bits_nz(dat6_actv_nz[49]),
.io_dat_actv_6_49_bits_data(dat6_actv_data[399:392]),

.io_dat_actv_6_50_valid(dat6_actv_pvld[50]),
.io_dat_actv_6_50_bits_nz(dat6_actv_nz[50]),
.io_dat_actv_6_50_bits_data(dat6_actv_data[407:400]),

.io_dat_actv_6_51_valid(dat6_actv_pvld[51]),
.io_dat_actv_6_51_bits_nz(dat6_actv_nz[51]),
.io_dat_actv_6_51_bits_data(dat6_actv_data[415:408]),

.io_dat_actv_6_52_valid(dat6_actv_pvld[52]),
.io_dat_actv_6_52_bits_nz(dat6_actv_nz[52]),
.io_dat_actv_6_52_bits_data(dat6_actv_data[423:416]),

.io_dat_actv_6_53_valid(dat6_actv_pvld[53]),
.io_dat_actv_6_53_bits_nz(dat6_actv_nz[53]),
.io_dat_actv_6_53_bits_data(dat6_actv_data[431:424]),

.io_dat_actv_6_54_valid(dat6_actv_pvld[54]),
.io_dat_actv_6_54_bits_nz(dat6_actv_nz[54]),
.io_dat_actv_6_54_bits_data(dat6_actv_data[439:432]),

.io_dat_actv_6_55_valid(dat6_actv_pvld[55]),
.io_dat_actv_6_55_bits_nz(dat6_actv_nz[55]),
.io_dat_actv_6_55_bits_data(dat6_actv_data[447:440]),

.io_dat_actv_6_56_valid(dat6_actv_pvld[56]),
.io_dat_actv_6_56_bits_nz(dat6_actv_nz[56]),
.io_dat_actv_6_56_bits_data(dat6_actv_data[455:448]),

.io_dat_actv_6_57_valid(dat6_actv_pvld[57]),
.io_dat_actv_6_57_bits_nz(dat6_actv_nz[57]),
.io_dat_actv_6_57_bits_data(dat6_actv_data[463:456]),

.io_dat_actv_6_58_valid(dat6_actv_pvld[58]),
.io_dat_actv_6_58_bits_nz(dat6_actv_nz[58]),
.io_dat_actv_6_58_bits_data(dat6_actv_data[471:464]),

.io_dat_actv_6_59_valid(dat6_actv_pvld[59]),
.io_dat_actv_6_59_bits_nz(dat6_actv_nz[59]),
.io_dat_actv_6_59_bits_data(dat6_actv_data[479:472]),

.io_dat_actv_6_60_valid(dat6_actv_pvld[60]),
.io_dat_actv_6_60_bits_nz(dat6_actv_nz[60]),
.io_dat_actv_6_60_bits_data(dat6_actv_data[487:480]),

.io_dat_actv_6_61_valid(dat6_actv_pvld[61]),
.io_dat_actv_6_61_bits_nz(dat6_actv_nz[61]),
.io_dat_actv_6_61_bits_data(dat6_actv_data[495:488]),

.io_dat_actv_6_62_valid(dat6_actv_pvld[62]),
.io_dat_actv_6_62_bits_nz(dat6_actv_nz[62]),
.io_dat_actv_6_62_bits_data(dat6_actv_data[503:496]),

.io_dat_actv_6_63_valid(dat6_actv_pvld[63]),
.io_dat_actv_6_63_bits_nz(dat6_actv_nz[63]),
.io_dat_actv_6_63_bits_data(dat6_actv_data[511:504]),

.io_dat_actv_7_0_valid(dat7_actv_pvld[0]),
.io_dat_actv_7_0_bits_nz(dat7_actv_nz[0]),
.io_dat_actv_7_0_bits_data(dat7_actv_data[7:0]),

.io_dat_actv_7_1_valid(dat7_actv_pvld[1]),
.io_dat_actv_7_1_bits_nz(dat7_actv_nz[1]),
.io_dat_actv_7_1_bits_data(dat7_actv_data[15:8]),

.io_dat_actv_7_2_valid(dat7_actv_pvld[2]),
.io_dat_actv_7_2_bits_nz(dat7_actv_nz[2]),
.io_dat_actv_7_2_bits_data(dat7_actv_data[23:16]),

.io_dat_actv_7_3_valid(dat7_actv_pvld[3]),
.io_dat_actv_7_3_bits_nz(dat7_actv_nz[3]),
.io_dat_actv_7_3_bits_data(dat7_actv_data[31:24]),

.io_dat_actv_7_4_valid(dat7_actv_pvld[4]),
.io_dat_actv_7_4_bits_nz(dat7_actv_nz[4]),
.io_dat_actv_7_4_bits_data(dat7_actv_data[39:32]),

.io_dat_actv_7_5_valid(dat7_actv_pvld[5]),
.io_dat_actv_7_5_bits_nz(dat7_actv_nz[5]),
.io_dat_actv_7_5_bits_data(dat7_actv_data[47:40]),

.io_dat_actv_7_6_valid(dat7_actv_pvld[6]),
.io_dat_actv_7_6_bits_nz(dat7_actv_nz[6]),
.io_dat_actv_7_6_bits_data(dat7_actv_data[55:48]),

.io_dat_actv_7_7_valid(dat7_actv_pvld[7]),
.io_dat_actv_7_7_bits_nz(dat7_actv_nz[7]),
.io_dat_actv_7_7_bits_data(dat7_actv_data[63:56]),

.io_dat_actv_7_8_valid(dat7_actv_pvld[8]),
.io_dat_actv_7_8_bits_nz(dat7_actv_nz[8]),
.io_dat_actv_7_8_bits_data(dat7_actv_data[71:64]),

.io_dat_actv_7_9_valid(dat7_actv_pvld[9]),
.io_dat_actv_7_9_bits_nz(dat7_actv_nz[9]),
.io_dat_actv_7_9_bits_data(dat7_actv_data[79:72]),

.io_dat_actv_7_10_valid(dat7_actv_pvld[10]),
.io_dat_actv_7_10_bits_nz(dat7_actv_nz[10]),
.io_dat_actv_7_10_bits_data(dat7_actv_data[87:80]),

.io_dat_actv_7_11_valid(dat7_actv_pvld[11]),
.io_dat_actv_7_11_bits_nz(dat7_actv_nz[11]),
.io_dat_actv_7_11_bits_data(dat7_actv_data[95:88]),

.io_dat_actv_7_12_valid(dat7_actv_pvld[12]),
.io_dat_actv_7_12_bits_nz(dat7_actv_nz[12]),
.io_dat_actv_7_12_bits_data(dat7_actv_data[103:96]),

.io_dat_actv_7_13_valid(dat7_actv_pvld[13]),
.io_dat_actv_7_13_bits_nz(dat7_actv_nz[13]),
.io_dat_actv_7_13_bits_data(dat7_actv_data[111:104]),

.io_dat_actv_7_14_valid(dat7_actv_pvld[14]),
.io_dat_actv_7_14_bits_nz(dat7_actv_nz[14]),
.io_dat_actv_7_14_bits_data(dat7_actv_data[119:112]),

.io_dat_actv_7_15_valid(dat7_actv_pvld[15]),
.io_dat_actv_7_15_bits_nz(dat7_actv_nz[15]),
.io_dat_actv_7_15_bits_data(dat7_actv_data[127:120]),

.io_dat_actv_7_16_valid(dat7_actv_pvld[16]),
.io_dat_actv_7_16_bits_nz(dat7_actv_nz[16]),
.io_dat_actv_7_16_bits_data(dat7_actv_data[135:128]),

.io_dat_actv_7_17_valid(dat7_actv_pvld[17]),
.io_dat_actv_7_17_bits_nz(dat7_actv_nz[17]),
.io_dat_actv_7_17_bits_data(dat7_actv_data[143:136]),

.io_dat_actv_7_18_valid(dat7_actv_pvld[18]),
.io_dat_actv_7_18_bits_nz(dat7_actv_nz[18]),
.io_dat_actv_7_18_bits_data(dat7_actv_data[151:144]),

.io_dat_actv_7_19_valid(dat7_actv_pvld[19]),
.io_dat_actv_7_19_bits_nz(dat7_actv_nz[19]),
.io_dat_actv_7_19_bits_data(dat7_actv_data[159:152]),

.io_dat_actv_7_20_valid(dat7_actv_pvld[20]),
.io_dat_actv_7_20_bits_nz(dat7_actv_nz[20]),
.io_dat_actv_7_20_bits_data(dat7_actv_data[167:160]),

.io_dat_actv_7_21_valid(dat7_actv_pvld[21]),
.io_dat_actv_7_21_bits_nz(dat7_actv_nz[21]),
.io_dat_actv_7_21_bits_data(dat7_actv_data[175:168]),

.io_dat_actv_7_22_valid(dat7_actv_pvld[22]),
.io_dat_actv_7_22_bits_nz(dat7_actv_nz[22]),
.io_dat_actv_7_22_bits_data(dat7_actv_data[183:176]),

.io_dat_actv_7_23_valid(dat7_actv_pvld[23]),
.io_dat_actv_7_23_bits_nz(dat7_actv_nz[23]),
.io_dat_actv_7_23_bits_data(dat7_actv_data[191:184]),

.io_dat_actv_7_24_valid(dat7_actv_pvld[24]),
.io_dat_actv_7_24_bits_nz(dat7_actv_nz[24]),
.io_dat_actv_7_24_bits_data(dat7_actv_data[199:192]),

.io_dat_actv_7_25_valid(dat7_actv_pvld[25]),
.io_dat_actv_7_25_bits_nz(dat7_actv_nz[25]),
.io_dat_actv_7_25_bits_data(dat7_actv_data[207:200]),

.io_dat_actv_7_26_valid(dat7_actv_pvld[26]),
.io_dat_actv_7_26_bits_nz(dat7_actv_nz[26]),
.io_dat_actv_7_26_bits_data(dat7_actv_data[215:208]),

.io_dat_actv_7_27_valid(dat7_actv_pvld[27]),
.io_dat_actv_7_27_bits_nz(dat7_actv_nz[27]),
.io_dat_actv_7_27_bits_data(dat7_actv_data[223:216]),

.io_dat_actv_7_28_valid(dat7_actv_pvld[28]),
.io_dat_actv_7_28_bits_nz(dat7_actv_nz[28]),
.io_dat_actv_7_28_bits_data(dat7_actv_data[231:224]),

.io_dat_actv_7_29_valid(dat7_actv_pvld[29]),
.io_dat_actv_7_29_bits_nz(dat7_actv_nz[29]),
.io_dat_actv_7_29_bits_data(dat7_actv_data[239:232]),

.io_dat_actv_7_30_valid(dat7_actv_pvld[30]),
.io_dat_actv_7_30_bits_nz(dat7_actv_nz[30]),
.io_dat_actv_7_30_bits_data(dat7_actv_data[247:240]),

.io_dat_actv_7_31_valid(dat7_actv_pvld[31]),
.io_dat_actv_7_31_bits_nz(dat7_actv_nz[31]),
.io_dat_actv_7_31_bits_data(dat7_actv_data[255:248]),

.io_dat_actv_7_32_valid(dat7_actv_pvld[32]),
.io_dat_actv_7_32_bits_nz(dat7_actv_nz[32]),
.io_dat_actv_7_32_bits_data(dat7_actv_data[263:256]),

.io_dat_actv_7_33_valid(dat7_actv_pvld[33]),
.io_dat_actv_7_33_bits_nz(dat7_actv_nz[33]),
.io_dat_actv_7_33_bits_data(dat7_actv_data[271:264]),

.io_dat_actv_7_34_valid(dat7_actv_pvld[34]),
.io_dat_actv_7_34_bits_nz(dat7_actv_nz[34]),
.io_dat_actv_7_34_bits_data(dat7_actv_data[279:272]),

.io_dat_actv_7_35_valid(dat7_actv_pvld[35]),
.io_dat_actv_7_35_bits_nz(dat7_actv_nz[35]),
.io_dat_actv_7_35_bits_data(dat7_actv_data[287:280]),

.io_dat_actv_7_36_valid(dat7_actv_pvld[36]),
.io_dat_actv_7_36_bits_nz(dat7_actv_nz[36]),
.io_dat_actv_7_36_bits_data(dat7_actv_data[295:288]),

.io_dat_actv_7_37_valid(dat7_actv_pvld[37]),
.io_dat_actv_7_37_bits_nz(dat7_actv_nz[37]),
.io_dat_actv_7_37_bits_data(dat7_actv_data[303:296]),

.io_dat_actv_7_38_valid(dat7_actv_pvld[38]),
.io_dat_actv_7_38_bits_nz(dat7_actv_nz[38]),
.io_dat_actv_7_38_bits_data(dat7_actv_data[311:304]),

.io_dat_actv_7_39_valid(dat7_actv_pvld[39]),
.io_dat_actv_7_39_bits_nz(dat7_actv_nz[39]),
.io_dat_actv_7_39_bits_data(dat7_actv_data[319:312]),

.io_dat_actv_7_40_valid(dat7_actv_pvld[40]),
.io_dat_actv_7_40_bits_nz(dat7_actv_nz[40]),
.io_dat_actv_7_40_bits_data(dat7_actv_data[327:320]),

.io_dat_actv_7_41_valid(dat7_actv_pvld[41]),
.io_dat_actv_7_41_bits_nz(dat7_actv_nz[41]),
.io_dat_actv_7_41_bits_data(dat7_actv_data[335:328]),

.io_dat_actv_7_42_valid(dat7_actv_pvld[42]),
.io_dat_actv_7_42_bits_nz(dat7_actv_nz[42]),
.io_dat_actv_7_42_bits_data(dat7_actv_data[343:336]),

.io_dat_actv_7_43_valid(dat7_actv_pvld[43]),
.io_dat_actv_7_43_bits_nz(dat7_actv_nz[43]),
.io_dat_actv_7_43_bits_data(dat7_actv_data[351:344]),

.io_dat_actv_7_44_valid(dat7_actv_pvld[44]),
.io_dat_actv_7_44_bits_nz(dat7_actv_nz[44]),
.io_dat_actv_7_44_bits_data(dat7_actv_data[359:352]),

.io_dat_actv_7_45_valid(dat7_actv_pvld[45]),
.io_dat_actv_7_45_bits_nz(dat7_actv_nz[45]),
.io_dat_actv_7_45_bits_data(dat7_actv_data[367:360]),

.io_dat_actv_7_46_valid(dat7_actv_pvld[46]),
.io_dat_actv_7_46_bits_nz(dat7_actv_nz[46]),
.io_dat_actv_7_46_bits_data(dat7_actv_data[375:368]),

.io_dat_actv_7_47_valid(dat7_actv_pvld[47]),
.io_dat_actv_7_47_bits_nz(dat7_actv_nz[47]),
.io_dat_actv_7_47_bits_data(dat7_actv_data[383:376]),

.io_dat_actv_7_48_valid(dat7_actv_pvld[48]),
.io_dat_actv_7_48_bits_nz(dat7_actv_nz[48]),
.io_dat_actv_7_48_bits_data(dat7_actv_data[391:384]),

.io_dat_actv_7_49_valid(dat7_actv_pvld[49]),
.io_dat_actv_7_49_bits_nz(dat7_actv_nz[49]),
.io_dat_actv_7_49_bits_data(dat7_actv_data[399:392]),

.io_dat_actv_7_50_valid(dat7_actv_pvld[50]),
.io_dat_actv_7_50_bits_nz(dat7_actv_nz[50]),
.io_dat_actv_7_50_bits_data(dat7_actv_data[407:400]),

.io_dat_actv_7_51_valid(dat7_actv_pvld[51]),
.io_dat_actv_7_51_bits_nz(dat7_actv_nz[51]),
.io_dat_actv_7_51_bits_data(dat7_actv_data[415:408]),

.io_dat_actv_7_52_valid(dat7_actv_pvld[52]),
.io_dat_actv_7_52_bits_nz(dat7_actv_nz[52]),
.io_dat_actv_7_52_bits_data(dat7_actv_data[423:416]),

.io_dat_actv_7_53_valid(dat7_actv_pvld[53]),
.io_dat_actv_7_53_bits_nz(dat7_actv_nz[53]),
.io_dat_actv_7_53_bits_data(dat7_actv_data[431:424]),

.io_dat_actv_7_54_valid(dat7_actv_pvld[54]),
.io_dat_actv_7_54_bits_nz(dat7_actv_nz[54]),
.io_dat_actv_7_54_bits_data(dat7_actv_data[439:432]),

.io_dat_actv_7_55_valid(dat7_actv_pvld[55]),
.io_dat_actv_7_55_bits_nz(dat7_actv_nz[55]),
.io_dat_actv_7_55_bits_data(dat7_actv_data[447:440]),

.io_dat_actv_7_56_valid(dat7_actv_pvld[56]),
.io_dat_actv_7_56_bits_nz(dat7_actv_nz[56]),
.io_dat_actv_7_56_bits_data(dat7_actv_data[455:448]),

.io_dat_actv_7_57_valid(dat7_actv_pvld[57]),
.io_dat_actv_7_57_bits_nz(dat7_actv_nz[57]),
.io_dat_actv_7_57_bits_data(dat7_actv_data[463:456]),

.io_dat_actv_7_58_valid(dat7_actv_pvld[58]),
.io_dat_actv_7_58_bits_nz(dat7_actv_nz[58]),
.io_dat_actv_7_58_bits_data(dat7_actv_data[471:464]),

.io_dat_actv_7_59_valid(dat7_actv_pvld[59]),
.io_dat_actv_7_59_bits_nz(dat7_actv_nz[59]),
.io_dat_actv_7_59_bits_data(dat7_actv_data[479:472]),

.io_dat_actv_7_60_valid(dat7_actv_pvld[60]),
.io_dat_actv_7_60_bits_nz(dat7_actv_nz[60]),
.io_dat_actv_7_60_bits_data(dat7_actv_data[487:480]),

.io_dat_actv_7_61_valid(dat7_actv_pvld[61]),
.io_dat_actv_7_61_bits_nz(dat7_actv_nz[61]),
.io_dat_actv_7_61_bits_data(dat7_actv_data[495:488]),

.io_dat_actv_7_62_valid(dat7_actv_pvld[62]),
.io_dat_actv_7_62_bits_nz(dat7_actv_nz[62]),
.io_dat_actv_7_62_bits_data(dat7_actv_data[503:496]),

.io_dat_actv_7_63_valid(dat7_actv_pvld[63]),
.io_dat_actv_7_63_bits_nz(dat7_actv_nz[63]),
.io_dat_actv_7_63_bits_data(dat7_actv_data[511:504]),

.io_dat_actv_8_0_valid(dat8_actv_pvld[0]),
.io_dat_actv_8_0_bits_nz(dat8_actv_nz[0]),
.io_dat_actv_8_0_bits_data(dat8_actv_data[7:0]),

.io_dat_actv_8_1_valid(dat8_actv_pvld[1]),
.io_dat_actv_8_1_bits_nz(dat8_actv_nz[1]),
.io_dat_actv_8_1_bits_data(dat8_actv_data[15:8]),

.io_dat_actv_8_2_valid(dat8_actv_pvld[2]),
.io_dat_actv_8_2_bits_nz(dat8_actv_nz[2]),
.io_dat_actv_8_2_bits_data(dat8_actv_data[23:16]),

.io_dat_actv_8_3_valid(dat8_actv_pvld[3]),
.io_dat_actv_8_3_bits_nz(dat8_actv_nz[3]),
.io_dat_actv_8_3_bits_data(dat8_actv_data[31:24]),

.io_dat_actv_8_4_valid(dat8_actv_pvld[4]),
.io_dat_actv_8_4_bits_nz(dat8_actv_nz[4]),
.io_dat_actv_8_4_bits_data(dat8_actv_data[39:32]),

.io_dat_actv_8_5_valid(dat8_actv_pvld[5]),
.io_dat_actv_8_5_bits_nz(dat8_actv_nz[5]),
.io_dat_actv_8_5_bits_data(dat8_actv_data[47:40]),

.io_dat_actv_8_6_valid(dat8_actv_pvld[6]),
.io_dat_actv_8_6_bits_nz(dat8_actv_nz[6]),
.io_dat_actv_8_6_bits_data(dat8_actv_data[55:48]),

.io_dat_actv_8_7_valid(dat8_actv_pvld[7]),
.io_dat_actv_8_7_bits_nz(dat8_actv_nz[7]),
.io_dat_actv_8_7_bits_data(dat8_actv_data[63:56]),

.io_dat_actv_8_8_valid(dat8_actv_pvld[8]),
.io_dat_actv_8_8_bits_nz(dat8_actv_nz[8]),
.io_dat_actv_8_8_bits_data(dat8_actv_data[71:64]),

.io_dat_actv_8_9_valid(dat8_actv_pvld[9]),
.io_dat_actv_8_9_bits_nz(dat8_actv_nz[9]),
.io_dat_actv_8_9_bits_data(dat8_actv_data[79:72]),

.io_dat_actv_8_10_valid(dat8_actv_pvld[10]),
.io_dat_actv_8_10_bits_nz(dat8_actv_nz[10]),
.io_dat_actv_8_10_bits_data(dat8_actv_data[87:80]),

.io_dat_actv_8_11_valid(dat8_actv_pvld[11]),
.io_dat_actv_8_11_bits_nz(dat8_actv_nz[11]),
.io_dat_actv_8_11_bits_data(dat8_actv_data[95:88]),

.io_dat_actv_8_12_valid(dat8_actv_pvld[12]),
.io_dat_actv_8_12_bits_nz(dat8_actv_nz[12]),
.io_dat_actv_8_12_bits_data(dat8_actv_data[103:96]),

.io_dat_actv_8_13_valid(dat8_actv_pvld[13]),
.io_dat_actv_8_13_bits_nz(dat8_actv_nz[13]),
.io_dat_actv_8_13_bits_data(dat8_actv_data[111:104]),

.io_dat_actv_8_14_valid(dat8_actv_pvld[14]),
.io_dat_actv_8_14_bits_nz(dat8_actv_nz[14]),
.io_dat_actv_8_14_bits_data(dat8_actv_data[119:112]),

.io_dat_actv_8_15_valid(dat8_actv_pvld[15]),
.io_dat_actv_8_15_bits_nz(dat8_actv_nz[15]),
.io_dat_actv_8_15_bits_data(dat8_actv_data[127:120]),

.io_dat_actv_8_16_valid(dat8_actv_pvld[16]),
.io_dat_actv_8_16_bits_nz(dat8_actv_nz[16]),
.io_dat_actv_8_16_bits_data(dat8_actv_data[135:128]),

.io_dat_actv_8_17_valid(dat8_actv_pvld[17]),
.io_dat_actv_8_17_bits_nz(dat8_actv_nz[17]),
.io_dat_actv_8_17_bits_data(dat8_actv_data[143:136]),

.io_dat_actv_8_18_valid(dat8_actv_pvld[18]),
.io_dat_actv_8_18_bits_nz(dat8_actv_nz[18]),
.io_dat_actv_8_18_bits_data(dat8_actv_data[151:144]),

.io_dat_actv_8_19_valid(dat8_actv_pvld[19]),
.io_dat_actv_8_19_bits_nz(dat8_actv_nz[19]),
.io_dat_actv_8_19_bits_data(dat8_actv_data[159:152]),

.io_dat_actv_8_20_valid(dat8_actv_pvld[20]),
.io_dat_actv_8_20_bits_nz(dat8_actv_nz[20]),
.io_dat_actv_8_20_bits_data(dat8_actv_data[167:160]),

.io_dat_actv_8_21_valid(dat8_actv_pvld[21]),
.io_dat_actv_8_21_bits_nz(dat8_actv_nz[21]),
.io_dat_actv_8_21_bits_data(dat8_actv_data[175:168]),

.io_dat_actv_8_22_valid(dat8_actv_pvld[22]),
.io_dat_actv_8_22_bits_nz(dat8_actv_nz[22]),
.io_dat_actv_8_22_bits_data(dat8_actv_data[183:176]),

.io_dat_actv_8_23_valid(dat8_actv_pvld[23]),
.io_dat_actv_8_23_bits_nz(dat8_actv_nz[23]),
.io_dat_actv_8_23_bits_data(dat8_actv_data[191:184]),

.io_dat_actv_8_24_valid(dat8_actv_pvld[24]),
.io_dat_actv_8_24_bits_nz(dat8_actv_nz[24]),
.io_dat_actv_8_24_bits_data(dat8_actv_data[199:192]),

.io_dat_actv_8_25_valid(dat8_actv_pvld[25]),
.io_dat_actv_8_25_bits_nz(dat8_actv_nz[25]),
.io_dat_actv_8_25_bits_data(dat8_actv_data[207:200]),

.io_dat_actv_8_26_valid(dat8_actv_pvld[26]),
.io_dat_actv_8_26_bits_nz(dat8_actv_nz[26]),
.io_dat_actv_8_26_bits_data(dat8_actv_data[215:208]),

.io_dat_actv_8_27_valid(dat8_actv_pvld[27]),
.io_dat_actv_8_27_bits_nz(dat8_actv_nz[27]),
.io_dat_actv_8_27_bits_data(dat8_actv_data[223:216]),

.io_dat_actv_8_28_valid(dat8_actv_pvld[28]),
.io_dat_actv_8_28_bits_nz(dat8_actv_nz[28]),
.io_dat_actv_8_28_bits_data(dat8_actv_data[231:224]),

.io_dat_actv_8_29_valid(dat8_actv_pvld[29]),
.io_dat_actv_8_29_bits_nz(dat8_actv_nz[29]),
.io_dat_actv_8_29_bits_data(dat8_actv_data[239:232]),

.io_dat_actv_8_30_valid(dat8_actv_pvld[30]),
.io_dat_actv_8_30_bits_nz(dat8_actv_nz[30]),
.io_dat_actv_8_30_bits_data(dat8_actv_data[247:240]),

.io_dat_actv_8_31_valid(dat8_actv_pvld[31]),
.io_dat_actv_8_31_bits_nz(dat8_actv_nz[31]),
.io_dat_actv_8_31_bits_data(dat8_actv_data[255:248]),

.io_dat_actv_8_32_valid(dat8_actv_pvld[32]),
.io_dat_actv_8_32_bits_nz(dat8_actv_nz[32]),
.io_dat_actv_8_32_bits_data(dat8_actv_data[263:256]),

.io_dat_actv_8_33_valid(dat8_actv_pvld[33]),
.io_dat_actv_8_33_bits_nz(dat8_actv_nz[33]),
.io_dat_actv_8_33_bits_data(dat8_actv_data[271:264]),

.io_dat_actv_8_34_valid(dat8_actv_pvld[34]),
.io_dat_actv_8_34_bits_nz(dat8_actv_nz[34]),
.io_dat_actv_8_34_bits_data(dat8_actv_data[279:272]),

.io_dat_actv_8_35_valid(dat8_actv_pvld[35]),
.io_dat_actv_8_35_bits_nz(dat8_actv_nz[35]),
.io_dat_actv_8_35_bits_data(dat8_actv_data[287:280]),

.io_dat_actv_8_36_valid(dat8_actv_pvld[36]),
.io_dat_actv_8_36_bits_nz(dat8_actv_nz[36]),
.io_dat_actv_8_36_bits_data(dat8_actv_data[295:288]),

.io_dat_actv_8_37_valid(dat8_actv_pvld[37]),
.io_dat_actv_8_37_bits_nz(dat8_actv_nz[37]),
.io_dat_actv_8_37_bits_data(dat8_actv_data[303:296]),

.io_dat_actv_8_38_valid(dat8_actv_pvld[38]),
.io_dat_actv_8_38_bits_nz(dat8_actv_nz[38]),
.io_dat_actv_8_38_bits_data(dat8_actv_data[311:304]),

.io_dat_actv_8_39_valid(dat8_actv_pvld[39]),
.io_dat_actv_8_39_bits_nz(dat8_actv_nz[39]),
.io_dat_actv_8_39_bits_data(dat8_actv_data[319:312]),

.io_dat_actv_8_40_valid(dat8_actv_pvld[40]),
.io_dat_actv_8_40_bits_nz(dat8_actv_nz[40]),
.io_dat_actv_8_40_bits_data(dat8_actv_data[327:320]),

.io_dat_actv_8_41_valid(dat8_actv_pvld[41]),
.io_dat_actv_8_41_bits_nz(dat8_actv_nz[41]),
.io_dat_actv_8_41_bits_data(dat8_actv_data[335:328]),

.io_dat_actv_8_42_valid(dat8_actv_pvld[42]),
.io_dat_actv_8_42_bits_nz(dat8_actv_nz[42]),
.io_dat_actv_8_42_bits_data(dat8_actv_data[343:336]),

.io_dat_actv_8_43_valid(dat8_actv_pvld[43]),
.io_dat_actv_8_43_bits_nz(dat8_actv_nz[43]),
.io_dat_actv_8_43_bits_data(dat8_actv_data[351:344]),

.io_dat_actv_8_44_valid(dat8_actv_pvld[44]),
.io_dat_actv_8_44_bits_nz(dat8_actv_nz[44]),
.io_dat_actv_8_44_bits_data(dat8_actv_data[359:352]),

.io_dat_actv_8_45_valid(dat8_actv_pvld[45]),
.io_dat_actv_8_45_bits_nz(dat8_actv_nz[45]),
.io_dat_actv_8_45_bits_data(dat8_actv_data[367:360]),

.io_dat_actv_8_46_valid(dat8_actv_pvld[46]),
.io_dat_actv_8_46_bits_nz(dat8_actv_nz[46]),
.io_dat_actv_8_46_bits_data(dat8_actv_data[375:368]),

.io_dat_actv_8_47_valid(dat8_actv_pvld[47]),
.io_dat_actv_8_47_bits_nz(dat8_actv_nz[47]),
.io_dat_actv_8_47_bits_data(dat8_actv_data[383:376]),

.io_dat_actv_8_48_valid(dat8_actv_pvld[48]),
.io_dat_actv_8_48_bits_nz(dat8_actv_nz[48]),
.io_dat_actv_8_48_bits_data(dat8_actv_data[391:384]),

.io_dat_actv_8_49_valid(dat8_actv_pvld[49]),
.io_dat_actv_8_49_bits_nz(dat8_actv_nz[49]),
.io_dat_actv_8_49_bits_data(dat8_actv_data[399:392]),

.io_dat_actv_8_50_valid(dat8_actv_pvld[50]),
.io_dat_actv_8_50_bits_nz(dat8_actv_nz[50]),
.io_dat_actv_8_50_bits_data(dat8_actv_data[407:400]),

.io_dat_actv_8_51_valid(dat8_actv_pvld[51]),
.io_dat_actv_8_51_bits_nz(dat8_actv_nz[51]),
.io_dat_actv_8_51_bits_data(dat8_actv_data[415:408]),

.io_dat_actv_8_52_valid(dat8_actv_pvld[52]),
.io_dat_actv_8_52_bits_nz(dat8_actv_nz[52]),
.io_dat_actv_8_52_bits_data(dat8_actv_data[423:416]),

.io_dat_actv_8_53_valid(dat8_actv_pvld[53]),
.io_dat_actv_8_53_bits_nz(dat8_actv_nz[53]),
.io_dat_actv_8_53_bits_data(dat8_actv_data[431:424]),

.io_dat_actv_8_54_valid(dat8_actv_pvld[54]),
.io_dat_actv_8_54_bits_nz(dat8_actv_nz[54]),
.io_dat_actv_8_54_bits_data(dat8_actv_data[439:432]),

.io_dat_actv_8_55_valid(dat8_actv_pvld[55]),
.io_dat_actv_8_55_bits_nz(dat8_actv_nz[55]),
.io_dat_actv_8_55_bits_data(dat8_actv_data[447:440]),

.io_dat_actv_8_56_valid(dat8_actv_pvld[56]),
.io_dat_actv_8_56_bits_nz(dat8_actv_nz[56]),
.io_dat_actv_8_56_bits_data(dat8_actv_data[455:448]),

.io_dat_actv_8_57_valid(dat8_actv_pvld[57]),
.io_dat_actv_8_57_bits_nz(dat8_actv_nz[57]),
.io_dat_actv_8_57_bits_data(dat8_actv_data[463:456]),

.io_dat_actv_8_58_valid(dat8_actv_pvld[58]),
.io_dat_actv_8_58_bits_nz(dat8_actv_nz[58]),
.io_dat_actv_8_58_bits_data(dat8_actv_data[471:464]),

.io_dat_actv_8_59_valid(dat8_actv_pvld[59]),
.io_dat_actv_8_59_bits_nz(dat8_actv_nz[59]),
.io_dat_actv_8_59_bits_data(dat8_actv_data[479:472]),

.io_dat_actv_8_60_valid(dat8_actv_pvld[60]),
.io_dat_actv_8_60_bits_nz(dat8_actv_nz[60]),
.io_dat_actv_8_60_bits_data(dat8_actv_data[487:480]),

.io_dat_actv_8_61_valid(dat8_actv_pvld[61]),
.io_dat_actv_8_61_bits_nz(dat8_actv_nz[61]),
.io_dat_actv_8_61_bits_data(dat8_actv_data[495:488]),

.io_dat_actv_8_62_valid(dat8_actv_pvld[62]),
.io_dat_actv_8_62_bits_nz(dat8_actv_nz[62]),
.io_dat_actv_8_62_bits_data(dat8_actv_data[503:496]),

.io_dat_actv_8_63_valid(dat8_actv_pvld[63]),
.io_dat_actv_8_63_bits_nz(dat8_actv_nz[63]),
.io_dat_actv_8_63_bits_data(dat8_actv_data[511:504]),

.io_dat_actv_9_0_valid(dat9_actv_pvld[0]),
.io_dat_actv_9_0_bits_nz(dat9_actv_nz[0]),
.io_dat_actv_9_0_bits_data(dat9_actv_data[7:0]),

.io_dat_actv_9_1_valid(dat9_actv_pvld[1]),
.io_dat_actv_9_1_bits_nz(dat9_actv_nz[1]),
.io_dat_actv_9_1_bits_data(dat9_actv_data[15:8]),

.io_dat_actv_9_2_valid(dat9_actv_pvld[2]),
.io_dat_actv_9_2_bits_nz(dat9_actv_nz[2]),
.io_dat_actv_9_2_bits_data(dat9_actv_data[23:16]),

.io_dat_actv_9_3_valid(dat9_actv_pvld[3]),
.io_dat_actv_9_3_bits_nz(dat9_actv_nz[3]),
.io_dat_actv_9_3_bits_data(dat9_actv_data[31:24]),

.io_dat_actv_9_4_valid(dat9_actv_pvld[4]),
.io_dat_actv_9_4_bits_nz(dat9_actv_nz[4]),
.io_dat_actv_9_4_bits_data(dat9_actv_data[39:32]),

.io_dat_actv_9_5_valid(dat9_actv_pvld[5]),
.io_dat_actv_9_5_bits_nz(dat9_actv_nz[5]),
.io_dat_actv_9_5_bits_data(dat9_actv_data[47:40]),

.io_dat_actv_9_6_valid(dat9_actv_pvld[6]),
.io_dat_actv_9_6_bits_nz(dat9_actv_nz[6]),
.io_dat_actv_9_6_bits_data(dat9_actv_data[55:48]),

.io_dat_actv_9_7_valid(dat9_actv_pvld[7]),
.io_dat_actv_9_7_bits_nz(dat9_actv_nz[7]),
.io_dat_actv_9_7_bits_data(dat9_actv_data[63:56]),

.io_dat_actv_9_8_valid(dat9_actv_pvld[8]),
.io_dat_actv_9_8_bits_nz(dat9_actv_nz[8]),
.io_dat_actv_9_8_bits_data(dat9_actv_data[71:64]),

.io_dat_actv_9_9_valid(dat9_actv_pvld[9]),
.io_dat_actv_9_9_bits_nz(dat9_actv_nz[9]),
.io_dat_actv_9_9_bits_data(dat9_actv_data[79:72]),

.io_dat_actv_9_10_valid(dat9_actv_pvld[10]),
.io_dat_actv_9_10_bits_nz(dat9_actv_nz[10]),
.io_dat_actv_9_10_bits_data(dat9_actv_data[87:80]),

.io_dat_actv_9_11_valid(dat9_actv_pvld[11]),
.io_dat_actv_9_11_bits_nz(dat9_actv_nz[11]),
.io_dat_actv_9_11_bits_data(dat9_actv_data[95:88]),

.io_dat_actv_9_12_valid(dat9_actv_pvld[12]),
.io_dat_actv_9_12_bits_nz(dat9_actv_nz[12]),
.io_dat_actv_9_12_bits_data(dat9_actv_data[103:96]),

.io_dat_actv_9_13_valid(dat9_actv_pvld[13]),
.io_dat_actv_9_13_bits_nz(dat9_actv_nz[13]),
.io_dat_actv_9_13_bits_data(dat9_actv_data[111:104]),

.io_dat_actv_9_14_valid(dat9_actv_pvld[14]),
.io_dat_actv_9_14_bits_nz(dat9_actv_nz[14]),
.io_dat_actv_9_14_bits_data(dat9_actv_data[119:112]),

.io_dat_actv_9_15_valid(dat9_actv_pvld[15]),
.io_dat_actv_9_15_bits_nz(dat9_actv_nz[15]),
.io_dat_actv_9_15_bits_data(dat9_actv_data[127:120]),

.io_dat_actv_9_16_valid(dat9_actv_pvld[16]),
.io_dat_actv_9_16_bits_nz(dat9_actv_nz[16]),
.io_dat_actv_9_16_bits_data(dat9_actv_data[135:128]),

.io_dat_actv_9_17_valid(dat9_actv_pvld[17]),
.io_dat_actv_9_17_bits_nz(dat9_actv_nz[17]),
.io_dat_actv_9_17_bits_data(dat9_actv_data[143:136]),

.io_dat_actv_9_18_valid(dat9_actv_pvld[18]),
.io_dat_actv_9_18_bits_nz(dat9_actv_nz[18]),
.io_dat_actv_9_18_bits_data(dat9_actv_data[151:144]),

.io_dat_actv_9_19_valid(dat9_actv_pvld[19]),
.io_dat_actv_9_19_bits_nz(dat9_actv_nz[19]),
.io_dat_actv_9_19_bits_data(dat9_actv_data[159:152]),

.io_dat_actv_9_20_valid(dat9_actv_pvld[20]),
.io_dat_actv_9_20_bits_nz(dat9_actv_nz[20]),
.io_dat_actv_9_20_bits_data(dat9_actv_data[167:160]),

.io_dat_actv_9_21_valid(dat9_actv_pvld[21]),
.io_dat_actv_9_21_bits_nz(dat9_actv_nz[21]),
.io_dat_actv_9_21_bits_data(dat9_actv_data[175:168]),

.io_dat_actv_9_22_valid(dat9_actv_pvld[22]),
.io_dat_actv_9_22_bits_nz(dat9_actv_nz[22]),
.io_dat_actv_9_22_bits_data(dat9_actv_data[183:176]),

.io_dat_actv_9_23_valid(dat9_actv_pvld[23]),
.io_dat_actv_9_23_bits_nz(dat9_actv_nz[23]),
.io_dat_actv_9_23_bits_data(dat9_actv_data[191:184]),

.io_dat_actv_9_24_valid(dat9_actv_pvld[24]),
.io_dat_actv_9_24_bits_nz(dat9_actv_nz[24]),
.io_dat_actv_9_24_bits_data(dat9_actv_data[199:192]),

.io_dat_actv_9_25_valid(dat9_actv_pvld[25]),
.io_dat_actv_9_25_bits_nz(dat9_actv_nz[25]),
.io_dat_actv_9_25_bits_data(dat9_actv_data[207:200]),

.io_dat_actv_9_26_valid(dat9_actv_pvld[26]),
.io_dat_actv_9_26_bits_nz(dat9_actv_nz[26]),
.io_dat_actv_9_26_bits_data(dat9_actv_data[215:208]),

.io_dat_actv_9_27_valid(dat9_actv_pvld[27]),
.io_dat_actv_9_27_bits_nz(dat9_actv_nz[27]),
.io_dat_actv_9_27_bits_data(dat9_actv_data[223:216]),

.io_dat_actv_9_28_valid(dat9_actv_pvld[28]),
.io_dat_actv_9_28_bits_nz(dat9_actv_nz[28]),
.io_dat_actv_9_28_bits_data(dat9_actv_data[231:224]),

.io_dat_actv_9_29_valid(dat9_actv_pvld[29]),
.io_dat_actv_9_29_bits_nz(dat9_actv_nz[29]),
.io_dat_actv_9_29_bits_data(dat9_actv_data[239:232]),

.io_dat_actv_9_30_valid(dat9_actv_pvld[30]),
.io_dat_actv_9_30_bits_nz(dat9_actv_nz[30]),
.io_dat_actv_9_30_bits_data(dat9_actv_data[247:240]),

.io_dat_actv_9_31_valid(dat9_actv_pvld[31]),
.io_dat_actv_9_31_bits_nz(dat9_actv_nz[31]),
.io_dat_actv_9_31_bits_data(dat9_actv_data[255:248]),

.io_dat_actv_9_32_valid(dat9_actv_pvld[32]),
.io_dat_actv_9_32_bits_nz(dat9_actv_nz[32]),
.io_dat_actv_9_32_bits_data(dat9_actv_data[263:256]),

.io_dat_actv_9_33_valid(dat9_actv_pvld[33]),
.io_dat_actv_9_33_bits_nz(dat9_actv_nz[33]),
.io_dat_actv_9_33_bits_data(dat9_actv_data[271:264]),

.io_dat_actv_9_34_valid(dat9_actv_pvld[34]),
.io_dat_actv_9_34_bits_nz(dat9_actv_nz[34]),
.io_dat_actv_9_34_bits_data(dat9_actv_data[279:272]),

.io_dat_actv_9_35_valid(dat9_actv_pvld[35]),
.io_dat_actv_9_35_bits_nz(dat9_actv_nz[35]),
.io_dat_actv_9_35_bits_data(dat9_actv_data[287:280]),

.io_dat_actv_9_36_valid(dat9_actv_pvld[36]),
.io_dat_actv_9_36_bits_nz(dat9_actv_nz[36]),
.io_dat_actv_9_36_bits_data(dat9_actv_data[295:288]),

.io_dat_actv_9_37_valid(dat9_actv_pvld[37]),
.io_dat_actv_9_37_bits_nz(dat9_actv_nz[37]),
.io_dat_actv_9_37_bits_data(dat9_actv_data[303:296]),

.io_dat_actv_9_38_valid(dat9_actv_pvld[38]),
.io_dat_actv_9_38_bits_nz(dat9_actv_nz[38]),
.io_dat_actv_9_38_bits_data(dat9_actv_data[311:304]),

.io_dat_actv_9_39_valid(dat9_actv_pvld[39]),
.io_dat_actv_9_39_bits_nz(dat9_actv_nz[39]),
.io_dat_actv_9_39_bits_data(dat9_actv_data[319:312]),

.io_dat_actv_9_40_valid(dat9_actv_pvld[40]),
.io_dat_actv_9_40_bits_nz(dat9_actv_nz[40]),
.io_dat_actv_9_40_bits_data(dat9_actv_data[327:320]),

.io_dat_actv_9_41_valid(dat9_actv_pvld[41]),
.io_dat_actv_9_41_bits_nz(dat9_actv_nz[41]),
.io_dat_actv_9_41_bits_data(dat9_actv_data[335:328]),

.io_dat_actv_9_42_valid(dat9_actv_pvld[42]),
.io_dat_actv_9_42_bits_nz(dat9_actv_nz[42]),
.io_dat_actv_9_42_bits_data(dat9_actv_data[343:336]),

.io_dat_actv_9_43_valid(dat9_actv_pvld[43]),
.io_dat_actv_9_43_bits_nz(dat9_actv_nz[43]),
.io_dat_actv_9_43_bits_data(dat9_actv_data[351:344]),

.io_dat_actv_9_44_valid(dat9_actv_pvld[44]),
.io_dat_actv_9_44_bits_nz(dat9_actv_nz[44]),
.io_dat_actv_9_44_bits_data(dat9_actv_data[359:352]),

.io_dat_actv_9_45_valid(dat9_actv_pvld[45]),
.io_dat_actv_9_45_bits_nz(dat9_actv_nz[45]),
.io_dat_actv_9_45_bits_data(dat9_actv_data[367:360]),

.io_dat_actv_9_46_valid(dat9_actv_pvld[46]),
.io_dat_actv_9_46_bits_nz(dat9_actv_nz[46]),
.io_dat_actv_9_46_bits_data(dat9_actv_data[375:368]),

.io_dat_actv_9_47_valid(dat9_actv_pvld[47]),
.io_dat_actv_9_47_bits_nz(dat9_actv_nz[47]),
.io_dat_actv_9_47_bits_data(dat9_actv_data[383:376]),

.io_dat_actv_9_48_valid(dat9_actv_pvld[48]),
.io_dat_actv_9_48_bits_nz(dat9_actv_nz[48]),
.io_dat_actv_9_48_bits_data(dat9_actv_data[391:384]),

.io_dat_actv_9_49_valid(dat9_actv_pvld[49]),
.io_dat_actv_9_49_bits_nz(dat9_actv_nz[49]),
.io_dat_actv_9_49_bits_data(dat9_actv_data[399:392]),

.io_dat_actv_9_50_valid(dat9_actv_pvld[50]),
.io_dat_actv_9_50_bits_nz(dat9_actv_nz[50]),
.io_dat_actv_9_50_bits_data(dat9_actv_data[407:400]),

.io_dat_actv_9_51_valid(dat9_actv_pvld[51]),
.io_dat_actv_9_51_bits_nz(dat9_actv_nz[51]),
.io_dat_actv_9_51_bits_data(dat9_actv_data[415:408]),

.io_dat_actv_9_52_valid(dat9_actv_pvld[52]),
.io_dat_actv_9_52_bits_nz(dat9_actv_nz[52]),
.io_dat_actv_9_52_bits_data(dat9_actv_data[423:416]),

.io_dat_actv_9_53_valid(dat9_actv_pvld[53]),
.io_dat_actv_9_53_bits_nz(dat9_actv_nz[53]),
.io_dat_actv_9_53_bits_data(dat9_actv_data[431:424]),

.io_dat_actv_9_54_valid(dat9_actv_pvld[54]),
.io_dat_actv_9_54_bits_nz(dat9_actv_nz[54]),
.io_dat_actv_9_54_bits_data(dat9_actv_data[439:432]),

.io_dat_actv_9_55_valid(dat9_actv_pvld[55]),
.io_dat_actv_9_55_bits_nz(dat9_actv_nz[55]),
.io_dat_actv_9_55_bits_data(dat9_actv_data[447:440]),

.io_dat_actv_9_56_valid(dat9_actv_pvld[56]),
.io_dat_actv_9_56_bits_nz(dat9_actv_nz[56]),
.io_dat_actv_9_56_bits_data(dat9_actv_data[455:448]),

.io_dat_actv_9_57_valid(dat9_actv_pvld[57]),
.io_dat_actv_9_57_bits_nz(dat9_actv_nz[57]),
.io_dat_actv_9_57_bits_data(dat9_actv_data[463:456]),

.io_dat_actv_9_58_valid(dat9_actv_pvld[58]),
.io_dat_actv_9_58_bits_nz(dat9_actv_nz[58]),
.io_dat_actv_9_58_bits_data(dat9_actv_data[471:464]),

.io_dat_actv_9_59_valid(dat9_actv_pvld[59]),
.io_dat_actv_9_59_bits_nz(dat9_actv_nz[59]),
.io_dat_actv_9_59_bits_data(dat9_actv_data[479:472]),

.io_dat_actv_9_60_valid(dat9_actv_pvld[60]),
.io_dat_actv_9_60_bits_nz(dat9_actv_nz[60]),
.io_dat_actv_9_60_bits_data(dat9_actv_data[487:480]),

.io_dat_actv_9_61_valid(dat9_actv_pvld[61]),
.io_dat_actv_9_61_bits_nz(dat9_actv_nz[61]),
.io_dat_actv_9_61_bits_data(dat9_actv_data[495:488]),

.io_dat_actv_9_62_valid(dat9_actv_pvld[62]),
.io_dat_actv_9_62_bits_nz(dat9_actv_nz[62]),
.io_dat_actv_9_62_bits_data(dat9_actv_data[503:496]),

.io_dat_actv_9_63_valid(dat9_actv_pvld[63]),
.io_dat_actv_9_63_bits_nz(dat9_actv_nz[63]),
.io_dat_actv_9_63_bits_data(dat9_actv_data[511:504]),

.io_dat_actv_10_0_valid(dat10_actv_pvld[0]),
.io_dat_actv_10_0_bits_nz(dat10_actv_nz[0]),
.io_dat_actv_10_0_bits_data(dat10_actv_data[7:0]),

.io_dat_actv_10_1_valid(dat10_actv_pvld[1]),
.io_dat_actv_10_1_bits_nz(dat10_actv_nz[1]),
.io_dat_actv_10_1_bits_data(dat10_actv_data[15:8]),

.io_dat_actv_10_2_valid(dat10_actv_pvld[2]),
.io_dat_actv_10_2_bits_nz(dat10_actv_nz[2]),
.io_dat_actv_10_2_bits_data(dat10_actv_data[23:16]),

.io_dat_actv_10_3_valid(dat10_actv_pvld[3]),
.io_dat_actv_10_3_bits_nz(dat10_actv_nz[3]),
.io_dat_actv_10_3_bits_data(dat10_actv_data[31:24]),

.io_dat_actv_10_4_valid(dat10_actv_pvld[4]),
.io_dat_actv_10_4_bits_nz(dat10_actv_nz[4]),
.io_dat_actv_10_4_bits_data(dat10_actv_data[39:32]),

.io_dat_actv_10_5_valid(dat10_actv_pvld[5]),
.io_dat_actv_10_5_bits_nz(dat10_actv_nz[5]),
.io_dat_actv_10_5_bits_data(dat10_actv_data[47:40]),

.io_dat_actv_10_6_valid(dat10_actv_pvld[6]),
.io_dat_actv_10_6_bits_nz(dat10_actv_nz[6]),
.io_dat_actv_10_6_bits_data(dat10_actv_data[55:48]),

.io_dat_actv_10_7_valid(dat10_actv_pvld[7]),
.io_dat_actv_10_7_bits_nz(dat10_actv_nz[7]),
.io_dat_actv_10_7_bits_data(dat10_actv_data[63:56]),

.io_dat_actv_10_8_valid(dat10_actv_pvld[8]),
.io_dat_actv_10_8_bits_nz(dat10_actv_nz[8]),
.io_dat_actv_10_8_bits_data(dat10_actv_data[71:64]),

.io_dat_actv_10_9_valid(dat10_actv_pvld[9]),
.io_dat_actv_10_9_bits_nz(dat10_actv_nz[9]),
.io_dat_actv_10_9_bits_data(dat10_actv_data[79:72]),

.io_dat_actv_10_10_valid(dat10_actv_pvld[10]),
.io_dat_actv_10_10_bits_nz(dat10_actv_nz[10]),
.io_dat_actv_10_10_bits_data(dat10_actv_data[87:80]),

.io_dat_actv_10_11_valid(dat10_actv_pvld[11]),
.io_dat_actv_10_11_bits_nz(dat10_actv_nz[11]),
.io_dat_actv_10_11_bits_data(dat10_actv_data[95:88]),

.io_dat_actv_10_12_valid(dat10_actv_pvld[12]),
.io_dat_actv_10_12_bits_nz(dat10_actv_nz[12]),
.io_dat_actv_10_12_bits_data(dat10_actv_data[103:96]),

.io_dat_actv_10_13_valid(dat10_actv_pvld[13]),
.io_dat_actv_10_13_bits_nz(dat10_actv_nz[13]),
.io_dat_actv_10_13_bits_data(dat10_actv_data[111:104]),

.io_dat_actv_10_14_valid(dat10_actv_pvld[14]),
.io_dat_actv_10_14_bits_nz(dat10_actv_nz[14]),
.io_dat_actv_10_14_bits_data(dat10_actv_data[119:112]),

.io_dat_actv_10_15_valid(dat10_actv_pvld[15]),
.io_dat_actv_10_15_bits_nz(dat10_actv_nz[15]),
.io_dat_actv_10_15_bits_data(dat10_actv_data[127:120]),

.io_dat_actv_10_16_valid(dat10_actv_pvld[16]),
.io_dat_actv_10_16_bits_nz(dat10_actv_nz[16]),
.io_dat_actv_10_16_bits_data(dat10_actv_data[135:128]),

.io_dat_actv_10_17_valid(dat10_actv_pvld[17]),
.io_dat_actv_10_17_bits_nz(dat10_actv_nz[17]),
.io_dat_actv_10_17_bits_data(dat10_actv_data[143:136]),

.io_dat_actv_10_18_valid(dat10_actv_pvld[18]),
.io_dat_actv_10_18_bits_nz(dat10_actv_nz[18]),
.io_dat_actv_10_18_bits_data(dat10_actv_data[151:144]),

.io_dat_actv_10_19_valid(dat10_actv_pvld[19]),
.io_dat_actv_10_19_bits_nz(dat10_actv_nz[19]),
.io_dat_actv_10_19_bits_data(dat10_actv_data[159:152]),

.io_dat_actv_10_20_valid(dat10_actv_pvld[20]),
.io_dat_actv_10_20_bits_nz(dat10_actv_nz[20]),
.io_dat_actv_10_20_bits_data(dat10_actv_data[167:160]),

.io_dat_actv_10_21_valid(dat10_actv_pvld[21]),
.io_dat_actv_10_21_bits_nz(dat10_actv_nz[21]),
.io_dat_actv_10_21_bits_data(dat10_actv_data[175:168]),

.io_dat_actv_10_22_valid(dat10_actv_pvld[22]),
.io_dat_actv_10_22_bits_nz(dat10_actv_nz[22]),
.io_dat_actv_10_22_bits_data(dat10_actv_data[183:176]),

.io_dat_actv_10_23_valid(dat10_actv_pvld[23]),
.io_dat_actv_10_23_bits_nz(dat10_actv_nz[23]),
.io_dat_actv_10_23_bits_data(dat10_actv_data[191:184]),

.io_dat_actv_10_24_valid(dat10_actv_pvld[24]),
.io_dat_actv_10_24_bits_nz(dat10_actv_nz[24]),
.io_dat_actv_10_24_bits_data(dat10_actv_data[199:192]),

.io_dat_actv_10_25_valid(dat10_actv_pvld[25]),
.io_dat_actv_10_25_bits_nz(dat10_actv_nz[25]),
.io_dat_actv_10_25_bits_data(dat10_actv_data[207:200]),

.io_dat_actv_10_26_valid(dat10_actv_pvld[26]),
.io_dat_actv_10_26_bits_nz(dat10_actv_nz[26]),
.io_dat_actv_10_26_bits_data(dat10_actv_data[215:208]),

.io_dat_actv_10_27_valid(dat10_actv_pvld[27]),
.io_dat_actv_10_27_bits_nz(dat10_actv_nz[27]),
.io_dat_actv_10_27_bits_data(dat10_actv_data[223:216]),

.io_dat_actv_10_28_valid(dat10_actv_pvld[28]),
.io_dat_actv_10_28_bits_nz(dat10_actv_nz[28]),
.io_dat_actv_10_28_bits_data(dat10_actv_data[231:224]),

.io_dat_actv_10_29_valid(dat10_actv_pvld[29]),
.io_dat_actv_10_29_bits_nz(dat10_actv_nz[29]),
.io_dat_actv_10_29_bits_data(dat10_actv_data[239:232]),

.io_dat_actv_10_30_valid(dat10_actv_pvld[30]),
.io_dat_actv_10_30_bits_nz(dat10_actv_nz[30]),
.io_dat_actv_10_30_bits_data(dat10_actv_data[247:240]),

.io_dat_actv_10_31_valid(dat10_actv_pvld[31]),
.io_dat_actv_10_31_bits_nz(dat10_actv_nz[31]),
.io_dat_actv_10_31_bits_data(dat10_actv_data[255:248]),

.io_dat_actv_10_32_valid(dat10_actv_pvld[32]),
.io_dat_actv_10_32_bits_nz(dat10_actv_nz[32]),
.io_dat_actv_10_32_bits_data(dat10_actv_data[263:256]),

.io_dat_actv_10_33_valid(dat10_actv_pvld[33]),
.io_dat_actv_10_33_bits_nz(dat10_actv_nz[33]),
.io_dat_actv_10_33_bits_data(dat10_actv_data[271:264]),

.io_dat_actv_10_34_valid(dat10_actv_pvld[34]),
.io_dat_actv_10_34_bits_nz(dat10_actv_nz[34]),
.io_dat_actv_10_34_bits_data(dat10_actv_data[279:272]),

.io_dat_actv_10_35_valid(dat10_actv_pvld[35]),
.io_dat_actv_10_35_bits_nz(dat10_actv_nz[35]),
.io_dat_actv_10_35_bits_data(dat10_actv_data[287:280]),

.io_dat_actv_10_36_valid(dat10_actv_pvld[36]),
.io_dat_actv_10_36_bits_nz(dat10_actv_nz[36]),
.io_dat_actv_10_36_bits_data(dat10_actv_data[295:288]),

.io_dat_actv_10_37_valid(dat10_actv_pvld[37]),
.io_dat_actv_10_37_bits_nz(dat10_actv_nz[37]),
.io_dat_actv_10_37_bits_data(dat10_actv_data[303:296]),

.io_dat_actv_10_38_valid(dat10_actv_pvld[38]),
.io_dat_actv_10_38_bits_nz(dat10_actv_nz[38]),
.io_dat_actv_10_38_bits_data(dat10_actv_data[311:304]),

.io_dat_actv_10_39_valid(dat10_actv_pvld[39]),
.io_dat_actv_10_39_bits_nz(dat10_actv_nz[39]),
.io_dat_actv_10_39_bits_data(dat10_actv_data[319:312]),

.io_dat_actv_10_40_valid(dat10_actv_pvld[40]),
.io_dat_actv_10_40_bits_nz(dat10_actv_nz[40]),
.io_dat_actv_10_40_bits_data(dat10_actv_data[327:320]),

.io_dat_actv_10_41_valid(dat10_actv_pvld[41]),
.io_dat_actv_10_41_bits_nz(dat10_actv_nz[41]),
.io_dat_actv_10_41_bits_data(dat10_actv_data[335:328]),

.io_dat_actv_10_42_valid(dat10_actv_pvld[42]),
.io_dat_actv_10_42_bits_nz(dat10_actv_nz[42]),
.io_dat_actv_10_42_bits_data(dat10_actv_data[343:336]),

.io_dat_actv_10_43_valid(dat10_actv_pvld[43]),
.io_dat_actv_10_43_bits_nz(dat10_actv_nz[43]),
.io_dat_actv_10_43_bits_data(dat10_actv_data[351:344]),

.io_dat_actv_10_44_valid(dat10_actv_pvld[44]),
.io_dat_actv_10_44_bits_nz(dat10_actv_nz[44]),
.io_dat_actv_10_44_bits_data(dat10_actv_data[359:352]),

.io_dat_actv_10_45_valid(dat10_actv_pvld[45]),
.io_dat_actv_10_45_bits_nz(dat10_actv_nz[45]),
.io_dat_actv_10_45_bits_data(dat10_actv_data[367:360]),

.io_dat_actv_10_46_valid(dat10_actv_pvld[46]),
.io_dat_actv_10_46_bits_nz(dat10_actv_nz[46]),
.io_dat_actv_10_46_bits_data(dat10_actv_data[375:368]),

.io_dat_actv_10_47_valid(dat10_actv_pvld[47]),
.io_dat_actv_10_47_bits_nz(dat10_actv_nz[47]),
.io_dat_actv_10_47_bits_data(dat10_actv_data[383:376]),

.io_dat_actv_10_48_valid(dat10_actv_pvld[48]),
.io_dat_actv_10_48_bits_nz(dat10_actv_nz[48]),
.io_dat_actv_10_48_bits_data(dat10_actv_data[391:384]),

.io_dat_actv_10_49_valid(dat10_actv_pvld[49]),
.io_dat_actv_10_49_bits_nz(dat10_actv_nz[49]),
.io_dat_actv_10_49_bits_data(dat10_actv_data[399:392]),

.io_dat_actv_10_50_valid(dat10_actv_pvld[50]),
.io_dat_actv_10_50_bits_nz(dat10_actv_nz[50]),
.io_dat_actv_10_50_bits_data(dat10_actv_data[407:400]),

.io_dat_actv_10_51_valid(dat10_actv_pvld[51]),
.io_dat_actv_10_51_bits_nz(dat10_actv_nz[51]),
.io_dat_actv_10_51_bits_data(dat10_actv_data[415:408]),

.io_dat_actv_10_52_valid(dat10_actv_pvld[52]),
.io_dat_actv_10_52_bits_nz(dat10_actv_nz[52]),
.io_dat_actv_10_52_bits_data(dat10_actv_data[423:416]),

.io_dat_actv_10_53_valid(dat10_actv_pvld[53]),
.io_dat_actv_10_53_bits_nz(dat10_actv_nz[53]),
.io_dat_actv_10_53_bits_data(dat10_actv_data[431:424]),

.io_dat_actv_10_54_valid(dat10_actv_pvld[54]),
.io_dat_actv_10_54_bits_nz(dat10_actv_nz[54]),
.io_dat_actv_10_54_bits_data(dat10_actv_data[439:432]),

.io_dat_actv_10_55_valid(dat10_actv_pvld[55]),
.io_dat_actv_10_55_bits_nz(dat10_actv_nz[55]),
.io_dat_actv_10_55_bits_data(dat10_actv_data[447:440]),

.io_dat_actv_10_56_valid(dat10_actv_pvld[56]),
.io_dat_actv_10_56_bits_nz(dat10_actv_nz[56]),
.io_dat_actv_10_56_bits_data(dat10_actv_data[455:448]),

.io_dat_actv_10_57_valid(dat10_actv_pvld[57]),
.io_dat_actv_10_57_bits_nz(dat10_actv_nz[57]),
.io_dat_actv_10_57_bits_data(dat10_actv_data[463:456]),

.io_dat_actv_10_58_valid(dat10_actv_pvld[58]),
.io_dat_actv_10_58_bits_nz(dat10_actv_nz[58]),
.io_dat_actv_10_58_bits_data(dat10_actv_data[471:464]),

.io_dat_actv_10_59_valid(dat10_actv_pvld[59]),
.io_dat_actv_10_59_bits_nz(dat10_actv_nz[59]),
.io_dat_actv_10_59_bits_data(dat10_actv_data[479:472]),

.io_dat_actv_10_60_valid(dat10_actv_pvld[60]),
.io_dat_actv_10_60_bits_nz(dat10_actv_nz[60]),
.io_dat_actv_10_60_bits_data(dat10_actv_data[487:480]),

.io_dat_actv_10_61_valid(dat10_actv_pvld[61]),
.io_dat_actv_10_61_bits_nz(dat10_actv_nz[61]),
.io_dat_actv_10_61_bits_data(dat10_actv_data[495:488]),

.io_dat_actv_10_62_valid(dat10_actv_pvld[62]),
.io_dat_actv_10_62_bits_nz(dat10_actv_nz[62]),
.io_dat_actv_10_62_bits_data(dat10_actv_data[503:496]),

.io_dat_actv_10_63_valid(dat10_actv_pvld[63]),
.io_dat_actv_10_63_bits_nz(dat10_actv_nz[63]),
.io_dat_actv_10_63_bits_data(dat10_actv_data[511:504]),

.io_dat_actv_11_0_valid(dat11_actv_pvld[0]),
.io_dat_actv_11_0_bits_nz(dat11_actv_nz[0]),
.io_dat_actv_11_0_bits_data(dat11_actv_data[7:0]),

.io_dat_actv_11_1_valid(dat11_actv_pvld[1]),
.io_dat_actv_11_1_bits_nz(dat11_actv_nz[1]),
.io_dat_actv_11_1_bits_data(dat11_actv_data[15:8]),

.io_dat_actv_11_2_valid(dat11_actv_pvld[2]),
.io_dat_actv_11_2_bits_nz(dat11_actv_nz[2]),
.io_dat_actv_11_2_bits_data(dat11_actv_data[23:16]),

.io_dat_actv_11_3_valid(dat11_actv_pvld[3]),
.io_dat_actv_11_3_bits_nz(dat11_actv_nz[3]),
.io_dat_actv_11_3_bits_data(dat11_actv_data[31:24]),

.io_dat_actv_11_4_valid(dat11_actv_pvld[4]),
.io_dat_actv_11_4_bits_nz(dat11_actv_nz[4]),
.io_dat_actv_11_4_bits_data(dat11_actv_data[39:32]),

.io_dat_actv_11_5_valid(dat11_actv_pvld[5]),
.io_dat_actv_11_5_bits_nz(dat11_actv_nz[5]),
.io_dat_actv_11_5_bits_data(dat11_actv_data[47:40]),

.io_dat_actv_11_6_valid(dat11_actv_pvld[6]),
.io_dat_actv_11_6_bits_nz(dat11_actv_nz[6]),
.io_dat_actv_11_6_bits_data(dat11_actv_data[55:48]),

.io_dat_actv_11_7_valid(dat11_actv_pvld[7]),
.io_dat_actv_11_7_bits_nz(dat11_actv_nz[7]),
.io_dat_actv_11_7_bits_data(dat11_actv_data[63:56]),

.io_dat_actv_11_8_valid(dat11_actv_pvld[8]),
.io_dat_actv_11_8_bits_nz(dat11_actv_nz[8]),
.io_dat_actv_11_8_bits_data(dat11_actv_data[71:64]),

.io_dat_actv_11_9_valid(dat11_actv_pvld[9]),
.io_dat_actv_11_9_bits_nz(dat11_actv_nz[9]),
.io_dat_actv_11_9_bits_data(dat11_actv_data[79:72]),

.io_dat_actv_11_10_valid(dat11_actv_pvld[10]),
.io_dat_actv_11_10_bits_nz(dat11_actv_nz[10]),
.io_dat_actv_11_10_bits_data(dat11_actv_data[87:80]),

.io_dat_actv_11_11_valid(dat11_actv_pvld[11]),
.io_dat_actv_11_11_bits_nz(dat11_actv_nz[11]),
.io_dat_actv_11_11_bits_data(dat11_actv_data[95:88]),

.io_dat_actv_11_12_valid(dat11_actv_pvld[12]),
.io_dat_actv_11_12_bits_nz(dat11_actv_nz[12]),
.io_dat_actv_11_12_bits_data(dat11_actv_data[103:96]),

.io_dat_actv_11_13_valid(dat11_actv_pvld[13]),
.io_dat_actv_11_13_bits_nz(dat11_actv_nz[13]),
.io_dat_actv_11_13_bits_data(dat11_actv_data[111:104]),

.io_dat_actv_11_14_valid(dat11_actv_pvld[14]),
.io_dat_actv_11_14_bits_nz(dat11_actv_nz[14]),
.io_dat_actv_11_14_bits_data(dat11_actv_data[119:112]),

.io_dat_actv_11_15_valid(dat11_actv_pvld[15]),
.io_dat_actv_11_15_bits_nz(dat11_actv_nz[15]),
.io_dat_actv_11_15_bits_data(dat11_actv_data[127:120]),

.io_dat_actv_11_16_valid(dat11_actv_pvld[16]),
.io_dat_actv_11_16_bits_nz(dat11_actv_nz[16]),
.io_dat_actv_11_16_bits_data(dat11_actv_data[135:128]),

.io_dat_actv_11_17_valid(dat11_actv_pvld[17]),
.io_dat_actv_11_17_bits_nz(dat11_actv_nz[17]),
.io_dat_actv_11_17_bits_data(dat11_actv_data[143:136]),

.io_dat_actv_11_18_valid(dat11_actv_pvld[18]),
.io_dat_actv_11_18_bits_nz(dat11_actv_nz[18]),
.io_dat_actv_11_18_bits_data(dat11_actv_data[151:144]),

.io_dat_actv_11_19_valid(dat11_actv_pvld[19]),
.io_dat_actv_11_19_bits_nz(dat11_actv_nz[19]),
.io_dat_actv_11_19_bits_data(dat11_actv_data[159:152]),

.io_dat_actv_11_20_valid(dat11_actv_pvld[20]),
.io_dat_actv_11_20_bits_nz(dat11_actv_nz[20]),
.io_dat_actv_11_20_bits_data(dat11_actv_data[167:160]),

.io_dat_actv_11_21_valid(dat11_actv_pvld[21]),
.io_dat_actv_11_21_bits_nz(dat11_actv_nz[21]),
.io_dat_actv_11_21_bits_data(dat11_actv_data[175:168]),

.io_dat_actv_11_22_valid(dat11_actv_pvld[22]),
.io_dat_actv_11_22_bits_nz(dat11_actv_nz[22]),
.io_dat_actv_11_22_bits_data(dat11_actv_data[183:176]),

.io_dat_actv_11_23_valid(dat11_actv_pvld[23]),
.io_dat_actv_11_23_bits_nz(dat11_actv_nz[23]),
.io_dat_actv_11_23_bits_data(dat11_actv_data[191:184]),

.io_dat_actv_11_24_valid(dat11_actv_pvld[24]),
.io_dat_actv_11_24_bits_nz(dat11_actv_nz[24]),
.io_dat_actv_11_24_bits_data(dat11_actv_data[199:192]),

.io_dat_actv_11_25_valid(dat11_actv_pvld[25]),
.io_dat_actv_11_25_bits_nz(dat11_actv_nz[25]),
.io_dat_actv_11_25_bits_data(dat11_actv_data[207:200]),

.io_dat_actv_11_26_valid(dat11_actv_pvld[26]),
.io_dat_actv_11_26_bits_nz(dat11_actv_nz[26]),
.io_dat_actv_11_26_bits_data(dat11_actv_data[215:208]),

.io_dat_actv_11_27_valid(dat11_actv_pvld[27]),
.io_dat_actv_11_27_bits_nz(dat11_actv_nz[27]),
.io_dat_actv_11_27_bits_data(dat11_actv_data[223:216]),

.io_dat_actv_11_28_valid(dat11_actv_pvld[28]),
.io_dat_actv_11_28_bits_nz(dat11_actv_nz[28]),
.io_dat_actv_11_28_bits_data(dat11_actv_data[231:224]),

.io_dat_actv_11_29_valid(dat11_actv_pvld[29]),
.io_dat_actv_11_29_bits_nz(dat11_actv_nz[29]),
.io_dat_actv_11_29_bits_data(dat11_actv_data[239:232]),

.io_dat_actv_11_30_valid(dat11_actv_pvld[30]),
.io_dat_actv_11_30_bits_nz(dat11_actv_nz[30]),
.io_dat_actv_11_30_bits_data(dat11_actv_data[247:240]),

.io_dat_actv_11_31_valid(dat11_actv_pvld[31]),
.io_dat_actv_11_31_bits_nz(dat11_actv_nz[31]),
.io_dat_actv_11_31_bits_data(dat11_actv_data[255:248]),

.io_dat_actv_11_32_valid(dat11_actv_pvld[32]),
.io_dat_actv_11_32_bits_nz(dat11_actv_nz[32]),
.io_dat_actv_11_32_bits_data(dat11_actv_data[263:256]),

.io_dat_actv_11_33_valid(dat11_actv_pvld[33]),
.io_dat_actv_11_33_bits_nz(dat11_actv_nz[33]),
.io_dat_actv_11_33_bits_data(dat11_actv_data[271:264]),

.io_dat_actv_11_34_valid(dat11_actv_pvld[34]),
.io_dat_actv_11_34_bits_nz(dat11_actv_nz[34]),
.io_dat_actv_11_34_bits_data(dat11_actv_data[279:272]),

.io_dat_actv_11_35_valid(dat11_actv_pvld[35]),
.io_dat_actv_11_35_bits_nz(dat11_actv_nz[35]),
.io_dat_actv_11_35_bits_data(dat11_actv_data[287:280]),

.io_dat_actv_11_36_valid(dat11_actv_pvld[36]),
.io_dat_actv_11_36_bits_nz(dat11_actv_nz[36]),
.io_dat_actv_11_36_bits_data(dat11_actv_data[295:288]),

.io_dat_actv_11_37_valid(dat11_actv_pvld[37]),
.io_dat_actv_11_37_bits_nz(dat11_actv_nz[37]),
.io_dat_actv_11_37_bits_data(dat11_actv_data[303:296]),

.io_dat_actv_11_38_valid(dat11_actv_pvld[38]),
.io_dat_actv_11_38_bits_nz(dat11_actv_nz[38]),
.io_dat_actv_11_38_bits_data(dat11_actv_data[311:304]),

.io_dat_actv_11_39_valid(dat11_actv_pvld[39]),
.io_dat_actv_11_39_bits_nz(dat11_actv_nz[39]),
.io_dat_actv_11_39_bits_data(dat11_actv_data[319:312]),

.io_dat_actv_11_40_valid(dat11_actv_pvld[40]),
.io_dat_actv_11_40_bits_nz(dat11_actv_nz[40]),
.io_dat_actv_11_40_bits_data(dat11_actv_data[327:320]),

.io_dat_actv_11_41_valid(dat11_actv_pvld[41]),
.io_dat_actv_11_41_bits_nz(dat11_actv_nz[41]),
.io_dat_actv_11_41_bits_data(dat11_actv_data[335:328]),

.io_dat_actv_11_42_valid(dat11_actv_pvld[42]),
.io_dat_actv_11_42_bits_nz(dat11_actv_nz[42]),
.io_dat_actv_11_42_bits_data(dat11_actv_data[343:336]),

.io_dat_actv_11_43_valid(dat11_actv_pvld[43]),
.io_dat_actv_11_43_bits_nz(dat11_actv_nz[43]),
.io_dat_actv_11_43_bits_data(dat11_actv_data[351:344]),

.io_dat_actv_11_44_valid(dat11_actv_pvld[44]),
.io_dat_actv_11_44_bits_nz(dat11_actv_nz[44]),
.io_dat_actv_11_44_bits_data(dat11_actv_data[359:352]),

.io_dat_actv_11_45_valid(dat11_actv_pvld[45]),
.io_dat_actv_11_45_bits_nz(dat11_actv_nz[45]),
.io_dat_actv_11_45_bits_data(dat11_actv_data[367:360]),

.io_dat_actv_11_46_valid(dat11_actv_pvld[46]),
.io_dat_actv_11_46_bits_nz(dat11_actv_nz[46]),
.io_dat_actv_11_46_bits_data(dat11_actv_data[375:368]),

.io_dat_actv_11_47_valid(dat11_actv_pvld[47]),
.io_dat_actv_11_47_bits_nz(dat11_actv_nz[47]),
.io_dat_actv_11_47_bits_data(dat11_actv_data[383:376]),

.io_dat_actv_11_48_valid(dat11_actv_pvld[48]),
.io_dat_actv_11_48_bits_nz(dat11_actv_nz[48]),
.io_dat_actv_11_48_bits_data(dat11_actv_data[391:384]),

.io_dat_actv_11_49_valid(dat11_actv_pvld[49]),
.io_dat_actv_11_49_bits_nz(dat11_actv_nz[49]),
.io_dat_actv_11_49_bits_data(dat11_actv_data[399:392]),

.io_dat_actv_11_50_valid(dat11_actv_pvld[50]),
.io_dat_actv_11_50_bits_nz(dat11_actv_nz[50]),
.io_dat_actv_11_50_bits_data(dat11_actv_data[407:400]),

.io_dat_actv_11_51_valid(dat11_actv_pvld[51]),
.io_dat_actv_11_51_bits_nz(dat11_actv_nz[51]),
.io_dat_actv_11_51_bits_data(dat11_actv_data[415:408]),

.io_dat_actv_11_52_valid(dat11_actv_pvld[52]),
.io_dat_actv_11_52_bits_nz(dat11_actv_nz[52]),
.io_dat_actv_11_52_bits_data(dat11_actv_data[423:416]),

.io_dat_actv_11_53_valid(dat11_actv_pvld[53]),
.io_dat_actv_11_53_bits_nz(dat11_actv_nz[53]),
.io_dat_actv_11_53_bits_data(dat11_actv_data[431:424]),

.io_dat_actv_11_54_valid(dat11_actv_pvld[54]),
.io_dat_actv_11_54_bits_nz(dat11_actv_nz[54]),
.io_dat_actv_11_54_bits_data(dat11_actv_data[439:432]),

.io_dat_actv_11_55_valid(dat11_actv_pvld[55]),
.io_dat_actv_11_55_bits_nz(dat11_actv_nz[55]),
.io_dat_actv_11_55_bits_data(dat11_actv_data[447:440]),

.io_dat_actv_11_56_valid(dat11_actv_pvld[56]),
.io_dat_actv_11_56_bits_nz(dat11_actv_nz[56]),
.io_dat_actv_11_56_bits_data(dat11_actv_data[455:448]),

.io_dat_actv_11_57_valid(dat11_actv_pvld[57]),
.io_dat_actv_11_57_bits_nz(dat11_actv_nz[57]),
.io_dat_actv_11_57_bits_data(dat11_actv_data[463:456]),

.io_dat_actv_11_58_valid(dat11_actv_pvld[58]),
.io_dat_actv_11_58_bits_nz(dat11_actv_nz[58]),
.io_dat_actv_11_58_bits_data(dat11_actv_data[471:464]),

.io_dat_actv_11_59_valid(dat11_actv_pvld[59]),
.io_dat_actv_11_59_bits_nz(dat11_actv_nz[59]),
.io_dat_actv_11_59_bits_data(dat11_actv_data[479:472]),

.io_dat_actv_11_60_valid(dat11_actv_pvld[60]),
.io_dat_actv_11_60_bits_nz(dat11_actv_nz[60]),
.io_dat_actv_11_60_bits_data(dat11_actv_data[487:480]),

.io_dat_actv_11_61_valid(dat11_actv_pvld[61]),
.io_dat_actv_11_61_bits_nz(dat11_actv_nz[61]),
.io_dat_actv_11_61_bits_data(dat11_actv_data[495:488]),

.io_dat_actv_11_62_valid(dat11_actv_pvld[62]),
.io_dat_actv_11_62_bits_nz(dat11_actv_nz[62]),
.io_dat_actv_11_62_bits_data(dat11_actv_data[503:496]),

.io_dat_actv_11_63_valid(dat11_actv_pvld[63]),
.io_dat_actv_11_63_bits_nz(dat11_actv_nz[63]),
.io_dat_actv_11_63_bits_data(dat11_actv_data[511:504]),

.io_dat_actv_12_0_valid(dat12_actv_pvld[0]),
.io_dat_actv_12_0_bits_nz(dat12_actv_nz[0]),
.io_dat_actv_12_0_bits_data(dat12_actv_data[7:0]),

.io_dat_actv_12_1_valid(dat12_actv_pvld[1]),
.io_dat_actv_12_1_bits_nz(dat12_actv_nz[1]),
.io_dat_actv_12_1_bits_data(dat12_actv_data[15:8]),

.io_dat_actv_12_2_valid(dat12_actv_pvld[2]),
.io_dat_actv_12_2_bits_nz(dat12_actv_nz[2]),
.io_dat_actv_12_2_bits_data(dat12_actv_data[23:16]),

.io_dat_actv_12_3_valid(dat12_actv_pvld[3]),
.io_dat_actv_12_3_bits_nz(dat12_actv_nz[3]),
.io_dat_actv_12_3_bits_data(dat12_actv_data[31:24]),

.io_dat_actv_12_4_valid(dat12_actv_pvld[4]),
.io_dat_actv_12_4_bits_nz(dat12_actv_nz[4]),
.io_dat_actv_12_4_bits_data(dat12_actv_data[39:32]),

.io_dat_actv_12_5_valid(dat12_actv_pvld[5]),
.io_dat_actv_12_5_bits_nz(dat12_actv_nz[5]),
.io_dat_actv_12_5_bits_data(dat12_actv_data[47:40]),

.io_dat_actv_12_6_valid(dat12_actv_pvld[6]),
.io_dat_actv_12_6_bits_nz(dat12_actv_nz[6]),
.io_dat_actv_12_6_bits_data(dat12_actv_data[55:48]),

.io_dat_actv_12_7_valid(dat12_actv_pvld[7]),
.io_dat_actv_12_7_bits_nz(dat12_actv_nz[7]),
.io_dat_actv_12_7_bits_data(dat12_actv_data[63:56]),

.io_dat_actv_12_8_valid(dat12_actv_pvld[8]),
.io_dat_actv_12_8_bits_nz(dat12_actv_nz[8]),
.io_dat_actv_12_8_bits_data(dat12_actv_data[71:64]),

.io_dat_actv_12_9_valid(dat12_actv_pvld[9]),
.io_dat_actv_12_9_bits_nz(dat12_actv_nz[9]),
.io_dat_actv_12_9_bits_data(dat12_actv_data[79:72]),

.io_dat_actv_12_10_valid(dat12_actv_pvld[10]),
.io_dat_actv_12_10_bits_nz(dat12_actv_nz[10]),
.io_dat_actv_12_10_bits_data(dat12_actv_data[87:80]),

.io_dat_actv_12_11_valid(dat12_actv_pvld[11]),
.io_dat_actv_12_11_bits_nz(dat12_actv_nz[11]),
.io_dat_actv_12_11_bits_data(dat12_actv_data[95:88]),

.io_dat_actv_12_12_valid(dat12_actv_pvld[12]),
.io_dat_actv_12_12_bits_nz(dat12_actv_nz[12]),
.io_dat_actv_12_12_bits_data(dat12_actv_data[103:96]),

.io_dat_actv_12_13_valid(dat12_actv_pvld[13]),
.io_dat_actv_12_13_bits_nz(dat12_actv_nz[13]),
.io_dat_actv_12_13_bits_data(dat12_actv_data[111:104]),

.io_dat_actv_12_14_valid(dat12_actv_pvld[14]),
.io_dat_actv_12_14_bits_nz(dat12_actv_nz[14]),
.io_dat_actv_12_14_bits_data(dat12_actv_data[119:112]),

.io_dat_actv_12_15_valid(dat12_actv_pvld[15]),
.io_dat_actv_12_15_bits_nz(dat12_actv_nz[15]),
.io_dat_actv_12_15_bits_data(dat12_actv_data[127:120]),

.io_dat_actv_12_16_valid(dat12_actv_pvld[16]),
.io_dat_actv_12_16_bits_nz(dat12_actv_nz[16]),
.io_dat_actv_12_16_bits_data(dat12_actv_data[135:128]),

.io_dat_actv_12_17_valid(dat12_actv_pvld[17]),
.io_dat_actv_12_17_bits_nz(dat12_actv_nz[17]),
.io_dat_actv_12_17_bits_data(dat12_actv_data[143:136]),

.io_dat_actv_12_18_valid(dat12_actv_pvld[18]),
.io_dat_actv_12_18_bits_nz(dat12_actv_nz[18]),
.io_dat_actv_12_18_bits_data(dat12_actv_data[151:144]),

.io_dat_actv_12_19_valid(dat12_actv_pvld[19]),
.io_dat_actv_12_19_bits_nz(dat12_actv_nz[19]),
.io_dat_actv_12_19_bits_data(dat12_actv_data[159:152]),

.io_dat_actv_12_20_valid(dat12_actv_pvld[20]),
.io_dat_actv_12_20_bits_nz(dat12_actv_nz[20]),
.io_dat_actv_12_20_bits_data(dat12_actv_data[167:160]),

.io_dat_actv_12_21_valid(dat12_actv_pvld[21]),
.io_dat_actv_12_21_bits_nz(dat12_actv_nz[21]),
.io_dat_actv_12_21_bits_data(dat12_actv_data[175:168]),

.io_dat_actv_12_22_valid(dat12_actv_pvld[22]),
.io_dat_actv_12_22_bits_nz(dat12_actv_nz[22]),
.io_dat_actv_12_22_bits_data(dat12_actv_data[183:176]),

.io_dat_actv_12_23_valid(dat12_actv_pvld[23]),
.io_dat_actv_12_23_bits_nz(dat12_actv_nz[23]),
.io_dat_actv_12_23_bits_data(dat12_actv_data[191:184]),

.io_dat_actv_12_24_valid(dat12_actv_pvld[24]),
.io_dat_actv_12_24_bits_nz(dat12_actv_nz[24]),
.io_dat_actv_12_24_bits_data(dat12_actv_data[199:192]),

.io_dat_actv_12_25_valid(dat12_actv_pvld[25]),
.io_dat_actv_12_25_bits_nz(dat12_actv_nz[25]),
.io_dat_actv_12_25_bits_data(dat12_actv_data[207:200]),

.io_dat_actv_12_26_valid(dat12_actv_pvld[26]),
.io_dat_actv_12_26_bits_nz(dat12_actv_nz[26]),
.io_dat_actv_12_26_bits_data(dat12_actv_data[215:208]),

.io_dat_actv_12_27_valid(dat12_actv_pvld[27]),
.io_dat_actv_12_27_bits_nz(dat12_actv_nz[27]),
.io_dat_actv_12_27_bits_data(dat12_actv_data[223:216]),

.io_dat_actv_12_28_valid(dat12_actv_pvld[28]),
.io_dat_actv_12_28_bits_nz(dat12_actv_nz[28]),
.io_dat_actv_12_28_bits_data(dat12_actv_data[231:224]),

.io_dat_actv_12_29_valid(dat12_actv_pvld[29]),
.io_dat_actv_12_29_bits_nz(dat12_actv_nz[29]),
.io_dat_actv_12_29_bits_data(dat12_actv_data[239:232]),

.io_dat_actv_12_30_valid(dat12_actv_pvld[30]),
.io_dat_actv_12_30_bits_nz(dat12_actv_nz[30]),
.io_dat_actv_12_30_bits_data(dat12_actv_data[247:240]),

.io_dat_actv_12_31_valid(dat12_actv_pvld[31]),
.io_dat_actv_12_31_bits_nz(dat12_actv_nz[31]),
.io_dat_actv_12_31_bits_data(dat12_actv_data[255:248]),

.io_dat_actv_12_32_valid(dat12_actv_pvld[32]),
.io_dat_actv_12_32_bits_nz(dat12_actv_nz[32]),
.io_dat_actv_12_32_bits_data(dat12_actv_data[263:256]),

.io_dat_actv_12_33_valid(dat12_actv_pvld[33]),
.io_dat_actv_12_33_bits_nz(dat12_actv_nz[33]),
.io_dat_actv_12_33_bits_data(dat12_actv_data[271:264]),

.io_dat_actv_12_34_valid(dat12_actv_pvld[34]),
.io_dat_actv_12_34_bits_nz(dat12_actv_nz[34]),
.io_dat_actv_12_34_bits_data(dat12_actv_data[279:272]),

.io_dat_actv_12_35_valid(dat12_actv_pvld[35]),
.io_dat_actv_12_35_bits_nz(dat12_actv_nz[35]),
.io_dat_actv_12_35_bits_data(dat12_actv_data[287:280]),

.io_dat_actv_12_36_valid(dat12_actv_pvld[36]),
.io_dat_actv_12_36_bits_nz(dat12_actv_nz[36]),
.io_dat_actv_12_36_bits_data(dat12_actv_data[295:288]),

.io_dat_actv_12_37_valid(dat12_actv_pvld[37]),
.io_dat_actv_12_37_bits_nz(dat12_actv_nz[37]),
.io_dat_actv_12_37_bits_data(dat12_actv_data[303:296]),

.io_dat_actv_12_38_valid(dat12_actv_pvld[38]),
.io_dat_actv_12_38_bits_nz(dat12_actv_nz[38]),
.io_dat_actv_12_38_bits_data(dat12_actv_data[311:304]),

.io_dat_actv_12_39_valid(dat12_actv_pvld[39]),
.io_dat_actv_12_39_bits_nz(dat12_actv_nz[39]),
.io_dat_actv_12_39_bits_data(dat12_actv_data[319:312]),

.io_dat_actv_12_40_valid(dat12_actv_pvld[40]),
.io_dat_actv_12_40_bits_nz(dat12_actv_nz[40]),
.io_dat_actv_12_40_bits_data(dat12_actv_data[327:320]),

.io_dat_actv_12_41_valid(dat12_actv_pvld[41]),
.io_dat_actv_12_41_bits_nz(dat12_actv_nz[41]),
.io_dat_actv_12_41_bits_data(dat12_actv_data[335:328]),

.io_dat_actv_12_42_valid(dat12_actv_pvld[42]),
.io_dat_actv_12_42_bits_nz(dat12_actv_nz[42]),
.io_dat_actv_12_42_bits_data(dat12_actv_data[343:336]),

.io_dat_actv_12_43_valid(dat12_actv_pvld[43]),
.io_dat_actv_12_43_bits_nz(dat12_actv_nz[43]),
.io_dat_actv_12_43_bits_data(dat12_actv_data[351:344]),

.io_dat_actv_12_44_valid(dat12_actv_pvld[44]),
.io_dat_actv_12_44_bits_nz(dat12_actv_nz[44]),
.io_dat_actv_12_44_bits_data(dat12_actv_data[359:352]),

.io_dat_actv_12_45_valid(dat12_actv_pvld[45]),
.io_dat_actv_12_45_bits_nz(dat12_actv_nz[45]),
.io_dat_actv_12_45_bits_data(dat12_actv_data[367:360]),

.io_dat_actv_12_46_valid(dat12_actv_pvld[46]),
.io_dat_actv_12_46_bits_nz(dat12_actv_nz[46]),
.io_dat_actv_12_46_bits_data(dat12_actv_data[375:368]),

.io_dat_actv_12_47_valid(dat12_actv_pvld[47]),
.io_dat_actv_12_47_bits_nz(dat12_actv_nz[47]),
.io_dat_actv_12_47_bits_data(dat12_actv_data[383:376]),

.io_dat_actv_12_48_valid(dat12_actv_pvld[48]),
.io_dat_actv_12_48_bits_nz(dat12_actv_nz[48]),
.io_dat_actv_12_48_bits_data(dat12_actv_data[391:384]),

.io_dat_actv_12_49_valid(dat12_actv_pvld[49]),
.io_dat_actv_12_49_bits_nz(dat12_actv_nz[49]),
.io_dat_actv_12_49_bits_data(dat12_actv_data[399:392]),

.io_dat_actv_12_50_valid(dat12_actv_pvld[50]),
.io_dat_actv_12_50_bits_nz(dat12_actv_nz[50]),
.io_dat_actv_12_50_bits_data(dat12_actv_data[407:400]),

.io_dat_actv_12_51_valid(dat12_actv_pvld[51]),
.io_dat_actv_12_51_bits_nz(dat12_actv_nz[51]),
.io_dat_actv_12_51_bits_data(dat12_actv_data[415:408]),

.io_dat_actv_12_52_valid(dat12_actv_pvld[52]),
.io_dat_actv_12_52_bits_nz(dat12_actv_nz[52]),
.io_dat_actv_12_52_bits_data(dat12_actv_data[423:416]),

.io_dat_actv_12_53_valid(dat12_actv_pvld[53]),
.io_dat_actv_12_53_bits_nz(dat12_actv_nz[53]),
.io_dat_actv_12_53_bits_data(dat12_actv_data[431:424]),

.io_dat_actv_12_54_valid(dat12_actv_pvld[54]),
.io_dat_actv_12_54_bits_nz(dat12_actv_nz[54]),
.io_dat_actv_12_54_bits_data(dat12_actv_data[439:432]),

.io_dat_actv_12_55_valid(dat12_actv_pvld[55]),
.io_dat_actv_12_55_bits_nz(dat12_actv_nz[55]),
.io_dat_actv_12_55_bits_data(dat12_actv_data[447:440]),

.io_dat_actv_12_56_valid(dat12_actv_pvld[56]),
.io_dat_actv_12_56_bits_nz(dat12_actv_nz[56]),
.io_dat_actv_12_56_bits_data(dat12_actv_data[455:448]),

.io_dat_actv_12_57_valid(dat12_actv_pvld[57]),
.io_dat_actv_12_57_bits_nz(dat12_actv_nz[57]),
.io_dat_actv_12_57_bits_data(dat12_actv_data[463:456]),

.io_dat_actv_12_58_valid(dat12_actv_pvld[58]),
.io_dat_actv_12_58_bits_nz(dat12_actv_nz[58]),
.io_dat_actv_12_58_bits_data(dat12_actv_data[471:464]),

.io_dat_actv_12_59_valid(dat12_actv_pvld[59]),
.io_dat_actv_12_59_bits_nz(dat12_actv_nz[59]),
.io_dat_actv_12_59_bits_data(dat12_actv_data[479:472]),

.io_dat_actv_12_60_valid(dat12_actv_pvld[60]),
.io_dat_actv_12_60_bits_nz(dat12_actv_nz[60]),
.io_dat_actv_12_60_bits_data(dat12_actv_data[487:480]),

.io_dat_actv_12_61_valid(dat12_actv_pvld[61]),
.io_dat_actv_12_61_bits_nz(dat12_actv_nz[61]),
.io_dat_actv_12_61_bits_data(dat12_actv_data[495:488]),

.io_dat_actv_12_62_valid(dat12_actv_pvld[62]),
.io_dat_actv_12_62_bits_nz(dat12_actv_nz[62]),
.io_dat_actv_12_62_bits_data(dat12_actv_data[503:496]),

.io_dat_actv_12_63_valid(dat12_actv_pvld[63]),
.io_dat_actv_12_63_bits_nz(dat12_actv_nz[63]),
.io_dat_actv_12_63_bits_data(dat12_actv_data[511:504]),

.io_dat_actv_13_0_valid(dat13_actv_pvld[0]),
.io_dat_actv_13_0_bits_nz(dat13_actv_nz[0]),
.io_dat_actv_13_0_bits_data(dat13_actv_data[7:0]),

.io_dat_actv_13_1_valid(dat13_actv_pvld[1]),
.io_dat_actv_13_1_bits_nz(dat13_actv_nz[1]),
.io_dat_actv_13_1_bits_data(dat13_actv_data[15:8]),

.io_dat_actv_13_2_valid(dat13_actv_pvld[2]),
.io_dat_actv_13_2_bits_nz(dat13_actv_nz[2]),
.io_dat_actv_13_2_bits_data(dat13_actv_data[23:16]),

.io_dat_actv_13_3_valid(dat13_actv_pvld[3]),
.io_dat_actv_13_3_bits_nz(dat13_actv_nz[3]),
.io_dat_actv_13_3_bits_data(dat13_actv_data[31:24]),

.io_dat_actv_13_4_valid(dat13_actv_pvld[4]),
.io_dat_actv_13_4_bits_nz(dat13_actv_nz[4]),
.io_dat_actv_13_4_bits_data(dat13_actv_data[39:32]),

.io_dat_actv_13_5_valid(dat13_actv_pvld[5]),
.io_dat_actv_13_5_bits_nz(dat13_actv_nz[5]),
.io_dat_actv_13_5_bits_data(dat13_actv_data[47:40]),

.io_dat_actv_13_6_valid(dat13_actv_pvld[6]),
.io_dat_actv_13_6_bits_nz(dat13_actv_nz[6]),
.io_dat_actv_13_6_bits_data(dat13_actv_data[55:48]),

.io_dat_actv_13_7_valid(dat13_actv_pvld[7]),
.io_dat_actv_13_7_bits_nz(dat13_actv_nz[7]),
.io_dat_actv_13_7_bits_data(dat13_actv_data[63:56]),

.io_dat_actv_13_8_valid(dat13_actv_pvld[8]),
.io_dat_actv_13_8_bits_nz(dat13_actv_nz[8]),
.io_dat_actv_13_8_bits_data(dat13_actv_data[71:64]),

.io_dat_actv_13_9_valid(dat13_actv_pvld[9]),
.io_dat_actv_13_9_bits_nz(dat13_actv_nz[9]),
.io_dat_actv_13_9_bits_data(dat13_actv_data[79:72]),

.io_dat_actv_13_10_valid(dat13_actv_pvld[10]),
.io_dat_actv_13_10_bits_nz(dat13_actv_nz[10]),
.io_dat_actv_13_10_bits_data(dat13_actv_data[87:80]),

.io_dat_actv_13_11_valid(dat13_actv_pvld[11]),
.io_dat_actv_13_11_bits_nz(dat13_actv_nz[11]),
.io_dat_actv_13_11_bits_data(dat13_actv_data[95:88]),

.io_dat_actv_13_12_valid(dat13_actv_pvld[12]),
.io_dat_actv_13_12_bits_nz(dat13_actv_nz[12]),
.io_dat_actv_13_12_bits_data(dat13_actv_data[103:96]),

.io_dat_actv_13_13_valid(dat13_actv_pvld[13]),
.io_dat_actv_13_13_bits_nz(dat13_actv_nz[13]),
.io_dat_actv_13_13_bits_data(dat13_actv_data[111:104]),

.io_dat_actv_13_14_valid(dat13_actv_pvld[14]),
.io_dat_actv_13_14_bits_nz(dat13_actv_nz[14]),
.io_dat_actv_13_14_bits_data(dat13_actv_data[119:112]),

.io_dat_actv_13_15_valid(dat13_actv_pvld[15]),
.io_dat_actv_13_15_bits_nz(dat13_actv_nz[15]),
.io_dat_actv_13_15_bits_data(dat13_actv_data[127:120]),

.io_dat_actv_13_16_valid(dat13_actv_pvld[16]),
.io_dat_actv_13_16_bits_nz(dat13_actv_nz[16]),
.io_dat_actv_13_16_bits_data(dat13_actv_data[135:128]),

.io_dat_actv_13_17_valid(dat13_actv_pvld[17]),
.io_dat_actv_13_17_bits_nz(dat13_actv_nz[17]),
.io_dat_actv_13_17_bits_data(dat13_actv_data[143:136]),

.io_dat_actv_13_18_valid(dat13_actv_pvld[18]),
.io_dat_actv_13_18_bits_nz(dat13_actv_nz[18]),
.io_dat_actv_13_18_bits_data(dat13_actv_data[151:144]),

.io_dat_actv_13_19_valid(dat13_actv_pvld[19]),
.io_dat_actv_13_19_bits_nz(dat13_actv_nz[19]),
.io_dat_actv_13_19_bits_data(dat13_actv_data[159:152]),

.io_dat_actv_13_20_valid(dat13_actv_pvld[20]),
.io_dat_actv_13_20_bits_nz(dat13_actv_nz[20]),
.io_dat_actv_13_20_bits_data(dat13_actv_data[167:160]),

.io_dat_actv_13_21_valid(dat13_actv_pvld[21]),
.io_dat_actv_13_21_bits_nz(dat13_actv_nz[21]),
.io_dat_actv_13_21_bits_data(dat13_actv_data[175:168]),

.io_dat_actv_13_22_valid(dat13_actv_pvld[22]),
.io_dat_actv_13_22_bits_nz(dat13_actv_nz[22]),
.io_dat_actv_13_22_bits_data(dat13_actv_data[183:176]),

.io_dat_actv_13_23_valid(dat13_actv_pvld[23]),
.io_dat_actv_13_23_bits_nz(dat13_actv_nz[23]),
.io_dat_actv_13_23_bits_data(dat13_actv_data[191:184]),

.io_dat_actv_13_24_valid(dat13_actv_pvld[24]),
.io_dat_actv_13_24_bits_nz(dat13_actv_nz[24]),
.io_dat_actv_13_24_bits_data(dat13_actv_data[199:192]),

.io_dat_actv_13_25_valid(dat13_actv_pvld[25]),
.io_dat_actv_13_25_bits_nz(dat13_actv_nz[25]),
.io_dat_actv_13_25_bits_data(dat13_actv_data[207:200]),

.io_dat_actv_13_26_valid(dat13_actv_pvld[26]),
.io_dat_actv_13_26_bits_nz(dat13_actv_nz[26]),
.io_dat_actv_13_26_bits_data(dat13_actv_data[215:208]),

.io_dat_actv_13_27_valid(dat13_actv_pvld[27]),
.io_dat_actv_13_27_bits_nz(dat13_actv_nz[27]),
.io_dat_actv_13_27_bits_data(dat13_actv_data[223:216]),

.io_dat_actv_13_28_valid(dat13_actv_pvld[28]),
.io_dat_actv_13_28_bits_nz(dat13_actv_nz[28]),
.io_dat_actv_13_28_bits_data(dat13_actv_data[231:224]),

.io_dat_actv_13_29_valid(dat13_actv_pvld[29]),
.io_dat_actv_13_29_bits_nz(dat13_actv_nz[29]),
.io_dat_actv_13_29_bits_data(dat13_actv_data[239:232]),

.io_dat_actv_13_30_valid(dat13_actv_pvld[30]),
.io_dat_actv_13_30_bits_nz(dat13_actv_nz[30]),
.io_dat_actv_13_30_bits_data(dat13_actv_data[247:240]),

.io_dat_actv_13_31_valid(dat13_actv_pvld[31]),
.io_dat_actv_13_31_bits_nz(dat13_actv_nz[31]),
.io_dat_actv_13_31_bits_data(dat13_actv_data[255:248]),

.io_dat_actv_13_32_valid(dat13_actv_pvld[32]),
.io_dat_actv_13_32_bits_nz(dat13_actv_nz[32]),
.io_dat_actv_13_32_bits_data(dat13_actv_data[263:256]),

.io_dat_actv_13_33_valid(dat13_actv_pvld[33]),
.io_dat_actv_13_33_bits_nz(dat13_actv_nz[33]),
.io_dat_actv_13_33_bits_data(dat13_actv_data[271:264]),

.io_dat_actv_13_34_valid(dat13_actv_pvld[34]),
.io_dat_actv_13_34_bits_nz(dat13_actv_nz[34]),
.io_dat_actv_13_34_bits_data(dat13_actv_data[279:272]),

.io_dat_actv_13_35_valid(dat13_actv_pvld[35]),
.io_dat_actv_13_35_bits_nz(dat13_actv_nz[35]),
.io_dat_actv_13_35_bits_data(dat13_actv_data[287:280]),

.io_dat_actv_13_36_valid(dat13_actv_pvld[36]),
.io_dat_actv_13_36_bits_nz(dat13_actv_nz[36]),
.io_dat_actv_13_36_bits_data(dat13_actv_data[295:288]),

.io_dat_actv_13_37_valid(dat13_actv_pvld[37]),
.io_dat_actv_13_37_bits_nz(dat13_actv_nz[37]),
.io_dat_actv_13_37_bits_data(dat13_actv_data[303:296]),

.io_dat_actv_13_38_valid(dat13_actv_pvld[38]),
.io_dat_actv_13_38_bits_nz(dat13_actv_nz[38]),
.io_dat_actv_13_38_bits_data(dat13_actv_data[311:304]),

.io_dat_actv_13_39_valid(dat13_actv_pvld[39]),
.io_dat_actv_13_39_bits_nz(dat13_actv_nz[39]),
.io_dat_actv_13_39_bits_data(dat13_actv_data[319:312]),

.io_dat_actv_13_40_valid(dat13_actv_pvld[40]),
.io_dat_actv_13_40_bits_nz(dat13_actv_nz[40]),
.io_dat_actv_13_40_bits_data(dat13_actv_data[327:320]),

.io_dat_actv_13_41_valid(dat13_actv_pvld[41]),
.io_dat_actv_13_41_bits_nz(dat13_actv_nz[41]),
.io_dat_actv_13_41_bits_data(dat13_actv_data[335:328]),

.io_dat_actv_13_42_valid(dat13_actv_pvld[42]),
.io_dat_actv_13_42_bits_nz(dat13_actv_nz[42]),
.io_dat_actv_13_42_bits_data(dat13_actv_data[343:336]),

.io_dat_actv_13_43_valid(dat13_actv_pvld[43]),
.io_dat_actv_13_43_bits_nz(dat13_actv_nz[43]),
.io_dat_actv_13_43_bits_data(dat13_actv_data[351:344]),

.io_dat_actv_13_44_valid(dat13_actv_pvld[44]),
.io_dat_actv_13_44_bits_nz(dat13_actv_nz[44]),
.io_dat_actv_13_44_bits_data(dat13_actv_data[359:352]),

.io_dat_actv_13_45_valid(dat13_actv_pvld[45]),
.io_dat_actv_13_45_bits_nz(dat13_actv_nz[45]),
.io_dat_actv_13_45_bits_data(dat13_actv_data[367:360]),

.io_dat_actv_13_46_valid(dat13_actv_pvld[46]),
.io_dat_actv_13_46_bits_nz(dat13_actv_nz[46]),
.io_dat_actv_13_46_bits_data(dat13_actv_data[375:368]),

.io_dat_actv_13_47_valid(dat13_actv_pvld[47]),
.io_dat_actv_13_47_bits_nz(dat13_actv_nz[47]),
.io_dat_actv_13_47_bits_data(dat13_actv_data[383:376]),

.io_dat_actv_13_48_valid(dat13_actv_pvld[48]),
.io_dat_actv_13_48_bits_nz(dat13_actv_nz[48]),
.io_dat_actv_13_48_bits_data(dat13_actv_data[391:384]),

.io_dat_actv_13_49_valid(dat13_actv_pvld[49]),
.io_dat_actv_13_49_bits_nz(dat13_actv_nz[49]),
.io_dat_actv_13_49_bits_data(dat13_actv_data[399:392]),

.io_dat_actv_13_50_valid(dat13_actv_pvld[50]),
.io_dat_actv_13_50_bits_nz(dat13_actv_nz[50]),
.io_dat_actv_13_50_bits_data(dat13_actv_data[407:400]),

.io_dat_actv_13_51_valid(dat13_actv_pvld[51]),
.io_dat_actv_13_51_bits_nz(dat13_actv_nz[51]),
.io_dat_actv_13_51_bits_data(dat13_actv_data[415:408]),

.io_dat_actv_13_52_valid(dat13_actv_pvld[52]),
.io_dat_actv_13_52_bits_nz(dat13_actv_nz[52]),
.io_dat_actv_13_52_bits_data(dat13_actv_data[423:416]),

.io_dat_actv_13_53_valid(dat13_actv_pvld[53]),
.io_dat_actv_13_53_bits_nz(dat13_actv_nz[53]),
.io_dat_actv_13_53_bits_data(dat13_actv_data[431:424]),

.io_dat_actv_13_54_valid(dat13_actv_pvld[54]),
.io_dat_actv_13_54_bits_nz(dat13_actv_nz[54]),
.io_dat_actv_13_54_bits_data(dat13_actv_data[439:432]),

.io_dat_actv_13_55_valid(dat13_actv_pvld[55]),
.io_dat_actv_13_55_bits_nz(dat13_actv_nz[55]),
.io_dat_actv_13_55_bits_data(dat13_actv_data[447:440]),

.io_dat_actv_13_56_valid(dat13_actv_pvld[56]),
.io_dat_actv_13_56_bits_nz(dat13_actv_nz[56]),
.io_dat_actv_13_56_bits_data(dat13_actv_data[455:448]),

.io_dat_actv_13_57_valid(dat13_actv_pvld[57]),
.io_dat_actv_13_57_bits_nz(dat13_actv_nz[57]),
.io_dat_actv_13_57_bits_data(dat13_actv_data[463:456]),

.io_dat_actv_13_58_valid(dat13_actv_pvld[58]),
.io_dat_actv_13_58_bits_nz(dat13_actv_nz[58]),
.io_dat_actv_13_58_bits_data(dat13_actv_data[471:464]),

.io_dat_actv_13_59_valid(dat13_actv_pvld[59]),
.io_dat_actv_13_59_bits_nz(dat13_actv_nz[59]),
.io_dat_actv_13_59_bits_data(dat13_actv_data[479:472]),

.io_dat_actv_13_60_valid(dat13_actv_pvld[60]),
.io_dat_actv_13_60_bits_nz(dat13_actv_nz[60]),
.io_dat_actv_13_60_bits_data(dat13_actv_data[487:480]),

.io_dat_actv_13_61_valid(dat13_actv_pvld[61]),
.io_dat_actv_13_61_bits_nz(dat13_actv_nz[61]),
.io_dat_actv_13_61_bits_data(dat13_actv_data[495:488]),

.io_dat_actv_13_62_valid(dat13_actv_pvld[62]),
.io_dat_actv_13_62_bits_nz(dat13_actv_nz[62]),
.io_dat_actv_13_62_bits_data(dat13_actv_data[503:496]),

.io_dat_actv_13_63_valid(dat13_actv_pvld[63]),
.io_dat_actv_13_63_bits_nz(dat13_actv_nz[63]),
.io_dat_actv_13_63_bits_data(dat13_actv_data[511:504]),

.io_dat_actv_14_0_valid(dat14_actv_pvld[0]),
.io_dat_actv_14_0_bits_nz(dat14_actv_nz[0]),
.io_dat_actv_14_0_bits_data(dat14_actv_data[7:0]),

.io_dat_actv_14_1_valid(dat14_actv_pvld[1]),
.io_dat_actv_14_1_bits_nz(dat14_actv_nz[1]),
.io_dat_actv_14_1_bits_data(dat14_actv_data[15:8]),

.io_dat_actv_14_2_valid(dat14_actv_pvld[2]),
.io_dat_actv_14_2_bits_nz(dat14_actv_nz[2]),
.io_dat_actv_14_2_bits_data(dat14_actv_data[23:16]),

.io_dat_actv_14_3_valid(dat14_actv_pvld[3]),
.io_dat_actv_14_3_bits_nz(dat14_actv_nz[3]),
.io_dat_actv_14_3_bits_data(dat14_actv_data[31:24]),

.io_dat_actv_14_4_valid(dat14_actv_pvld[4]),
.io_dat_actv_14_4_bits_nz(dat14_actv_nz[4]),
.io_dat_actv_14_4_bits_data(dat14_actv_data[39:32]),

.io_dat_actv_14_5_valid(dat14_actv_pvld[5]),
.io_dat_actv_14_5_bits_nz(dat14_actv_nz[5]),
.io_dat_actv_14_5_bits_data(dat14_actv_data[47:40]),

.io_dat_actv_14_6_valid(dat14_actv_pvld[6]),
.io_dat_actv_14_6_bits_nz(dat14_actv_nz[6]),
.io_dat_actv_14_6_bits_data(dat14_actv_data[55:48]),

.io_dat_actv_14_7_valid(dat14_actv_pvld[7]),
.io_dat_actv_14_7_bits_nz(dat14_actv_nz[7]),
.io_dat_actv_14_7_bits_data(dat14_actv_data[63:56]),

.io_dat_actv_14_8_valid(dat14_actv_pvld[8]),
.io_dat_actv_14_8_bits_nz(dat14_actv_nz[8]),
.io_dat_actv_14_8_bits_data(dat14_actv_data[71:64]),

.io_dat_actv_14_9_valid(dat14_actv_pvld[9]),
.io_dat_actv_14_9_bits_nz(dat14_actv_nz[9]),
.io_dat_actv_14_9_bits_data(dat14_actv_data[79:72]),

.io_dat_actv_14_10_valid(dat14_actv_pvld[10]),
.io_dat_actv_14_10_bits_nz(dat14_actv_nz[10]),
.io_dat_actv_14_10_bits_data(dat14_actv_data[87:80]),

.io_dat_actv_14_11_valid(dat14_actv_pvld[11]),
.io_dat_actv_14_11_bits_nz(dat14_actv_nz[11]),
.io_dat_actv_14_11_bits_data(dat14_actv_data[95:88]),

.io_dat_actv_14_12_valid(dat14_actv_pvld[12]),
.io_dat_actv_14_12_bits_nz(dat14_actv_nz[12]),
.io_dat_actv_14_12_bits_data(dat14_actv_data[103:96]),

.io_dat_actv_14_13_valid(dat14_actv_pvld[13]),
.io_dat_actv_14_13_bits_nz(dat14_actv_nz[13]),
.io_dat_actv_14_13_bits_data(dat14_actv_data[111:104]),

.io_dat_actv_14_14_valid(dat14_actv_pvld[14]),
.io_dat_actv_14_14_bits_nz(dat14_actv_nz[14]),
.io_dat_actv_14_14_bits_data(dat14_actv_data[119:112]),

.io_dat_actv_14_15_valid(dat14_actv_pvld[15]),
.io_dat_actv_14_15_bits_nz(dat14_actv_nz[15]),
.io_dat_actv_14_15_bits_data(dat14_actv_data[127:120]),

.io_dat_actv_14_16_valid(dat14_actv_pvld[16]),
.io_dat_actv_14_16_bits_nz(dat14_actv_nz[16]),
.io_dat_actv_14_16_bits_data(dat14_actv_data[135:128]),

.io_dat_actv_14_17_valid(dat14_actv_pvld[17]),
.io_dat_actv_14_17_bits_nz(dat14_actv_nz[17]),
.io_dat_actv_14_17_bits_data(dat14_actv_data[143:136]),

.io_dat_actv_14_18_valid(dat14_actv_pvld[18]),
.io_dat_actv_14_18_bits_nz(dat14_actv_nz[18]),
.io_dat_actv_14_18_bits_data(dat14_actv_data[151:144]),

.io_dat_actv_14_19_valid(dat14_actv_pvld[19]),
.io_dat_actv_14_19_bits_nz(dat14_actv_nz[19]),
.io_dat_actv_14_19_bits_data(dat14_actv_data[159:152]),

.io_dat_actv_14_20_valid(dat14_actv_pvld[20]),
.io_dat_actv_14_20_bits_nz(dat14_actv_nz[20]),
.io_dat_actv_14_20_bits_data(dat14_actv_data[167:160]),

.io_dat_actv_14_21_valid(dat14_actv_pvld[21]),
.io_dat_actv_14_21_bits_nz(dat14_actv_nz[21]),
.io_dat_actv_14_21_bits_data(dat14_actv_data[175:168]),

.io_dat_actv_14_22_valid(dat14_actv_pvld[22]),
.io_dat_actv_14_22_bits_nz(dat14_actv_nz[22]),
.io_dat_actv_14_22_bits_data(dat14_actv_data[183:176]),

.io_dat_actv_14_23_valid(dat14_actv_pvld[23]),
.io_dat_actv_14_23_bits_nz(dat14_actv_nz[23]),
.io_dat_actv_14_23_bits_data(dat14_actv_data[191:184]),

.io_dat_actv_14_24_valid(dat14_actv_pvld[24]),
.io_dat_actv_14_24_bits_nz(dat14_actv_nz[24]),
.io_dat_actv_14_24_bits_data(dat14_actv_data[199:192]),

.io_dat_actv_14_25_valid(dat14_actv_pvld[25]),
.io_dat_actv_14_25_bits_nz(dat14_actv_nz[25]),
.io_dat_actv_14_25_bits_data(dat14_actv_data[207:200]),

.io_dat_actv_14_26_valid(dat14_actv_pvld[26]),
.io_dat_actv_14_26_bits_nz(dat14_actv_nz[26]),
.io_dat_actv_14_26_bits_data(dat14_actv_data[215:208]),

.io_dat_actv_14_27_valid(dat14_actv_pvld[27]),
.io_dat_actv_14_27_bits_nz(dat14_actv_nz[27]),
.io_dat_actv_14_27_bits_data(dat14_actv_data[223:216]),

.io_dat_actv_14_28_valid(dat14_actv_pvld[28]),
.io_dat_actv_14_28_bits_nz(dat14_actv_nz[28]),
.io_dat_actv_14_28_bits_data(dat14_actv_data[231:224]),

.io_dat_actv_14_29_valid(dat14_actv_pvld[29]),
.io_dat_actv_14_29_bits_nz(dat14_actv_nz[29]),
.io_dat_actv_14_29_bits_data(dat14_actv_data[239:232]),

.io_dat_actv_14_30_valid(dat14_actv_pvld[30]),
.io_dat_actv_14_30_bits_nz(dat14_actv_nz[30]),
.io_dat_actv_14_30_bits_data(dat14_actv_data[247:240]),

.io_dat_actv_14_31_valid(dat14_actv_pvld[31]),
.io_dat_actv_14_31_bits_nz(dat14_actv_nz[31]),
.io_dat_actv_14_31_bits_data(dat14_actv_data[255:248]),

.io_dat_actv_14_32_valid(dat14_actv_pvld[32]),
.io_dat_actv_14_32_bits_nz(dat14_actv_nz[32]),
.io_dat_actv_14_32_bits_data(dat14_actv_data[263:256]),

.io_dat_actv_14_33_valid(dat14_actv_pvld[33]),
.io_dat_actv_14_33_bits_nz(dat14_actv_nz[33]),
.io_dat_actv_14_33_bits_data(dat14_actv_data[271:264]),

.io_dat_actv_14_34_valid(dat14_actv_pvld[34]),
.io_dat_actv_14_34_bits_nz(dat14_actv_nz[34]),
.io_dat_actv_14_34_bits_data(dat14_actv_data[279:272]),

.io_dat_actv_14_35_valid(dat14_actv_pvld[35]),
.io_dat_actv_14_35_bits_nz(dat14_actv_nz[35]),
.io_dat_actv_14_35_bits_data(dat14_actv_data[287:280]),

.io_dat_actv_14_36_valid(dat14_actv_pvld[36]),
.io_dat_actv_14_36_bits_nz(dat14_actv_nz[36]),
.io_dat_actv_14_36_bits_data(dat14_actv_data[295:288]),

.io_dat_actv_14_37_valid(dat14_actv_pvld[37]),
.io_dat_actv_14_37_bits_nz(dat14_actv_nz[37]),
.io_dat_actv_14_37_bits_data(dat14_actv_data[303:296]),

.io_dat_actv_14_38_valid(dat14_actv_pvld[38]),
.io_dat_actv_14_38_bits_nz(dat14_actv_nz[38]),
.io_dat_actv_14_38_bits_data(dat14_actv_data[311:304]),

.io_dat_actv_14_39_valid(dat14_actv_pvld[39]),
.io_dat_actv_14_39_bits_nz(dat14_actv_nz[39]),
.io_dat_actv_14_39_bits_data(dat14_actv_data[319:312]),

.io_dat_actv_14_40_valid(dat14_actv_pvld[40]),
.io_dat_actv_14_40_bits_nz(dat14_actv_nz[40]),
.io_dat_actv_14_40_bits_data(dat14_actv_data[327:320]),

.io_dat_actv_14_41_valid(dat14_actv_pvld[41]),
.io_dat_actv_14_41_bits_nz(dat14_actv_nz[41]),
.io_dat_actv_14_41_bits_data(dat14_actv_data[335:328]),

.io_dat_actv_14_42_valid(dat14_actv_pvld[42]),
.io_dat_actv_14_42_bits_nz(dat14_actv_nz[42]),
.io_dat_actv_14_42_bits_data(dat14_actv_data[343:336]),

.io_dat_actv_14_43_valid(dat14_actv_pvld[43]),
.io_dat_actv_14_43_bits_nz(dat14_actv_nz[43]),
.io_dat_actv_14_43_bits_data(dat14_actv_data[351:344]),

.io_dat_actv_14_44_valid(dat14_actv_pvld[44]),
.io_dat_actv_14_44_bits_nz(dat14_actv_nz[44]),
.io_dat_actv_14_44_bits_data(dat14_actv_data[359:352]),

.io_dat_actv_14_45_valid(dat14_actv_pvld[45]),
.io_dat_actv_14_45_bits_nz(dat14_actv_nz[45]),
.io_dat_actv_14_45_bits_data(dat14_actv_data[367:360]),

.io_dat_actv_14_46_valid(dat14_actv_pvld[46]),
.io_dat_actv_14_46_bits_nz(dat14_actv_nz[46]),
.io_dat_actv_14_46_bits_data(dat14_actv_data[375:368]),

.io_dat_actv_14_47_valid(dat14_actv_pvld[47]),
.io_dat_actv_14_47_bits_nz(dat14_actv_nz[47]),
.io_dat_actv_14_47_bits_data(dat14_actv_data[383:376]),

.io_dat_actv_14_48_valid(dat14_actv_pvld[48]),
.io_dat_actv_14_48_bits_nz(dat14_actv_nz[48]),
.io_dat_actv_14_48_bits_data(dat14_actv_data[391:384]),

.io_dat_actv_14_49_valid(dat14_actv_pvld[49]),
.io_dat_actv_14_49_bits_nz(dat14_actv_nz[49]),
.io_dat_actv_14_49_bits_data(dat14_actv_data[399:392]),

.io_dat_actv_14_50_valid(dat14_actv_pvld[50]),
.io_dat_actv_14_50_bits_nz(dat14_actv_nz[50]),
.io_dat_actv_14_50_bits_data(dat14_actv_data[407:400]),

.io_dat_actv_14_51_valid(dat14_actv_pvld[51]),
.io_dat_actv_14_51_bits_nz(dat14_actv_nz[51]),
.io_dat_actv_14_51_bits_data(dat14_actv_data[415:408]),

.io_dat_actv_14_52_valid(dat14_actv_pvld[52]),
.io_dat_actv_14_52_bits_nz(dat14_actv_nz[52]),
.io_dat_actv_14_52_bits_data(dat14_actv_data[423:416]),

.io_dat_actv_14_53_valid(dat14_actv_pvld[53]),
.io_dat_actv_14_53_bits_nz(dat14_actv_nz[53]),
.io_dat_actv_14_53_bits_data(dat14_actv_data[431:424]),

.io_dat_actv_14_54_valid(dat14_actv_pvld[54]),
.io_dat_actv_14_54_bits_nz(dat14_actv_nz[54]),
.io_dat_actv_14_54_bits_data(dat14_actv_data[439:432]),

.io_dat_actv_14_55_valid(dat14_actv_pvld[55]),
.io_dat_actv_14_55_bits_nz(dat14_actv_nz[55]),
.io_dat_actv_14_55_bits_data(dat14_actv_data[447:440]),

.io_dat_actv_14_56_valid(dat14_actv_pvld[56]),
.io_dat_actv_14_56_bits_nz(dat14_actv_nz[56]),
.io_dat_actv_14_56_bits_data(dat14_actv_data[455:448]),

.io_dat_actv_14_57_valid(dat14_actv_pvld[57]),
.io_dat_actv_14_57_bits_nz(dat14_actv_nz[57]),
.io_dat_actv_14_57_bits_data(dat14_actv_data[463:456]),

.io_dat_actv_14_58_valid(dat14_actv_pvld[58]),
.io_dat_actv_14_58_bits_nz(dat14_actv_nz[58]),
.io_dat_actv_14_58_bits_data(dat14_actv_data[471:464]),

.io_dat_actv_14_59_valid(dat14_actv_pvld[59]),
.io_dat_actv_14_59_bits_nz(dat14_actv_nz[59]),
.io_dat_actv_14_59_bits_data(dat14_actv_data[479:472]),

.io_dat_actv_14_60_valid(dat14_actv_pvld[60]),
.io_dat_actv_14_60_bits_nz(dat14_actv_nz[60]),
.io_dat_actv_14_60_bits_data(dat14_actv_data[487:480]),

.io_dat_actv_14_61_valid(dat14_actv_pvld[61]),
.io_dat_actv_14_61_bits_nz(dat14_actv_nz[61]),
.io_dat_actv_14_61_bits_data(dat14_actv_data[495:488]),

.io_dat_actv_14_62_valid(dat14_actv_pvld[62]),
.io_dat_actv_14_62_bits_nz(dat14_actv_nz[62]),
.io_dat_actv_14_62_bits_data(dat14_actv_data[503:496]),

.io_dat_actv_14_63_valid(dat14_actv_pvld[63]),
.io_dat_actv_14_63_bits_nz(dat14_actv_nz[63]),
.io_dat_actv_14_63_bits_data(dat14_actv_data[511:504]),

.io_dat_actv_15_0_valid(dat15_actv_pvld[0]),
.io_dat_actv_15_0_bits_nz(dat15_actv_nz[0]),
.io_dat_actv_15_0_bits_data(dat15_actv_data[7:0]),

.io_dat_actv_15_1_valid(dat15_actv_pvld[1]),
.io_dat_actv_15_1_bits_nz(dat15_actv_nz[1]),
.io_dat_actv_15_1_bits_data(dat15_actv_data[15:8]),

.io_dat_actv_15_2_valid(dat15_actv_pvld[2]),
.io_dat_actv_15_2_bits_nz(dat15_actv_nz[2]),
.io_dat_actv_15_2_bits_data(dat15_actv_data[23:16]),

.io_dat_actv_15_3_valid(dat15_actv_pvld[3]),
.io_dat_actv_15_3_bits_nz(dat15_actv_nz[3]),
.io_dat_actv_15_3_bits_data(dat15_actv_data[31:24]),

.io_dat_actv_15_4_valid(dat15_actv_pvld[4]),
.io_dat_actv_15_4_bits_nz(dat15_actv_nz[4]),
.io_dat_actv_15_4_bits_data(dat15_actv_data[39:32]),

.io_dat_actv_15_5_valid(dat15_actv_pvld[5]),
.io_dat_actv_15_5_bits_nz(dat15_actv_nz[5]),
.io_dat_actv_15_5_bits_data(dat15_actv_data[47:40]),

.io_dat_actv_15_6_valid(dat15_actv_pvld[6]),
.io_dat_actv_15_6_bits_nz(dat15_actv_nz[6]),
.io_dat_actv_15_6_bits_data(dat15_actv_data[55:48]),

.io_dat_actv_15_7_valid(dat15_actv_pvld[7]),
.io_dat_actv_15_7_bits_nz(dat15_actv_nz[7]),
.io_dat_actv_15_7_bits_data(dat15_actv_data[63:56]),

.io_dat_actv_15_8_valid(dat15_actv_pvld[8]),
.io_dat_actv_15_8_bits_nz(dat15_actv_nz[8]),
.io_dat_actv_15_8_bits_data(dat15_actv_data[71:64]),

.io_dat_actv_15_9_valid(dat15_actv_pvld[9]),
.io_dat_actv_15_9_bits_nz(dat15_actv_nz[9]),
.io_dat_actv_15_9_bits_data(dat15_actv_data[79:72]),

.io_dat_actv_15_10_valid(dat15_actv_pvld[10]),
.io_dat_actv_15_10_bits_nz(dat15_actv_nz[10]),
.io_dat_actv_15_10_bits_data(dat15_actv_data[87:80]),

.io_dat_actv_15_11_valid(dat15_actv_pvld[11]),
.io_dat_actv_15_11_bits_nz(dat15_actv_nz[11]),
.io_dat_actv_15_11_bits_data(dat15_actv_data[95:88]),

.io_dat_actv_15_12_valid(dat15_actv_pvld[12]),
.io_dat_actv_15_12_bits_nz(dat15_actv_nz[12]),
.io_dat_actv_15_12_bits_data(dat15_actv_data[103:96]),

.io_dat_actv_15_13_valid(dat15_actv_pvld[13]),
.io_dat_actv_15_13_bits_nz(dat15_actv_nz[13]),
.io_dat_actv_15_13_bits_data(dat15_actv_data[111:104]),

.io_dat_actv_15_14_valid(dat15_actv_pvld[14]),
.io_dat_actv_15_14_bits_nz(dat15_actv_nz[14]),
.io_dat_actv_15_14_bits_data(dat15_actv_data[119:112]),

.io_dat_actv_15_15_valid(dat15_actv_pvld[15]),
.io_dat_actv_15_15_bits_nz(dat15_actv_nz[15]),
.io_dat_actv_15_15_bits_data(dat15_actv_data[127:120]),

.io_dat_actv_15_16_valid(dat15_actv_pvld[16]),
.io_dat_actv_15_16_bits_nz(dat15_actv_nz[16]),
.io_dat_actv_15_16_bits_data(dat15_actv_data[135:128]),

.io_dat_actv_15_17_valid(dat15_actv_pvld[17]),
.io_dat_actv_15_17_bits_nz(dat15_actv_nz[17]),
.io_dat_actv_15_17_bits_data(dat15_actv_data[143:136]),

.io_dat_actv_15_18_valid(dat15_actv_pvld[18]),
.io_dat_actv_15_18_bits_nz(dat15_actv_nz[18]),
.io_dat_actv_15_18_bits_data(dat15_actv_data[151:144]),

.io_dat_actv_15_19_valid(dat15_actv_pvld[19]),
.io_dat_actv_15_19_bits_nz(dat15_actv_nz[19]),
.io_dat_actv_15_19_bits_data(dat15_actv_data[159:152]),

.io_dat_actv_15_20_valid(dat15_actv_pvld[20]),
.io_dat_actv_15_20_bits_nz(dat15_actv_nz[20]),
.io_dat_actv_15_20_bits_data(dat15_actv_data[167:160]),

.io_dat_actv_15_21_valid(dat15_actv_pvld[21]),
.io_dat_actv_15_21_bits_nz(dat15_actv_nz[21]),
.io_dat_actv_15_21_bits_data(dat15_actv_data[175:168]),

.io_dat_actv_15_22_valid(dat15_actv_pvld[22]),
.io_dat_actv_15_22_bits_nz(dat15_actv_nz[22]),
.io_dat_actv_15_22_bits_data(dat15_actv_data[183:176]),

.io_dat_actv_15_23_valid(dat15_actv_pvld[23]),
.io_dat_actv_15_23_bits_nz(dat15_actv_nz[23]),
.io_dat_actv_15_23_bits_data(dat15_actv_data[191:184]),

.io_dat_actv_15_24_valid(dat15_actv_pvld[24]),
.io_dat_actv_15_24_bits_nz(dat15_actv_nz[24]),
.io_dat_actv_15_24_bits_data(dat15_actv_data[199:192]),

.io_dat_actv_15_25_valid(dat15_actv_pvld[25]),
.io_dat_actv_15_25_bits_nz(dat15_actv_nz[25]),
.io_dat_actv_15_25_bits_data(dat15_actv_data[207:200]),

.io_dat_actv_15_26_valid(dat15_actv_pvld[26]),
.io_dat_actv_15_26_bits_nz(dat15_actv_nz[26]),
.io_dat_actv_15_26_bits_data(dat15_actv_data[215:208]),

.io_dat_actv_15_27_valid(dat15_actv_pvld[27]),
.io_dat_actv_15_27_bits_nz(dat15_actv_nz[27]),
.io_dat_actv_15_27_bits_data(dat15_actv_data[223:216]),

.io_dat_actv_15_28_valid(dat15_actv_pvld[28]),
.io_dat_actv_15_28_bits_nz(dat15_actv_nz[28]),
.io_dat_actv_15_28_bits_data(dat15_actv_data[231:224]),

.io_dat_actv_15_29_valid(dat15_actv_pvld[29]),
.io_dat_actv_15_29_bits_nz(dat15_actv_nz[29]),
.io_dat_actv_15_29_bits_data(dat15_actv_data[239:232]),

.io_dat_actv_15_30_valid(dat15_actv_pvld[30]),
.io_dat_actv_15_30_bits_nz(dat15_actv_nz[30]),
.io_dat_actv_15_30_bits_data(dat15_actv_data[247:240]),

.io_dat_actv_15_31_valid(dat15_actv_pvld[31]),
.io_dat_actv_15_31_bits_nz(dat15_actv_nz[31]),
.io_dat_actv_15_31_bits_data(dat15_actv_data[255:248]),

.io_dat_actv_15_32_valid(dat15_actv_pvld[32]),
.io_dat_actv_15_32_bits_nz(dat15_actv_nz[32]),
.io_dat_actv_15_32_bits_data(dat15_actv_data[263:256]),

.io_dat_actv_15_33_valid(dat15_actv_pvld[33]),
.io_dat_actv_15_33_bits_nz(dat15_actv_nz[33]),
.io_dat_actv_15_33_bits_data(dat15_actv_data[271:264]),

.io_dat_actv_15_34_valid(dat15_actv_pvld[34]),
.io_dat_actv_15_34_bits_nz(dat15_actv_nz[34]),
.io_dat_actv_15_34_bits_data(dat15_actv_data[279:272]),

.io_dat_actv_15_35_valid(dat15_actv_pvld[35]),
.io_dat_actv_15_35_bits_nz(dat15_actv_nz[35]),
.io_dat_actv_15_35_bits_data(dat15_actv_data[287:280]),

.io_dat_actv_15_36_valid(dat15_actv_pvld[36]),
.io_dat_actv_15_36_bits_nz(dat15_actv_nz[36]),
.io_dat_actv_15_36_bits_data(dat15_actv_data[295:288]),

.io_dat_actv_15_37_valid(dat15_actv_pvld[37]),
.io_dat_actv_15_37_bits_nz(dat15_actv_nz[37]),
.io_dat_actv_15_37_bits_data(dat15_actv_data[303:296]),

.io_dat_actv_15_38_valid(dat15_actv_pvld[38]),
.io_dat_actv_15_38_bits_nz(dat15_actv_nz[38]),
.io_dat_actv_15_38_bits_data(dat15_actv_data[311:304]),

.io_dat_actv_15_39_valid(dat15_actv_pvld[39]),
.io_dat_actv_15_39_bits_nz(dat15_actv_nz[39]),
.io_dat_actv_15_39_bits_data(dat15_actv_data[319:312]),

.io_dat_actv_15_40_valid(dat15_actv_pvld[40]),
.io_dat_actv_15_40_bits_nz(dat15_actv_nz[40]),
.io_dat_actv_15_40_bits_data(dat15_actv_data[327:320]),

.io_dat_actv_15_41_valid(dat15_actv_pvld[41]),
.io_dat_actv_15_41_bits_nz(dat15_actv_nz[41]),
.io_dat_actv_15_41_bits_data(dat15_actv_data[335:328]),

.io_dat_actv_15_42_valid(dat15_actv_pvld[42]),
.io_dat_actv_15_42_bits_nz(dat15_actv_nz[42]),
.io_dat_actv_15_42_bits_data(dat15_actv_data[343:336]),

.io_dat_actv_15_43_valid(dat15_actv_pvld[43]),
.io_dat_actv_15_43_bits_nz(dat15_actv_nz[43]),
.io_dat_actv_15_43_bits_data(dat15_actv_data[351:344]),

.io_dat_actv_15_44_valid(dat15_actv_pvld[44]),
.io_dat_actv_15_44_bits_nz(dat15_actv_nz[44]),
.io_dat_actv_15_44_bits_data(dat15_actv_data[359:352]),

.io_dat_actv_15_45_valid(dat15_actv_pvld[45]),
.io_dat_actv_15_45_bits_nz(dat15_actv_nz[45]),
.io_dat_actv_15_45_bits_data(dat15_actv_data[367:360]),

.io_dat_actv_15_46_valid(dat15_actv_pvld[46]),
.io_dat_actv_15_46_bits_nz(dat15_actv_nz[46]),
.io_dat_actv_15_46_bits_data(dat15_actv_data[375:368]),

.io_dat_actv_15_47_valid(dat15_actv_pvld[47]),
.io_dat_actv_15_47_bits_nz(dat15_actv_nz[47]),
.io_dat_actv_15_47_bits_data(dat15_actv_data[383:376]),

.io_dat_actv_15_48_valid(dat15_actv_pvld[48]),
.io_dat_actv_15_48_bits_nz(dat15_actv_nz[48]),
.io_dat_actv_15_48_bits_data(dat15_actv_data[391:384]),

.io_dat_actv_15_49_valid(dat15_actv_pvld[49]),
.io_dat_actv_15_49_bits_nz(dat15_actv_nz[49]),
.io_dat_actv_15_49_bits_data(dat15_actv_data[399:392]),

.io_dat_actv_15_50_valid(dat15_actv_pvld[50]),
.io_dat_actv_15_50_bits_nz(dat15_actv_nz[50]),
.io_dat_actv_15_50_bits_data(dat15_actv_data[407:400]),

.io_dat_actv_15_51_valid(dat15_actv_pvld[51]),
.io_dat_actv_15_51_bits_nz(dat15_actv_nz[51]),
.io_dat_actv_15_51_bits_data(dat15_actv_data[415:408]),

.io_dat_actv_15_52_valid(dat15_actv_pvld[52]),
.io_dat_actv_15_52_bits_nz(dat15_actv_nz[52]),
.io_dat_actv_15_52_bits_data(dat15_actv_data[423:416]),

.io_dat_actv_15_53_valid(dat15_actv_pvld[53]),
.io_dat_actv_15_53_bits_nz(dat15_actv_nz[53]),
.io_dat_actv_15_53_bits_data(dat15_actv_data[431:424]),

.io_dat_actv_15_54_valid(dat15_actv_pvld[54]),
.io_dat_actv_15_54_bits_nz(dat15_actv_nz[54]),
.io_dat_actv_15_54_bits_data(dat15_actv_data[439:432]),

.io_dat_actv_15_55_valid(dat15_actv_pvld[55]),
.io_dat_actv_15_55_bits_nz(dat15_actv_nz[55]),
.io_dat_actv_15_55_bits_data(dat15_actv_data[447:440]),

.io_dat_actv_15_56_valid(dat15_actv_pvld[56]),
.io_dat_actv_15_56_bits_nz(dat15_actv_nz[56]),
.io_dat_actv_15_56_bits_data(dat15_actv_data[455:448]),

.io_dat_actv_15_57_valid(dat15_actv_pvld[57]),
.io_dat_actv_15_57_bits_nz(dat15_actv_nz[57]),
.io_dat_actv_15_57_bits_data(dat15_actv_data[463:456]),

.io_dat_actv_15_58_valid(dat15_actv_pvld[58]),
.io_dat_actv_15_58_bits_nz(dat15_actv_nz[58]),
.io_dat_actv_15_58_bits_data(dat15_actv_data[471:464]),

.io_dat_actv_15_59_valid(dat15_actv_pvld[59]),
.io_dat_actv_15_59_bits_nz(dat15_actv_nz[59]),
.io_dat_actv_15_59_bits_data(dat15_actv_data[479:472]),

.io_dat_actv_15_60_valid(dat15_actv_pvld[60]),
.io_dat_actv_15_60_bits_nz(dat15_actv_nz[60]),
.io_dat_actv_15_60_bits_data(dat15_actv_data[487:480]),

.io_dat_actv_15_61_valid(dat15_actv_pvld[61]),
.io_dat_actv_15_61_bits_nz(dat15_actv_nz[61]),
.io_dat_actv_15_61_bits_data(dat15_actv_data[495:488]),

.io_dat_actv_15_62_valid(dat15_actv_pvld[62]),
.io_dat_actv_15_62_bits_nz(dat15_actv_nz[62]),
.io_dat_actv_15_62_bits_data(dat15_actv_data[503:496]),

.io_dat_actv_15_63_valid(dat15_actv_pvld[63]),
.io_dat_actv_15_63_bits_nz(dat15_actv_nz[63]),
.io_dat_actv_15_63_bits_data(dat15_actv_data[511:504]),

    .io_wt_actv_0_0_valid(wt0_actv_pvld[0]),
.io_wt_actv_0_0_bits_nz(wt0_actv_nz[0]),
.io_wt_actv_0_0_bits_data(wt0_actv_data[7:0]),

.io_wt_actv_0_1_valid(wt0_actv_pvld[1]),
.io_wt_actv_0_1_bits_nz(wt0_actv_nz[1]),
.io_wt_actv_0_1_bits_data(wt0_actv_data[15:8]),

.io_wt_actv_0_2_valid(wt0_actv_pvld[2]),
.io_wt_actv_0_2_bits_nz(wt0_actv_nz[2]),
.io_wt_actv_0_2_bits_data(wt0_actv_data[23:16]),

.io_wt_actv_0_3_valid(wt0_actv_pvld[3]),
.io_wt_actv_0_3_bits_nz(wt0_actv_nz[3]),
.io_wt_actv_0_3_bits_data(wt0_actv_data[31:24]),

.io_wt_actv_0_4_valid(wt0_actv_pvld[4]),
.io_wt_actv_0_4_bits_nz(wt0_actv_nz[4]),
.io_wt_actv_0_4_bits_data(wt0_actv_data[39:32]),

.io_wt_actv_0_5_valid(wt0_actv_pvld[5]),
.io_wt_actv_0_5_bits_nz(wt0_actv_nz[5]),
.io_wt_actv_0_5_bits_data(wt0_actv_data[47:40]),

.io_wt_actv_0_6_valid(wt0_actv_pvld[6]),
.io_wt_actv_0_6_bits_nz(wt0_actv_nz[6]),
.io_wt_actv_0_6_bits_data(wt0_actv_data[55:48]),

.io_wt_actv_0_7_valid(wt0_actv_pvld[7]),
.io_wt_actv_0_7_bits_nz(wt0_actv_nz[7]),
.io_wt_actv_0_7_bits_data(wt0_actv_data[63:56]),

.io_wt_actv_0_8_valid(wt0_actv_pvld[8]),
.io_wt_actv_0_8_bits_nz(wt0_actv_nz[8]),
.io_wt_actv_0_8_bits_data(wt0_actv_data[71:64]),

.io_wt_actv_0_9_valid(wt0_actv_pvld[9]),
.io_wt_actv_0_9_bits_nz(wt0_actv_nz[9]),
.io_wt_actv_0_9_bits_data(wt0_actv_data[79:72]),

.io_wt_actv_0_10_valid(wt0_actv_pvld[10]),
.io_wt_actv_0_10_bits_nz(wt0_actv_nz[10]),
.io_wt_actv_0_10_bits_data(wt0_actv_data[87:80]),

.io_wt_actv_0_11_valid(wt0_actv_pvld[11]),
.io_wt_actv_0_11_bits_nz(wt0_actv_nz[11]),
.io_wt_actv_0_11_bits_data(wt0_actv_data[95:88]),

.io_wt_actv_0_12_valid(wt0_actv_pvld[12]),
.io_wt_actv_0_12_bits_nz(wt0_actv_nz[12]),
.io_wt_actv_0_12_bits_data(wt0_actv_data[103:96]),

.io_wt_actv_0_13_valid(wt0_actv_pvld[13]),
.io_wt_actv_0_13_bits_nz(wt0_actv_nz[13]),
.io_wt_actv_0_13_bits_data(wt0_actv_data[111:104]),

.io_wt_actv_0_14_valid(wt0_actv_pvld[14]),
.io_wt_actv_0_14_bits_nz(wt0_actv_nz[14]),
.io_wt_actv_0_14_bits_data(wt0_actv_data[119:112]),

.io_wt_actv_0_15_valid(wt0_actv_pvld[15]),
.io_wt_actv_0_15_bits_nz(wt0_actv_nz[15]),
.io_wt_actv_0_15_bits_data(wt0_actv_data[127:120]),

.io_wt_actv_0_16_valid(wt0_actv_pvld[16]),
.io_wt_actv_0_16_bits_nz(wt0_actv_nz[16]),
.io_wt_actv_0_16_bits_data(wt0_actv_data[135:128]),

.io_wt_actv_0_17_valid(wt0_actv_pvld[17]),
.io_wt_actv_0_17_bits_nz(wt0_actv_nz[17]),
.io_wt_actv_0_17_bits_data(wt0_actv_data[143:136]),

.io_wt_actv_0_18_valid(wt0_actv_pvld[18]),
.io_wt_actv_0_18_bits_nz(wt0_actv_nz[18]),
.io_wt_actv_0_18_bits_data(wt0_actv_data[151:144]),

.io_wt_actv_0_19_valid(wt0_actv_pvld[19]),
.io_wt_actv_0_19_bits_nz(wt0_actv_nz[19]),
.io_wt_actv_0_19_bits_data(wt0_actv_data[159:152]),

.io_wt_actv_0_20_valid(wt0_actv_pvld[20]),
.io_wt_actv_0_20_bits_nz(wt0_actv_nz[20]),
.io_wt_actv_0_20_bits_data(wt0_actv_data[167:160]),

.io_wt_actv_0_21_valid(wt0_actv_pvld[21]),
.io_wt_actv_0_21_bits_nz(wt0_actv_nz[21]),
.io_wt_actv_0_21_bits_data(wt0_actv_data[175:168]),

.io_wt_actv_0_22_valid(wt0_actv_pvld[22]),
.io_wt_actv_0_22_bits_nz(wt0_actv_nz[22]),
.io_wt_actv_0_22_bits_data(wt0_actv_data[183:176]),

.io_wt_actv_0_23_valid(wt0_actv_pvld[23]),
.io_wt_actv_0_23_bits_nz(wt0_actv_nz[23]),
.io_wt_actv_0_23_bits_data(wt0_actv_data[191:184]),

.io_wt_actv_0_24_valid(wt0_actv_pvld[24]),
.io_wt_actv_0_24_bits_nz(wt0_actv_nz[24]),
.io_wt_actv_0_24_bits_data(wt0_actv_data[199:192]),

.io_wt_actv_0_25_valid(wt0_actv_pvld[25]),
.io_wt_actv_0_25_bits_nz(wt0_actv_nz[25]),
.io_wt_actv_0_25_bits_data(wt0_actv_data[207:200]),

.io_wt_actv_0_26_valid(wt0_actv_pvld[26]),
.io_wt_actv_0_26_bits_nz(wt0_actv_nz[26]),
.io_wt_actv_0_26_bits_data(wt0_actv_data[215:208]),

.io_wt_actv_0_27_valid(wt0_actv_pvld[27]),
.io_wt_actv_0_27_bits_nz(wt0_actv_nz[27]),
.io_wt_actv_0_27_bits_data(wt0_actv_data[223:216]),

.io_wt_actv_0_28_valid(wt0_actv_pvld[28]),
.io_wt_actv_0_28_bits_nz(wt0_actv_nz[28]),
.io_wt_actv_0_28_bits_data(wt0_actv_data[231:224]),

.io_wt_actv_0_29_valid(wt0_actv_pvld[29]),
.io_wt_actv_0_29_bits_nz(wt0_actv_nz[29]),
.io_wt_actv_0_29_bits_data(wt0_actv_data[239:232]),

.io_wt_actv_0_30_valid(wt0_actv_pvld[30]),
.io_wt_actv_0_30_bits_nz(wt0_actv_nz[30]),
.io_wt_actv_0_30_bits_data(wt0_actv_data[247:240]),

.io_wt_actv_0_31_valid(wt0_actv_pvld[31]),
.io_wt_actv_0_31_bits_nz(wt0_actv_nz[31]),
.io_wt_actv_0_31_bits_data(wt0_actv_data[255:248]),

.io_wt_actv_0_32_valid(wt0_actv_pvld[32]),
.io_wt_actv_0_32_bits_nz(wt0_actv_nz[32]),
.io_wt_actv_0_32_bits_data(wt0_actv_data[263:256]),

.io_wt_actv_0_33_valid(wt0_actv_pvld[33]),
.io_wt_actv_0_33_bits_nz(wt0_actv_nz[33]),
.io_wt_actv_0_33_bits_data(wt0_actv_data[271:264]),

.io_wt_actv_0_34_valid(wt0_actv_pvld[34]),
.io_wt_actv_0_34_bits_nz(wt0_actv_nz[34]),
.io_wt_actv_0_34_bits_data(wt0_actv_data[279:272]),

.io_wt_actv_0_35_valid(wt0_actv_pvld[35]),
.io_wt_actv_0_35_bits_nz(wt0_actv_nz[35]),
.io_wt_actv_0_35_bits_data(wt0_actv_data[287:280]),

.io_wt_actv_0_36_valid(wt0_actv_pvld[36]),
.io_wt_actv_0_36_bits_nz(wt0_actv_nz[36]),
.io_wt_actv_0_36_bits_data(wt0_actv_data[295:288]),

.io_wt_actv_0_37_valid(wt0_actv_pvld[37]),
.io_wt_actv_0_37_bits_nz(wt0_actv_nz[37]),
.io_wt_actv_0_37_bits_data(wt0_actv_data[303:296]),

.io_wt_actv_0_38_valid(wt0_actv_pvld[38]),
.io_wt_actv_0_38_bits_nz(wt0_actv_nz[38]),
.io_wt_actv_0_38_bits_data(wt0_actv_data[311:304]),

.io_wt_actv_0_39_valid(wt0_actv_pvld[39]),
.io_wt_actv_0_39_bits_nz(wt0_actv_nz[39]),
.io_wt_actv_0_39_bits_data(wt0_actv_data[319:312]),

.io_wt_actv_0_40_valid(wt0_actv_pvld[40]),
.io_wt_actv_0_40_bits_nz(wt0_actv_nz[40]),
.io_wt_actv_0_40_bits_data(wt0_actv_data[327:320]),

.io_wt_actv_0_41_valid(wt0_actv_pvld[41]),
.io_wt_actv_0_41_bits_nz(wt0_actv_nz[41]),
.io_wt_actv_0_41_bits_data(wt0_actv_data[335:328]),

.io_wt_actv_0_42_valid(wt0_actv_pvld[42]),
.io_wt_actv_0_42_bits_nz(wt0_actv_nz[42]),
.io_wt_actv_0_42_bits_data(wt0_actv_data[343:336]),

.io_wt_actv_0_43_valid(wt0_actv_pvld[43]),
.io_wt_actv_0_43_bits_nz(wt0_actv_nz[43]),
.io_wt_actv_0_43_bits_data(wt0_actv_data[351:344]),

.io_wt_actv_0_44_valid(wt0_actv_pvld[44]),
.io_wt_actv_0_44_bits_nz(wt0_actv_nz[44]),
.io_wt_actv_0_44_bits_data(wt0_actv_data[359:352]),

.io_wt_actv_0_45_valid(wt0_actv_pvld[45]),
.io_wt_actv_0_45_bits_nz(wt0_actv_nz[45]),
.io_wt_actv_0_45_bits_data(wt0_actv_data[367:360]),

.io_wt_actv_0_46_valid(wt0_actv_pvld[46]),
.io_wt_actv_0_46_bits_nz(wt0_actv_nz[46]),
.io_wt_actv_0_46_bits_data(wt0_actv_data[375:368]),

.io_wt_actv_0_47_valid(wt0_actv_pvld[47]),
.io_wt_actv_0_47_bits_nz(wt0_actv_nz[47]),
.io_wt_actv_0_47_bits_data(wt0_actv_data[383:376]),

.io_wt_actv_0_48_valid(wt0_actv_pvld[48]),
.io_wt_actv_0_48_bits_nz(wt0_actv_nz[48]),
.io_wt_actv_0_48_bits_data(wt0_actv_data[391:384]),

.io_wt_actv_0_49_valid(wt0_actv_pvld[49]),
.io_wt_actv_0_49_bits_nz(wt0_actv_nz[49]),
.io_wt_actv_0_49_bits_data(wt0_actv_data[399:392]),

.io_wt_actv_0_50_valid(wt0_actv_pvld[50]),
.io_wt_actv_0_50_bits_nz(wt0_actv_nz[50]),
.io_wt_actv_0_50_bits_data(wt0_actv_data[407:400]),

.io_wt_actv_0_51_valid(wt0_actv_pvld[51]),
.io_wt_actv_0_51_bits_nz(wt0_actv_nz[51]),
.io_wt_actv_0_51_bits_data(wt0_actv_data[415:408]),

.io_wt_actv_0_52_valid(wt0_actv_pvld[52]),
.io_wt_actv_0_52_bits_nz(wt0_actv_nz[52]),
.io_wt_actv_0_52_bits_data(wt0_actv_data[423:416]),

.io_wt_actv_0_53_valid(wt0_actv_pvld[53]),
.io_wt_actv_0_53_bits_nz(wt0_actv_nz[53]),
.io_wt_actv_0_53_bits_data(wt0_actv_data[431:424]),

.io_wt_actv_0_54_valid(wt0_actv_pvld[54]),
.io_wt_actv_0_54_bits_nz(wt0_actv_nz[54]),
.io_wt_actv_0_54_bits_data(wt0_actv_data[439:432]),

.io_wt_actv_0_55_valid(wt0_actv_pvld[55]),
.io_wt_actv_0_55_bits_nz(wt0_actv_nz[55]),
.io_wt_actv_0_55_bits_data(wt0_actv_data[447:440]),

.io_wt_actv_0_56_valid(wt0_actv_pvld[56]),
.io_wt_actv_0_56_bits_nz(wt0_actv_nz[56]),
.io_wt_actv_0_56_bits_data(wt0_actv_data[455:448]),

.io_wt_actv_0_57_valid(wt0_actv_pvld[57]),
.io_wt_actv_0_57_bits_nz(wt0_actv_nz[57]),
.io_wt_actv_0_57_bits_data(wt0_actv_data[463:456]),

.io_wt_actv_0_58_valid(wt0_actv_pvld[58]),
.io_wt_actv_0_58_bits_nz(wt0_actv_nz[58]),
.io_wt_actv_0_58_bits_data(wt0_actv_data[471:464]),

.io_wt_actv_0_59_valid(wt0_actv_pvld[59]),
.io_wt_actv_0_59_bits_nz(wt0_actv_nz[59]),
.io_wt_actv_0_59_bits_data(wt0_actv_data[479:472]),

.io_wt_actv_0_60_valid(wt0_actv_pvld[60]),
.io_wt_actv_0_60_bits_nz(wt0_actv_nz[60]),
.io_wt_actv_0_60_bits_data(wt0_actv_data[487:480]),

.io_wt_actv_0_61_valid(wt0_actv_pvld[61]),
.io_wt_actv_0_61_bits_nz(wt0_actv_nz[61]),
.io_wt_actv_0_61_bits_data(wt0_actv_data[495:488]),

.io_wt_actv_0_62_valid(wt0_actv_pvld[62]),
.io_wt_actv_0_62_bits_nz(wt0_actv_nz[62]),
.io_wt_actv_0_62_bits_data(wt0_actv_data[503:496]),

.io_wt_actv_0_63_valid(wt0_actv_pvld[63]),
.io_wt_actv_0_63_bits_nz(wt0_actv_nz[63]),
.io_wt_actv_0_63_bits_data(wt0_actv_data[511:504]),

.io_wt_actv_1_0_valid(wt1_actv_pvld[0]),
.io_wt_actv_1_0_bits_nz(wt1_actv_nz[0]),
.io_wt_actv_1_0_bits_data(wt1_actv_data[7:0]),

.io_wt_actv_1_1_valid(wt1_actv_pvld[1]),
.io_wt_actv_1_1_bits_nz(wt1_actv_nz[1]),
.io_wt_actv_1_1_bits_data(wt1_actv_data[15:8]),

.io_wt_actv_1_2_valid(wt1_actv_pvld[2]),
.io_wt_actv_1_2_bits_nz(wt1_actv_nz[2]),
.io_wt_actv_1_2_bits_data(wt1_actv_data[23:16]),

.io_wt_actv_1_3_valid(wt1_actv_pvld[3]),
.io_wt_actv_1_3_bits_nz(wt1_actv_nz[3]),
.io_wt_actv_1_3_bits_data(wt1_actv_data[31:24]),

.io_wt_actv_1_4_valid(wt1_actv_pvld[4]),
.io_wt_actv_1_4_bits_nz(wt1_actv_nz[4]),
.io_wt_actv_1_4_bits_data(wt1_actv_data[39:32]),

.io_wt_actv_1_5_valid(wt1_actv_pvld[5]),
.io_wt_actv_1_5_bits_nz(wt1_actv_nz[5]),
.io_wt_actv_1_5_bits_data(wt1_actv_data[47:40]),

.io_wt_actv_1_6_valid(wt1_actv_pvld[6]),
.io_wt_actv_1_6_bits_nz(wt1_actv_nz[6]),
.io_wt_actv_1_6_bits_data(wt1_actv_data[55:48]),

.io_wt_actv_1_7_valid(wt1_actv_pvld[7]),
.io_wt_actv_1_7_bits_nz(wt1_actv_nz[7]),
.io_wt_actv_1_7_bits_data(wt1_actv_data[63:56]),

.io_wt_actv_1_8_valid(wt1_actv_pvld[8]),
.io_wt_actv_1_8_bits_nz(wt1_actv_nz[8]),
.io_wt_actv_1_8_bits_data(wt1_actv_data[71:64]),

.io_wt_actv_1_9_valid(wt1_actv_pvld[9]),
.io_wt_actv_1_9_bits_nz(wt1_actv_nz[9]),
.io_wt_actv_1_9_bits_data(wt1_actv_data[79:72]),

.io_wt_actv_1_10_valid(wt1_actv_pvld[10]),
.io_wt_actv_1_10_bits_nz(wt1_actv_nz[10]),
.io_wt_actv_1_10_bits_data(wt1_actv_data[87:80]),

.io_wt_actv_1_11_valid(wt1_actv_pvld[11]),
.io_wt_actv_1_11_bits_nz(wt1_actv_nz[11]),
.io_wt_actv_1_11_bits_data(wt1_actv_data[95:88]),

.io_wt_actv_1_12_valid(wt1_actv_pvld[12]),
.io_wt_actv_1_12_bits_nz(wt1_actv_nz[12]),
.io_wt_actv_1_12_bits_data(wt1_actv_data[103:96]),

.io_wt_actv_1_13_valid(wt1_actv_pvld[13]),
.io_wt_actv_1_13_bits_nz(wt1_actv_nz[13]),
.io_wt_actv_1_13_bits_data(wt1_actv_data[111:104]),

.io_wt_actv_1_14_valid(wt1_actv_pvld[14]),
.io_wt_actv_1_14_bits_nz(wt1_actv_nz[14]),
.io_wt_actv_1_14_bits_data(wt1_actv_data[119:112]),

.io_wt_actv_1_15_valid(wt1_actv_pvld[15]),
.io_wt_actv_1_15_bits_nz(wt1_actv_nz[15]),
.io_wt_actv_1_15_bits_data(wt1_actv_data[127:120]),

.io_wt_actv_1_16_valid(wt1_actv_pvld[16]),
.io_wt_actv_1_16_bits_nz(wt1_actv_nz[16]),
.io_wt_actv_1_16_bits_data(wt1_actv_data[135:128]),

.io_wt_actv_1_17_valid(wt1_actv_pvld[17]),
.io_wt_actv_1_17_bits_nz(wt1_actv_nz[17]),
.io_wt_actv_1_17_bits_data(wt1_actv_data[143:136]),

.io_wt_actv_1_18_valid(wt1_actv_pvld[18]),
.io_wt_actv_1_18_bits_nz(wt1_actv_nz[18]),
.io_wt_actv_1_18_bits_data(wt1_actv_data[151:144]),

.io_wt_actv_1_19_valid(wt1_actv_pvld[19]),
.io_wt_actv_1_19_bits_nz(wt1_actv_nz[19]),
.io_wt_actv_1_19_bits_data(wt1_actv_data[159:152]),

.io_wt_actv_1_20_valid(wt1_actv_pvld[20]),
.io_wt_actv_1_20_bits_nz(wt1_actv_nz[20]),
.io_wt_actv_1_20_bits_data(wt1_actv_data[167:160]),

.io_wt_actv_1_21_valid(wt1_actv_pvld[21]),
.io_wt_actv_1_21_bits_nz(wt1_actv_nz[21]),
.io_wt_actv_1_21_bits_data(wt1_actv_data[175:168]),

.io_wt_actv_1_22_valid(wt1_actv_pvld[22]),
.io_wt_actv_1_22_bits_nz(wt1_actv_nz[22]),
.io_wt_actv_1_22_bits_data(wt1_actv_data[183:176]),

.io_wt_actv_1_23_valid(wt1_actv_pvld[23]),
.io_wt_actv_1_23_bits_nz(wt1_actv_nz[23]),
.io_wt_actv_1_23_bits_data(wt1_actv_data[191:184]),

.io_wt_actv_1_24_valid(wt1_actv_pvld[24]),
.io_wt_actv_1_24_bits_nz(wt1_actv_nz[24]),
.io_wt_actv_1_24_bits_data(wt1_actv_data[199:192]),

.io_wt_actv_1_25_valid(wt1_actv_pvld[25]),
.io_wt_actv_1_25_bits_nz(wt1_actv_nz[25]),
.io_wt_actv_1_25_bits_data(wt1_actv_data[207:200]),

.io_wt_actv_1_26_valid(wt1_actv_pvld[26]),
.io_wt_actv_1_26_bits_nz(wt1_actv_nz[26]),
.io_wt_actv_1_26_bits_data(wt1_actv_data[215:208]),

.io_wt_actv_1_27_valid(wt1_actv_pvld[27]),
.io_wt_actv_1_27_bits_nz(wt1_actv_nz[27]),
.io_wt_actv_1_27_bits_data(wt1_actv_data[223:216]),

.io_wt_actv_1_28_valid(wt1_actv_pvld[28]),
.io_wt_actv_1_28_bits_nz(wt1_actv_nz[28]),
.io_wt_actv_1_28_bits_data(wt1_actv_data[231:224]),

.io_wt_actv_1_29_valid(wt1_actv_pvld[29]),
.io_wt_actv_1_29_bits_nz(wt1_actv_nz[29]),
.io_wt_actv_1_29_bits_data(wt1_actv_data[239:232]),

.io_wt_actv_1_30_valid(wt1_actv_pvld[30]),
.io_wt_actv_1_30_bits_nz(wt1_actv_nz[30]),
.io_wt_actv_1_30_bits_data(wt1_actv_data[247:240]),

.io_wt_actv_1_31_valid(wt1_actv_pvld[31]),
.io_wt_actv_1_31_bits_nz(wt1_actv_nz[31]),
.io_wt_actv_1_31_bits_data(wt1_actv_data[255:248]),

.io_wt_actv_1_32_valid(wt1_actv_pvld[32]),
.io_wt_actv_1_32_bits_nz(wt1_actv_nz[32]),
.io_wt_actv_1_32_bits_data(wt1_actv_data[263:256]),

.io_wt_actv_1_33_valid(wt1_actv_pvld[33]),
.io_wt_actv_1_33_bits_nz(wt1_actv_nz[33]),
.io_wt_actv_1_33_bits_data(wt1_actv_data[271:264]),

.io_wt_actv_1_34_valid(wt1_actv_pvld[34]),
.io_wt_actv_1_34_bits_nz(wt1_actv_nz[34]),
.io_wt_actv_1_34_bits_data(wt1_actv_data[279:272]),

.io_wt_actv_1_35_valid(wt1_actv_pvld[35]),
.io_wt_actv_1_35_bits_nz(wt1_actv_nz[35]),
.io_wt_actv_1_35_bits_data(wt1_actv_data[287:280]),

.io_wt_actv_1_36_valid(wt1_actv_pvld[36]),
.io_wt_actv_1_36_bits_nz(wt1_actv_nz[36]),
.io_wt_actv_1_36_bits_data(wt1_actv_data[295:288]),

.io_wt_actv_1_37_valid(wt1_actv_pvld[37]),
.io_wt_actv_1_37_bits_nz(wt1_actv_nz[37]),
.io_wt_actv_1_37_bits_data(wt1_actv_data[303:296]),

.io_wt_actv_1_38_valid(wt1_actv_pvld[38]),
.io_wt_actv_1_38_bits_nz(wt1_actv_nz[38]),
.io_wt_actv_1_38_bits_data(wt1_actv_data[311:304]),

.io_wt_actv_1_39_valid(wt1_actv_pvld[39]),
.io_wt_actv_1_39_bits_nz(wt1_actv_nz[39]),
.io_wt_actv_1_39_bits_data(wt1_actv_data[319:312]),

.io_wt_actv_1_40_valid(wt1_actv_pvld[40]),
.io_wt_actv_1_40_bits_nz(wt1_actv_nz[40]),
.io_wt_actv_1_40_bits_data(wt1_actv_data[327:320]),

.io_wt_actv_1_41_valid(wt1_actv_pvld[41]),
.io_wt_actv_1_41_bits_nz(wt1_actv_nz[41]),
.io_wt_actv_1_41_bits_data(wt1_actv_data[335:328]),

.io_wt_actv_1_42_valid(wt1_actv_pvld[42]),
.io_wt_actv_1_42_bits_nz(wt1_actv_nz[42]),
.io_wt_actv_1_42_bits_data(wt1_actv_data[343:336]),

.io_wt_actv_1_43_valid(wt1_actv_pvld[43]),
.io_wt_actv_1_43_bits_nz(wt1_actv_nz[43]),
.io_wt_actv_1_43_bits_data(wt1_actv_data[351:344]),

.io_wt_actv_1_44_valid(wt1_actv_pvld[44]),
.io_wt_actv_1_44_bits_nz(wt1_actv_nz[44]),
.io_wt_actv_1_44_bits_data(wt1_actv_data[359:352]),

.io_wt_actv_1_45_valid(wt1_actv_pvld[45]),
.io_wt_actv_1_45_bits_nz(wt1_actv_nz[45]),
.io_wt_actv_1_45_bits_data(wt1_actv_data[367:360]),

.io_wt_actv_1_46_valid(wt1_actv_pvld[46]),
.io_wt_actv_1_46_bits_nz(wt1_actv_nz[46]),
.io_wt_actv_1_46_bits_data(wt1_actv_data[375:368]),

.io_wt_actv_1_47_valid(wt1_actv_pvld[47]),
.io_wt_actv_1_47_bits_nz(wt1_actv_nz[47]),
.io_wt_actv_1_47_bits_data(wt1_actv_data[383:376]),

.io_wt_actv_1_48_valid(wt1_actv_pvld[48]),
.io_wt_actv_1_48_bits_nz(wt1_actv_nz[48]),
.io_wt_actv_1_48_bits_data(wt1_actv_data[391:384]),

.io_wt_actv_1_49_valid(wt1_actv_pvld[49]),
.io_wt_actv_1_49_bits_nz(wt1_actv_nz[49]),
.io_wt_actv_1_49_bits_data(wt1_actv_data[399:392]),

.io_wt_actv_1_50_valid(wt1_actv_pvld[50]),
.io_wt_actv_1_50_bits_nz(wt1_actv_nz[50]),
.io_wt_actv_1_50_bits_data(wt1_actv_data[407:400]),

.io_wt_actv_1_51_valid(wt1_actv_pvld[51]),
.io_wt_actv_1_51_bits_nz(wt1_actv_nz[51]),
.io_wt_actv_1_51_bits_data(wt1_actv_data[415:408]),

.io_wt_actv_1_52_valid(wt1_actv_pvld[52]),
.io_wt_actv_1_52_bits_nz(wt1_actv_nz[52]),
.io_wt_actv_1_52_bits_data(wt1_actv_data[423:416]),

.io_wt_actv_1_53_valid(wt1_actv_pvld[53]),
.io_wt_actv_1_53_bits_nz(wt1_actv_nz[53]),
.io_wt_actv_1_53_bits_data(wt1_actv_data[431:424]),

.io_wt_actv_1_54_valid(wt1_actv_pvld[54]),
.io_wt_actv_1_54_bits_nz(wt1_actv_nz[54]),
.io_wt_actv_1_54_bits_data(wt1_actv_data[439:432]),

.io_wt_actv_1_55_valid(wt1_actv_pvld[55]),
.io_wt_actv_1_55_bits_nz(wt1_actv_nz[55]),
.io_wt_actv_1_55_bits_data(wt1_actv_data[447:440]),

.io_wt_actv_1_56_valid(wt1_actv_pvld[56]),
.io_wt_actv_1_56_bits_nz(wt1_actv_nz[56]),
.io_wt_actv_1_56_bits_data(wt1_actv_data[455:448]),

.io_wt_actv_1_57_valid(wt1_actv_pvld[57]),
.io_wt_actv_1_57_bits_nz(wt1_actv_nz[57]),
.io_wt_actv_1_57_bits_data(wt1_actv_data[463:456]),

.io_wt_actv_1_58_valid(wt1_actv_pvld[58]),
.io_wt_actv_1_58_bits_nz(wt1_actv_nz[58]),
.io_wt_actv_1_58_bits_data(wt1_actv_data[471:464]),

.io_wt_actv_1_59_valid(wt1_actv_pvld[59]),
.io_wt_actv_1_59_bits_nz(wt1_actv_nz[59]),
.io_wt_actv_1_59_bits_data(wt1_actv_data[479:472]),

.io_wt_actv_1_60_valid(wt1_actv_pvld[60]),
.io_wt_actv_1_60_bits_nz(wt1_actv_nz[60]),
.io_wt_actv_1_60_bits_data(wt1_actv_data[487:480]),

.io_wt_actv_1_61_valid(wt1_actv_pvld[61]),
.io_wt_actv_1_61_bits_nz(wt1_actv_nz[61]),
.io_wt_actv_1_61_bits_data(wt1_actv_data[495:488]),

.io_wt_actv_1_62_valid(wt1_actv_pvld[62]),
.io_wt_actv_1_62_bits_nz(wt1_actv_nz[62]),
.io_wt_actv_1_62_bits_data(wt1_actv_data[503:496]),

.io_wt_actv_1_63_valid(wt1_actv_pvld[63]),
.io_wt_actv_1_63_bits_nz(wt1_actv_nz[63]),
.io_wt_actv_1_63_bits_data(wt1_actv_data[511:504]),

.io_wt_actv_2_0_valid(wt2_actv_pvld[0]),
.io_wt_actv_2_0_bits_nz(wt2_actv_nz[0]),
.io_wt_actv_2_0_bits_data(wt2_actv_data[7:0]),

.io_wt_actv_2_1_valid(wt2_actv_pvld[1]),
.io_wt_actv_2_1_bits_nz(wt2_actv_nz[1]),
.io_wt_actv_2_1_bits_data(wt2_actv_data[15:8]),

.io_wt_actv_2_2_valid(wt2_actv_pvld[2]),
.io_wt_actv_2_2_bits_nz(wt2_actv_nz[2]),
.io_wt_actv_2_2_bits_data(wt2_actv_data[23:16]),

.io_wt_actv_2_3_valid(wt2_actv_pvld[3]),
.io_wt_actv_2_3_bits_nz(wt2_actv_nz[3]),
.io_wt_actv_2_3_bits_data(wt2_actv_data[31:24]),

.io_wt_actv_2_4_valid(wt2_actv_pvld[4]),
.io_wt_actv_2_4_bits_nz(wt2_actv_nz[4]),
.io_wt_actv_2_4_bits_data(wt2_actv_data[39:32]),

.io_wt_actv_2_5_valid(wt2_actv_pvld[5]),
.io_wt_actv_2_5_bits_nz(wt2_actv_nz[5]),
.io_wt_actv_2_5_bits_data(wt2_actv_data[47:40]),

.io_wt_actv_2_6_valid(wt2_actv_pvld[6]),
.io_wt_actv_2_6_bits_nz(wt2_actv_nz[6]),
.io_wt_actv_2_6_bits_data(wt2_actv_data[55:48]),

.io_wt_actv_2_7_valid(wt2_actv_pvld[7]),
.io_wt_actv_2_7_bits_nz(wt2_actv_nz[7]),
.io_wt_actv_2_7_bits_data(wt2_actv_data[63:56]),

.io_wt_actv_2_8_valid(wt2_actv_pvld[8]),
.io_wt_actv_2_8_bits_nz(wt2_actv_nz[8]),
.io_wt_actv_2_8_bits_data(wt2_actv_data[71:64]),

.io_wt_actv_2_9_valid(wt2_actv_pvld[9]),
.io_wt_actv_2_9_bits_nz(wt2_actv_nz[9]),
.io_wt_actv_2_9_bits_data(wt2_actv_data[79:72]),

.io_wt_actv_2_10_valid(wt2_actv_pvld[10]),
.io_wt_actv_2_10_bits_nz(wt2_actv_nz[10]),
.io_wt_actv_2_10_bits_data(wt2_actv_data[87:80]),

.io_wt_actv_2_11_valid(wt2_actv_pvld[11]),
.io_wt_actv_2_11_bits_nz(wt2_actv_nz[11]),
.io_wt_actv_2_11_bits_data(wt2_actv_data[95:88]),

.io_wt_actv_2_12_valid(wt2_actv_pvld[12]),
.io_wt_actv_2_12_bits_nz(wt2_actv_nz[12]),
.io_wt_actv_2_12_bits_data(wt2_actv_data[103:96]),

.io_wt_actv_2_13_valid(wt2_actv_pvld[13]),
.io_wt_actv_2_13_bits_nz(wt2_actv_nz[13]),
.io_wt_actv_2_13_bits_data(wt2_actv_data[111:104]),

.io_wt_actv_2_14_valid(wt2_actv_pvld[14]),
.io_wt_actv_2_14_bits_nz(wt2_actv_nz[14]),
.io_wt_actv_2_14_bits_data(wt2_actv_data[119:112]),

.io_wt_actv_2_15_valid(wt2_actv_pvld[15]),
.io_wt_actv_2_15_bits_nz(wt2_actv_nz[15]),
.io_wt_actv_2_15_bits_data(wt2_actv_data[127:120]),

.io_wt_actv_2_16_valid(wt2_actv_pvld[16]),
.io_wt_actv_2_16_bits_nz(wt2_actv_nz[16]),
.io_wt_actv_2_16_bits_data(wt2_actv_data[135:128]),

.io_wt_actv_2_17_valid(wt2_actv_pvld[17]),
.io_wt_actv_2_17_bits_nz(wt2_actv_nz[17]),
.io_wt_actv_2_17_bits_data(wt2_actv_data[143:136]),

.io_wt_actv_2_18_valid(wt2_actv_pvld[18]),
.io_wt_actv_2_18_bits_nz(wt2_actv_nz[18]),
.io_wt_actv_2_18_bits_data(wt2_actv_data[151:144]),

.io_wt_actv_2_19_valid(wt2_actv_pvld[19]),
.io_wt_actv_2_19_bits_nz(wt2_actv_nz[19]),
.io_wt_actv_2_19_bits_data(wt2_actv_data[159:152]),

.io_wt_actv_2_20_valid(wt2_actv_pvld[20]),
.io_wt_actv_2_20_bits_nz(wt2_actv_nz[20]),
.io_wt_actv_2_20_bits_data(wt2_actv_data[167:160]),

.io_wt_actv_2_21_valid(wt2_actv_pvld[21]),
.io_wt_actv_2_21_bits_nz(wt2_actv_nz[21]),
.io_wt_actv_2_21_bits_data(wt2_actv_data[175:168]),

.io_wt_actv_2_22_valid(wt2_actv_pvld[22]),
.io_wt_actv_2_22_bits_nz(wt2_actv_nz[22]),
.io_wt_actv_2_22_bits_data(wt2_actv_data[183:176]),

.io_wt_actv_2_23_valid(wt2_actv_pvld[23]),
.io_wt_actv_2_23_bits_nz(wt2_actv_nz[23]),
.io_wt_actv_2_23_bits_data(wt2_actv_data[191:184]),

.io_wt_actv_2_24_valid(wt2_actv_pvld[24]),
.io_wt_actv_2_24_bits_nz(wt2_actv_nz[24]),
.io_wt_actv_2_24_bits_data(wt2_actv_data[199:192]),

.io_wt_actv_2_25_valid(wt2_actv_pvld[25]),
.io_wt_actv_2_25_bits_nz(wt2_actv_nz[25]),
.io_wt_actv_2_25_bits_data(wt2_actv_data[207:200]),

.io_wt_actv_2_26_valid(wt2_actv_pvld[26]),
.io_wt_actv_2_26_bits_nz(wt2_actv_nz[26]),
.io_wt_actv_2_26_bits_data(wt2_actv_data[215:208]),

.io_wt_actv_2_27_valid(wt2_actv_pvld[27]),
.io_wt_actv_2_27_bits_nz(wt2_actv_nz[27]),
.io_wt_actv_2_27_bits_data(wt2_actv_data[223:216]),

.io_wt_actv_2_28_valid(wt2_actv_pvld[28]),
.io_wt_actv_2_28_bits_nz(wt2_actv_nz[28]),
.io_wt_actv_2_28_bits_data(wt2_actv_data[231:224]),

.io_wt_actv_2_29_valid(wt2_actv_pvld[29]),
.io_wt_actv_2_29_bits_nz(wt2_actv_nz[29]),
.io_wt_actv_2_29_bits_data(wt2_actv_data[239:232]),

.io_wt_actv_2_30_valid(wt2_actv_pvld[30]),
.io_wt_actv_2_30_bits_nz(wt2_actv_nz[30]),
.io_wt_actv_2_30_bits_data(wt2_actv_data[247:240]),

.io_wt_actv_2_31_valid(wt2_actv_pvld[31]),
.io_wt_actv_2_31_bits_nz(wt2_actv_nz[31]),
.io_wt_actv_2_31_bits_data(wt2_actv_data[255:248]),

.io_wt_actv_2_32_valid(wt2_actv_pvld[32]),
.io_wt_actv_2_32_bits_nz(wt2_actv_nz[32]),
.io_wt_actv_2_32_bits_data(wt2_actv_data[263:256]),

.io_wt_actv_2_33_valid(wt2_actv_pvld[33]),
.io_wt_actv_2_33_bits_nz(wt2_actv_nz[33]),
.io_wt_actv_2_33_bits_data(wt2_actv_data[271:264]),

.io_wt_actv_2_34_valid(wt2_actv_pvld[34]),
.io_wt_actv_2_34_bits_nz(wt2_actv_nz[34]),
.io_wt_actv_2_34_bits_data(wt2_actv_data[279:272]),

.io_wt_actv_2_35_valid(wt2_actv_pvld[35]),
.io_wt_actv_2_35_bits_nz(wt2_actv_nz[35]),
.io_wt_actv_2_35_bits_data(wt2_actv_data[287:280]),

.io_wt_actv_2_36_valid(wt2_actv_pvld[36]),
.io_wt_actv_2_36_bits_nz(wt2_actv_nz[36]),
.io_wt_actv_2_36_bits_data(wt2_actv_data[295:288]),

.io_wt_actv_2_37_valid(wt2_actv_pvld[37]),
.io_wt_actv_2_37_bits_nz(wt2_actv_nz[37]),
.io_wt_actv_2_37_bits_data(wt2_actv_data[303:296]),

.io_wt_actv_2_38_valid(wt2_actv_pvld[38]),
.io_wt_actv_2_38_bits_nz(wt2_actv_nz[38]),
.io_wt_actv_2_38_bits_data(wt2_actv_data[311:304]),

.io_wt_actv_2_39_valid(wt2_actv_pvld[39]),
.io_wt_actv_2_39_bits_nz(wt2_actv_nz[39]),
.io_wt_actv_2_39_bits_data(wt2_actv_data[319:312]),

.io_wt_actv_2_40_valid(wt2_actv_pvld[40]),
.io_wt_actv_2_40_bits_nz(wt2_actv_nz[40]),
.io_wt_actv_2_40_bits_data(wt2_actv_data[327:320]),

.io_wt_actv_2_41_valid(wt2_actv_pvld[41]),
.io_wt_actv_2_41_bits_nz(wt2_actv_nz[41]),
.io_wt_actv_2_41_bits_data(wt2_actv_data[335:328]),

.io_wt_actv_2_42_valid(wt2_actv_pvld[42]),
.io_wt_actv_2_42_bits_nz(wt2_actv_nz[42]),
.io_wt_actv_2_42_bits_data(wt2_actv_data[343:336]),

.io_wt_actv_2_43_valid(wt2_actv_pvld[43]),
.io_wt_actv_2_43_bits_nz(wt2_actv_nz[43]),
.io_wt_actv_2_43_bits_data(wt2_actv_data[351:344]),

.io_wt_actv_2_44_valid(wt2_actv_pvld[44]),
.io_wt_actv_2_44_bits_nz(wt2_actv_nz[44]),
.io_wt_actv_2_44_bits_data(wt2_actv_data[359:352]),

.io_wt_actv_2_45_valid(wt2_actv_pvld[45]),
.io_wt_actv_2_45_bits_nz(wt2_actv_nz[45]),
.io_wt_actv_2_45_bits_data(wt2_actv_data[367:360]),

.io_wt_actv_2_46_valid(wt2_actv_pvld[46]),
.io_wt_actv_2_46_bits_nz(wt2_actv_nz[46]),
.io_wt_actv_2_46_bits_data(wt2_actv_data[375:368]),

.io_wt_actv_2_47_valid(wt2_actv_pvld[47]),
.io_wt_actv_2_47_bits_nz(wt2_actv_nz[47]),
.io_wt_actv_2_47_bits_data(wt2_actv_data[383:376]),

.io_wt_actv_2_48_valid(wt2_actv_pvld[48]),
.io_wt_actv_2_48_bits_nz(wt2_actv_nz[48]),
.io_wt_actv_2_48_bits_data(wt2_actv_data[391:384]),

.io_wt_actv_2_49_valid(wt2_actv_pvld[49]),
.io_wt_actv_2_49_bits_nz(wt2_actv_nz[49]),
.io_wt_actv_2_49_bits_data(wt2_actv_data[399:392]),

.io_wt_actv_2_50_valid(wt2_actv_pvld[50]),
.io_wt_actv_2_50_bits_nz(wt2_actv_nz[50]),
.io_wt_actv_2_50_bits_data(wt2_actv_data[407:400]),

.io_wt_actv_2_51_valid(wt2_actv_pvld[51]),
.io_wt_actv_2_51_bits_nz(wt2_actv_nz[51]),
.io_wt_actv_2_51_bits_data(wt2_actv_data[415:408]),

.io_wt_actv_2_52_valid(wt2_actv_pvld[52]),
.io_wt_actv_2_52_bits_nz(wt2_actv_nz[52]),
.io_wt_actv_2_52_bits_data(wt2_actv_data[423:416]),

.io_wt_actv_2_53_valid(wt2_actv_pvld[53]),
.io_wt_actv_2_53_bits_nz(wt2_actv_nz[53]),
.io_wt_actv_2_53_bits_data(wt2_actv_data[431:424]),

.io_wt_actv_2_54_valid(wt2_actv_pvld[54]),
.io_wt_actv_2_54_bits_nz(wt2_actv_nz[54]),
.io_wt_actv_2_54_bits_data(wt2_actv_data[439:432]),

.io_wt_actv_2_55_valid(wt2_actv_pvld[55]),
.io_wt_actv_2_55_bits_nz(wt2_actv_nz[55]),
.io_wt_actv_2_55_bits_data(wt2_actv_data[447:440]),

.io_wt_actv_2_56_valid(wt2_actv_pvld[56]),
.io_wt_actv_2_56_bits_nz(wt2_actv_nz[56]),
.io_wt_actv_2_56_bits_data(wt2_actv_data[455:448]),

.io_wt_actv_2_57_valid(wt2_actv_pvld[57]),
.io_wt_actv_2_57_bits_nz(wt2_actv_nz[57]),
.io_wt_actv_2_57_bits_data(wt2_actv_data[463:456]),

.io_wt_actv_2_58_valid(wt2_actv_pvld[58]),
.io_wt_actv_2_58_bits_nz(wt2_actv_nz[58]),
.io_wt_actv_2_58_bits_data(wt2_actv_data[471:464]),

.io_wt_actv_2_59_valid(wt2_actv_pvld[59]),
.io_wt_actv_2_59_bits_nz(wt2_actv_nz[59]),
.io_wt_actv_2_59_bits_data(wt2_actv_data[479:472]),

.io_wt_actv_2_60_valid(wt2_actv_pvld[60]),
.io_wt_actv_2_60_bits_nz(wt2_actv_nz[60]),
.io_wt_actv_2_60_bits_data(wt2_actv_data[487:480]),

.io_wt_actv_2_61_valid(wt2_actv_pvld[61]),
.io_wt_actv_2_61_bits_nz(wt2_actv_nz[61]),
.io_wt_actv_2_61_bits_data(wt2_actv_data[495:488]),

.io_wt_actv_2_62_valid(wt2_actv_pvld[62]),
.io_wt_actv_2_62_bits_nz(wt2_actv_nz[62]),
.io_wt_actv_2_62_bits_data(wt2_actv_data[503:496]),

.io_wt_actv_2_63_valid(wt2_actv_pvld[63]),
.io_wt_actv_2_63_bits_nz(wt2_actv_nz[63]),
.io_wt_actv_2_63_bits_data(wt2_actv_data[511:504]),

.io_wt_actv_3_0_valid(wt3_actv_pvld[0]),
.io_wt_actv_3_0_bits_nz(wt3_actv_nz[0]),
.io_wt_actv_3_0_bits_data(wt3_actv_data[7:0]),

.io_wt_actv_3_1_valid(wt3_actv_pvld[1]),
.io_wt_actv_3_1_bits_nz(wt3_actv_nz[1]),
.io_wt_actv_3_1_bits_data(wt3_actv_data[15:8]),

.io_wt_actv_3_2_valid(wt3_actv_pvld[2]),
.io_wt_actv_3_2_bits_nz(wt3_actv_nz[2]),
.io_wt_actv_3_2_bits_data(wt3_actv_data[23:16]),

.io_wt_actv_3_3_valid(wt3_actv_pvld[3]),
.io_wt_actv_3_3_bits_nz(wt3_actv_nz[3]),
.io_wt_actv_3_3_bits_data(wt3_actv_data[31:24]),

.io_wt_actv_3_4_valid(wt3_actv_pvld[4]),
.io_wt_actv_3_4_bits_nz(wt3_actv_nz[4]),
.io_wt_actv_3_4_bits_data(wt3_actv_data[39:32]),

.io_wt_actv_3_5_valid(wt3_actv_pvld[5]),
.io_wt_actv_3_5_bits_nz(wt3_actv_nz[5]),
.io_wt_actv_3_5_bits_data(wt3_actv_data[47:40]),

.io_wt_actv_3_6_valid(wt3_actv_pvld[6]),
.io_wt_actv_3_6_bits_nz(wt3_actv_nz[6]),
.io_wt_actv_3_6_bits_data(wt3_actv_data[55:48]),

.io_wt_actv_3_7_valid(wt3_actv_pvld[7]),
.io_wt_actv_3_7_bits_nz(wt3_actv_nz[7]),
.io_wt_actv_3_7_bits_data(wt3_actv_data[63:56]),

.io_wt_actv_3_8_valid(wt3_actv_pvld[8]),
.io_wt_actv_3_8_bits_nz(wt3_actv_nz[8]),
.io_wt_actv_3_8_bits_data(wt3_actv_data[71:64]),

.io_wt_actv_3_9_valid(wt3_actv_pvld[9]),
.io_wt_actv_3_9_bits_nz(wt3_actv_nz[9]),
.io_wt_actv_3_9_bits_data(wt3_actv_data[79:72]),

.io_wt_actv_3_10_valid(wt3_actv_pvld[10]),
.io_wt_actv_3_10_bits_nz(wt3_actv_nz[10]),
.io_wt_actv_3_10_bits_data(wt3_actv_data[87:80]),

.io_wt_actv_3_11_valid(wt3_actv_pvld[11]),
.io_wt_actv_3_11_bits_nz(wt3_actv_nz[11]),
.io_wt_actv_3_11_bits_data(wt3_actv_data[95:88]),

.io_wt_actv_3_12_valid(wt3_actv_pvld[12]),
.io_wt_actv_3_12_bits_nz(wt3_actv_nz[12]),
.io_wt_actv_3_12_bits_data(wt3_actv_data[103:96]),

.io_wt_actv_3_13_valid(wt3_actv_pvld[13]),
.io_wt_actv_3_13_bits_nz(wt3_actv_nz[13]),
.io_wt_actv_3_13_bits_data(wt3_actv_data[111:104]),

.io_wt_actv_3_14_valid(wt3_actv_pvld[14]),
.io_wt_actv_3_14_bits_nz(wt3_actv_nz[14]),
.io_wt_actv_3_14_bits_data(wt3_actv_data[119:112]),

.io_wt_actv_3_15_valid(wt3_actv_pvld[15]),
.io_wt_actv_3_15_bits_nz(wt3_actv_nz[15]),
.io_wt_actv_3_15_bits_data(wt3_actv_data[127:120]),

.io_wt_actv_3_16_valid(wt3_actv_pvld[16]),
.io_wt_actv_3_16_bits_nz(wt3_actv_nz[16]),
.io_wt_actv_3_16_bits_data(wt3_actv_data[135:128]),

.io_wt_actv_3_17_valid(wt3_actv_pvld[17]),
.io_wt_actv_3_17_bits_nz(wt3_actv_nz[17]),
.io_wt_actv_3_17_bits_data(wt3_actv_data[143:136]),

.io_wt_actv_3_18_valid(wt3_actv_pvld[18]),
.io_wt_actv_3_18_bits_nz(wt3_actv_nz[18]),
.io_wt_actv_3_18_bits_data(wt3_actv_data[151:144]),

.io_wt_actv_3_19_valid(wt3_actv_pvld[19]),
.io_wt_actv_3_19_bits_nz(wt3_actv_nz[19]),
.io_wt_actv_3_19_bits_data(wt3_actv_data[159:152]),

.io_wt_actv_3_20_valid(wt3_actv_pvld[20]),
.io_wt_actv_3_20_bits_nz(wt3_actv_nz[20]),
.io_wt_actv_3_20_bits_data(wt3_actv_data[167:160]),

.io_wt_actv_3_21_valid(wt3_actv_pvld[21]),
.io_wt_actv_3_21_bits_nz(wt3_actv_nz[21]),
.io_wt_actv_3_21_bits_data(wt3_actv_data[175:168]),

.io_wt_actv_3_22_valid(wt3_actv_pvld[22]),
.io_wt_actv_3_22_bits_nz(wt3_actv_nz[22]),
.io_wt_actv_3_22_bits_data(wt3_actv_data[183:176]),

.io_wt_actv_3_23_valid(wt3_actv_pvld[23]),
.io_wt_actv_3_23_bits_nz(wt3_actv_nz[23]),
.io_wt_actv_3_23_bits_data(wt3_actv_data[191:184]),

.io_wt_actv_3_24_valid(wt3_actv_pvld[24]),
.io_wt_actv_3_24_bits_nz(wt3_actv_nz[24]),
.io_wt_actv_3_24_bits_data(wt3_actv_data[199:192]),

.io_wt_actv_3_25_valid(wt3_actv_pvld[25]),
.io_wt_actv_3_25_bits_nz(wt3_actv_nz[25]),
.io_wt_actv_3_25_bits_data(wt3_actv_data[207:200]),

.io_wt_actv_3_26_valid(wt3_actv_pvld[26]),
.io_wt_actv_3_26_bits_nz(wt3_actv_nz[26]),
.io_wt_actv_3_26_bits_data(wt3_actv_data[215:208]),

.io_wt_actv_3_27_valid(wt3_actv_pvld[27]),
.io_wt_actv_3_27_bits_nz(wt3_actv_nz[27]),
.io_wt_actv_3_27_bits_data(wt3_actv_data[223:216]),

.io_wt_actv_3_28_valid(wt3_actv_pvld[28]),
.io_wt_actv_3_28_bits_nz(wt3_actv_nz[28]),
.io_wt_actv_3_28_bits_data(wt3_actv_data[231:224]),

.io_wt_actv_3_29_valid(wt3_actv_pvld[29]),
.io_wt_actv_3_29_bits_nz(wt3_actv_nz[29]),
.io_wt_actv_3_29_bits_data(wt3_actv_data[239:232]),

.io_wt_actv_3_30_valid(wt3_actv_pvld[30]),
.io_wt_actv_3_30_bits_nz(wt3_actv_nz[30]),
.io_wt_actv_3_30_bits_data(wt3_actv_data[247:240]),

.io_wt_actv_3_31_valid(wt3_actv_pvld[31]),
.io_wt_actv_3_31_bits_nz(wt3_actv_nz[31]),
.io_wt_actv_3_31_bits_data(wt3_actv_data[255:248]),

.io_wt_actv_3_32_valid(wt3_actv_pvld[32]),
.io_wt_actv_3_32_bits_nz(wt3_actv_nz[32]),
.io_wt_actv_3_32_bits_data(wt3_actv_data[263:256]),

.io_wt_actv_3_33_valid(wt3_actv_pvld[33]),
.io_wt_actv_3_33_bits_nz(wt3_actv_nz[33]),
.io_wt_actv_3_33_bits_data(wt3_actv_data[271:264]),

.io_wt_actv_3_34_valid(wt3_actv_pvld[34]),
.io_wt_actv_3_34_bits_nz(wt3_actv_nz[34]),
.io_wt_actv_3_34_bits_data(wt3_actv_data[279:272]),

.io_wt_actv_3_35_valid(wt3_actv_pvld[35]),
.io_wt_actv_3_35_bits_nz(wt3_actv_nz[35]),
.io_wt_actv_3_35_bits_data(wt3_actv_data[287:280]),

.io_wt_actv_3_36_valid(wt3_actv_pvld[36]),
.io_wt_actv_3_36_bits_nz(wt3_actv_nz[36]),
.io_wt_actv_3_36_bits_data(wt3_actv_data[295:288]),

.io_wt_actv_3_37_valid(wt3_actv_pvld[37]),
.io_wt_actv_3_37_bits_nz(wt3_actv_nz[37]),
.io_wt_actv_3_37_bits_data(wt3_actv_data[303:296]),

.io_wt_actv_3_38_valid(wt3_actv_pvld[38]),
.io_wt_actv_3_38_bits_nz(wt3_actv_nz[38]),
.io_wt_actv_3_38_bits_data(wt3_actv_data[311:304]),

.io_wt_actv_3_39_valid(wt3_actv_pvld[39]),
.io_wt_actv_3_39_bits_nz(wt3_actv_nz[39]),
.io_wt_actv_3_39_bits_data(wt3_actv_data[319:312]),

.io_wt_actv_3_40_valid(wt3_actv_pvld[40]),
.io_wt_actv_3_40_bits_nz(wt3_actv_nz[40]),
.io_wt_actv_3_40_bits_data(wt3_actv_data[327:320]),

.io_wt_actv_3_41_valid(wt3_actv_pvld[41]),
.io_wt_actv_3_41_bits_nz(wt3_actv_nz[41]),
.io_wt_actv_3_41_bits_data(wt3_actv_data[335:328]),

.io_wt_actv_3_42_valid(wt3_actv_pvld[42]),
.io_wt_actv_3_42_bits_nz(wt3_actv_nz[42]),
.io_wt_actv_3_42_bits_data(wt3_actv_data[343:336]),

.io_wt_actv_3_43_valid(wt3_actv_pvld[43]),
.io_wt_actv_3_43_bits_nz(wt3_actv_nz[43]),
.io_wt_actv_3_43_bits_data(wt3_actv_data[351:344]),

.io_wt_actv_3_44_valid(wt3_actv_pvld[44]),
.io_wt_actv_3_44_bits_nz(wt3_actv_nz[44]),
.io_wt_actv_3_44_bits_data(wt3_actv_data[359:352]),

.io_wt_actv_3_45_valid(wt3_actv_pvld[45]),
.io_wt_actv_3_45_bits_nz(wt3_actv_nz[45]),
.io_wt_actv_3_45_bits_data(wt3_actv_data[367:360]),

.io_wt_actv_3_46_valid(wt3_actv_pvld[46]),
.io_wt_actv_3_46_bits_nz(wt3_actv_nz[46]),
.io_wt_actv_3_46_bits_data(wt3_actv_data[375:368]),

.io_wt_actv_3_47_valid(wt3_actv_pvld[47]),
.io_wt_actv_3_47_bits_nz(wt3_actv_nz[47]),
.io_wt_actv_3_47_bits_data(wt3_actv_data[383:376]),

.io_wt_actv_3_48_valid(wt3_actv_pvld[48]),
.io_wt_actv_3_48_bits_nz(wt3_actv_nz[48]),
.io_wt_actv_3_48_bits_data(wt3_actv_data[391:384]),

.io_wt_actv_3_49_valid(wt3_actv_pvld[49]),
.io_wt_actv_3_49_bits_nz(wt3_actv_nz[49]),
.io_wt_actv_3_49_bits_data(wt3_actv_data[399:392]),

.io_wt_actv_3_50_valid(wt3_actv_pvld[50]),
.io_wt_actv_3_50_bits_nz(wt3_actv_nz[50]),
.io_wt_actv_3_50_bits_data(wt3_actv_data[407:400]),

.io_wt_actv_3_51_valid(wt3_actv_pvld[51]),
.io_wt_actv_3_51_bits_nz(wt3_actv_nz[51]),
.io_wt_actv_3_51_bits_data(wt3_actv_data[415:408]),

.io_wt_actv_3_52_valid(wt3_actv_pvld[52]),
.io_wt_actv_3_52_bits_nz(wt3_actv_nz[52]),
.io_wt_actv_3_52_bits_data(wt3_actv_data[423:416]),

.io_wt_actv_3_53_valid(wt3_actv_pvld[53]),
.io_wt_actv_3_53_bits_nz(wt3_actv_nz[53]),
.io_wt_actv_3_53_bits_data(wt3_actv_data[431:424]),

.io_wt_actv_3_54_valid(wt3_actv_pvld[54]),
.io_wt_actv_3_54_bits_nz(wt3_actv_nz[54]),
.io_wt_actv_3_54_bits_data(wt3_actv_data[439:432]),

.io_wt_actv_3_55_valid(wt3_actv_pvld[55]),
.io_wt_actv_3_55_bits_nz(wt3_actv_nz[55]),
.io_wt_actv_3_55_bits_data(wt3_actv_data[447:440]),

.io_wt_actv_3_56_valid(wt3_actv_pvld[56]),
.io_wt_actv_3_56_bits_nz(wt3_actv_nz[56]),
.io_wt_actv_3_56_bits_data(wt3_actv_data[455:448]),

.io_wt_actv_3_57_valid(wt3_actv_pvld[57]),
.io_wt_actv_3_57_bits_nz(wt3_actv_nz[57]),
.io_wt_actv_3_57_bits_data(wt3_actv_data[463:456]),

.io_wt_actv_3_58_valid(wt3_actv_pvld[58]),
.io_wt_actv_3_58_bits_nz(wt3_actv_nz[58]),
.io_wt_actv_3_58_bits_data(wt3_actv_data[471:464]),

.io_wt_actv_3_59_valid(wt3_actv_pvld[59]),
.io_wt_actv_3_59_bits_nz(wt3_actv_nz[59]),
.io_wt_actv_3_59_bits_data(wt3_actv_data[479:472]),

.io_wt_actv_3_60_valid(wt3_actv_pvld[60]),
.io_wt_actv_3_60_bits_nz(wt3_actv_nz[60]),
.io_wt_actv_3_60_bits_data(wt3_actv_data[487:480]),

.io_wt_actv_3_61_valid(wt3_actv_pvld[61]),
.io_wt_actv_3_61_bits_nz(wt3_actv_nz[61]),
.io_wt_actv_3_61_bits_data(wt3_actv_data[495:488]),

.io_wt_actv_3_62_valid(wt3_actv_pvld[62]),
.io_wt_actv_3_62_bits_nz(wt3_actv_nz[62]),
.io_wt_actv_3_62_bits_data(wt3_actv_data[503:496]),

.io_wt_actv_3_63_valid(wt3_actv_pvld[63]),
.io_wt_actv_3_63_bits_nz(wt3_actv_nz[63]),
.io_wt_actv_3_63_bits_data(wt3_actv_data[511:504]),

.io_wt_actv_4_0_valid(wt4_actv_pvld[0]),
.io_wt_actv_4_0_bits_nz(wt4_actv_nz[0]),
.io_wt_actv_4_0_bits_data(wt4_actv_data[7:0]),

.io_wt_actv_4_1_valid(wt4_actv_pvld[1]),
.io_wt_actv_4_1_bits_nz(wt4_actv_nz[1]),
.io_wt_actv_4_1_bits_data(wt4_actv_data[15:8]),

.io_wt_actv_4_2_valid(wt4_actv_pvld[2]),
.io_wt_actv_4_2_bits_nz(wt4_actv_nz[2]),
.io_wt_actv_4_2_bits_data(wt4_actv_data[23:16]),

.io_wt_actv_4_3_valid(wt4_actv_pvld[3]),
.io_wt_actv_4_3_bits_nz(wt4_actv_nz[3]),
.io_wt_actv_4_3_bits_data(wt4_actv_data[31:24]),

.io_wt_actv_4_4_valid(wt4_actv_pvld[4]),
.io_wt_actv_4_4_bits_nz(wt4_actv_nz[4]),
.io_wt_actv_4_4_bits_data(wt4_actv_data[39:32]),

.io_wt_actv_4_5_valid(wt4_actv_pvld[5]),
.io_wt_actv_4_5_bits_nz(wt4_actv_nz[5]),
.io_wt_actv_4_5_bits_data(wt4_actv_data[47:40]),

.io_wt_actv_4_6_valid(wt4_actv_pvld[6]),
.io_wt_actv_4_6_bits_nz(wt4_actv_nz[6]),
.io_wt_actv_4_6_bits_data(wt4_actv_data[55:48]),

.io_wt_actv_4_7_valid(wt4_actv_pvld[7]),
.io_wt_actv_4_7_bits_nz(wt4_actv_nz[7]),
.io_wt_actv_4_7_bits_data(wt4_actv_data[63:56]),

.io_wt_actv_4_8_valid(wt4_actv_pvld[8]),
.io_wt_actv_4_8_bits_nz(wt4_actv_nz[8]),
.io_wt_actv_4_8_bits_data(wt4_actv_data[71:64]),

.io_wt_actv_4_9_valid(wt4_actv_pvld[9]),
.io_wt_actv_4_9_bits_nz(wt4_actv_nz[9]),
.io_wt_actv_4_9_bits_data(wt4_actv_data[79:72]),

.io_wt_actv_4_10_valid(wt4_actv_pvld[10]),
.io_wt_actv_4_10_bits_nz(wt4_actv_nz[10]),
.io_wt_actv_4_10_bits_data(wt4_actv_data[87:80]),

.io_wt_actv_4_11_valid(wt4_actv_pvld[11]),
.io_wt_actv_4_11_bits_nz(wt4_actv_nz[11]),
.io_wt_actv_4_11_bits_data(wt4_actv_data[95:88]),

.io_wt_actv_4_12_valid(wt4_actv_pvld[12]),
.io_wt_actv_4_12_bits_nz(wt4_actv_nz[12]),
.io_wt_actv_4_12_bits_data(wt4_actv_data[103:96]),

.io_wt_actv_4_13_valid(wt4_actv_pvld[13]),
.io_wt_actv_4_13_bits_nz(wt4_actv_nz[13]),
.io_wt_actv_4_13_bits_data(wt4_actv_data[111:104]),

.io_wt_actv_4_14_valid(wt4_actv_pvld[14]),
.io_wt_actv_4_14_bits_nz(wt4_actv_nz[14]),
.io_wt_actv_4_14_bits_data(wt4_actv_data[119:112]),

.io_wt_actv_4_15_valid(wt4_actv_pvld[15]),
.io_wt_actv_4_15_bits_nz(wt4_actv_nz[15]),
.io_wt_actv_4_15_bits_data(wt4_actv_data[127:120]),

.io_wt_actv_4_16_valid(wt4_actv_pvld[16]),
.io_wt_actv_4_16_bits_nz(wt4_actv_nz[16]),
.io_wt_actv_4_16_bits_data(wt4_actv_data[135:128]),

.io_wt_actv_4_17_valid(wt4_actv_pvld[17]),
.io_wt_actv_4_17_bits_nz(wt4_actv_nz[17]),
.io_wt_actv_4_17_bits_data(wt4_actv_data[143:136]),

.io_wt_actv_4_18_valid(wt4_actv_pvld[18]),
.io_wt_actv_4_18_bits_nz(wt4_actv_nz[18]),
.io_wt_actv_4_18_bits_data(wt4_actv_data[151:144]),

.io_wt_actv_4_19_valid(wt4_actv_pvld[19]),
.io_wt_actv_4_19_bits_nz(wt4_actv_nz[19]),
.io_wt_actv_4_19_bits_data(wt4_actv_data[159:152]),

.io_wt_actv_4_20_valid(wt4_actv_pvld[20]),
.io_wt_actv_4_20_bits_nz(wt4_actv_nz[20]),
.io_wt_actv_4_20_bits_data(wt4_actv_data[167:160]),

.io_wt_actv_4_21_valid(wt4_actv_pvld[21]),
.io_wt_actv_4_21_bits_nz(wt4_actv_nz[21]),
.io_wt_actv_4_21_bits_data(wt4_actv_data[175:168]),

.io_wt_actv_4_22_valid(wt4_actv_pvld[22]),
.io_wt_actv_4_22_bits_nz(wt4_actv_nz[22]),
.io_wt_actv_4_22_bits_data(wt4_actv_data[183:176]),

.io_wt_actv_4_23_valid(wt4_actv_pvld[23]),
.io_wt_actv_4_23_bits_nz(wt4_actv_nz[23]),
.io_wt_actv_4_23_bits_data(wt4_actv_data[191:184]),

.io_wt_actv_4_24_valid(wt4_actv_pvld[24]),
.io_wt_actv_4_24_bits_nz(wt4_actv_nz[24]),
.io_wt_actv_4_24_bits_data(wt4_actv_data[199:192]),

.io_wt_actv_4_25_valid(wt4_actv_pvld[25]),
.io_wt_actv_4_25_bits_nz(wt4_actv_nz[25]),
.io_wt_actv_4_25_bits_data(wt4_actv_data[207:200]),

.io_wt_actv_4_26_valid(wt4_actv_pvld[26]),
.io_wt_actv_4_26_bits_nz(wt4_actv_nz[26]),
.io_wt_actv_4_26_bits_data(wt4_actv_data[215:208]),

.io_wt_actv_4_27_valid(wt4_actv_pvld[27]),
.io_wt_actv_4_27_bits_nz(wt4_actv_nz[27]),
.io_wt_actv_4_27_bits_data(wt4_actv_data[223:216]),

.io_wt_actv_4_28_valid(wt4_actv_pvld[28]),
.io_wt_actv_4_28_bits_nz(wt4_actv_nz[28]),
.io_wt_actv_4_28_bits_data(wt4_actv_data[231:224]),

.io_wt_actv_4_29_valid(wt4_actv_pvld[29]),
.io_wt_actv_4_29_bits_nz(wt4_actv_nz[29]),
.io_wt_actv_4_29_bits_data(wt4_actv_data[239:232]),

.io_wt_actv_4_30_valid(wt4_actv_pvld[30]),
.io_wt_actv_4_30_bits_nz(wt4_actv_nz[30]),
.io_wt_actv_4_30_bits_data(wt4_actv_data[247:240]),

.io_wt_actv_4_31_valid(wt4_actv_pvld[31]),
.io_wt_actv_4_31_bits_nz(wt4_actv_nz[31]),
.io_wt_actv_4_31_bits_data(wt4_actv_data[255:248]),

.io_wt_actv_4_32_valid(wt4_actv_pvld[32]),
.io_wt_actv_4_32_bits_nz(wt4_actv_nz[32]),
.io_wt_actv_4_32_bits_data(wt4_actv_data[263:256]),

.io_wt_actv_4_33_valid(wt4_actv_pvld[33]),
.io_wt_actv_4_33_bits_nz(wt4_actv_nz[33]),
.io_wt_actv_4_33_bits_data(wt4_actv_data[271:264]),

.io_wt_actv_4_34_valid(wt4_actv_pvld[34]),
.io_wt_actv_4_34_bits_nz(wt4_actv_nz[34]),
.io_wt_actv_4_34_bits_data(wt4_actv_data[279:272]),

.io_wt_actv_4_35_valid(wt4_actv_pvld[35]),
.io_wt_actv_4_35_bits_nz(wt4_actv_nz[35]),
.io_wt_actv_4_35_bits_data(wt4_actv_data[287:280]),

.io_wt_actv_4_36_valid(wt4_actv_pvld[36]),
.io_wt_actv_4_36_bits_nz(wt4_actv_nz[36]),
.io_wt_actv_4_36_bits_data(wt4_actv_data[295:288]),

.io_wt_actv_4_37_valid(wt4_actv_pvld[37]),
.io_wt_actv_4_37_bits_nz(wt4_actv_nz[37]),
.io_wt_actv_4_37_bits_data(wt4_actv_data[303:296]),

.io_wt_actv_4_38_valid(wt4_actv_pvld[38]),
.io_wt_actv_4_38_bits_nz(wt4_actv_nz[38]),
.io_wt_actv_4_38_bits_data(wt4_actv_data[311:304]),

.io_wt_actv_4_39_valid(wt4_actv_pvld[39]),
.io_wt_actv_4_39_bits_nz(wt4_actv_nz[39]),
.io_wt_actv_4_39_bits_data(wt4_actv_data[319:312]),

.io_wt_actv_4_40_valid(wt4_actv_pvld[40]),
.io_wt_actv_4_40_bits_nz(wt4_actv_nz[40]),
.io_wt_actv_4_40_bits_data(wt4_actv_data[327:320]),

.io_wt_actv_4_41_valid(wt4_actv_pvld[41]),
.io_wt_actv_4_41_bits_nz(wt4_actv_nz[41]),
.io_wt_actv_4_41_bits_data(wt4_actv_data[335:328]),

.io_wt_actv_4_42_valid(wt4_actv_pvld[42]),
.io_wt_actv_4_42_bits_nz(wt4_actv_nz[42]),
.io_wt_actv_4_42_bits_data(wt4_actv_data[343:336]),

.io_wt_actv_4_43_valid(wt4_actv_pvld[43]),
.io_wt_actv_4_43_bits_nz(wt4_actv_nz[43]),
.io_wt_actv_4_43_bits_data(wt4_actv_data[351:344]),

.io_wt_actv_4_44_valid(wt4_actv_pvld[44]),
.io_wt_actv_4_44_bits_nz(wt4_actv_nz[44]),
.io_wt_actv_4_44_bits_data(wt4_actv_data[359:352]),

.io_wt_actv_4_45_valid(wt4_actv_pvld[45]),
.io_wt_actv_4_45_bits_nz(wt4_actv_nz[45]),
.io_wt_actv_4_45_bits_data(wt4_actv_data[367:360]),

.io_wt_actv_4_46_valid(wt4_actv_pvld[46]),
.io_wt_actv_4_46_bits_nz(wt4_actv_nz[46]),
.io_wt_actv_4_46_bits_data(wt4_actv_data[375:368]),

.io_wt_actv_4_47_valid(wt4_actv_pvld[47]),
.io_wt_actv_4_47_bits_nz(wt4_actv_nz[47]),
.io_wt_actv_4_47_bits_data(wt4_actv_data[383:376]),

.io_wt_actv_4_48_valid(wt4_actv_pvld[48]),
.io_wt_actv_4_48_bits_nz(wt4_actv_nz[48]),
.io_wt_actv_4_48_bits_data(wt4_actv_data[391:384]),

.io_wt_actv_4_49_valid(wt4_actv_pvld[49]),
.io_wt_actv_4_49_bits_nz(wt4_actv_nz[49]),
.io_wt_actv_4_49_bits_data(wt4_actv_data[399:392]),

.io_wt_actv_4_50_valid(wt4_actv_pvld[50]),
.io_wt_actv_4_50_bits_nz(wt4_actv_nz[50]),
.io_wt_actv_4_50_bits_data(wt4_actv_data[407:400]),

.io_wt_actv_4_51_valid(wt4_actv_pvld[51]),
.io_wt_actv_4_51_bits_nz(wt4_actv_nz[51]),
.io_wt_actv_4_51_bits_data(wt4_actv_data[415:408]),

.io_wt_actv_4_52_valid(wt4_actv_pvld[52]),
.io_wt_actv_4_52_bits_nz(wt4_actv_nz[52]),
.io_wt_actv_4_52_bits_data(wt4_actv_data[423:416]),

.io_wt_actv_4_53_valid(wt4_actv_pvld[53]),
.io_wt_actv_4_53_bits_nz(wt4_actv_nz[53]),
.io_wt_actv_4_53_bits_data(wt4_actv_data[431:424]),

.io_wt_actv_4_54_valid(wt4_actv_pvld[54]),
.io_wt_actv_4_54_bits_nz(wt4_actv_nz[54]),
.io_wt_actv_4_54_bits_data(wt4_actv_data[439:432]),

.io_wt_actv_4_55_valid(wt4_actv_pvld[55]),
.io_wt_actv_4_55_bits_nz(wt4_actv_nz[55]),
.io_wt_actv_4_55_bits_data(wt4_actv_data[447:440]),

.io_wt_actv_4_56_valid(wt4_actv_pvld[56]),
.io_wt_actv_4_56_bits_nz(wt4_actv_nz[56]),
.io_wt_actv_4_56_bits_data(wt4_actv_data[455:448]),

.io_wt_actv_4_57_valid(wt4_actv_pvld[57]),
.io_wt_actv_4_57_bits_nz(wt4_actv_nz[57]),
.io_wt_actv_4_57_bits_data(wt4_actv_data[463:456]),

.io_wt_actv_4_58_valid(wt4_actv_pvld[58]),
.io_wt_actv_4_58_bits_nz(wt4_actv_nz[58]),
.io_wt_actv_4_58_bits_data(wt4_actv_data[471:464]),

.io_wt_actv_4_59_valid(wt4_actv_pvld[59]),
.io_wt_actv_4_59_bits_nz(wt4_actv_nz[59]),
.io_wt_actv_4_59_bits_data(wt4_actv_data[479:472]),

.io_wt_actv_4_60_valid(wt4_actv_pvld[60]),
.io_wt_actv_4_60_bits_nz(wt4_actv_nz[60]),
.io_wt_actv_4_60_bits_data(wt4_actv_data[487:480]),

.io_wt_actv_4_61_valid(wt4_actv_pvld[61]),
.io_wt_actv_4_61_bits_nz(wt4_actv_nz[61]),
.io_wt_actv_4_61_bits_data(wt4_actv_data[495:488]),

.io_wt_actv_4_62_valid(wt4_actv_pvld[62]),
.io_wt_actv_4_62_bits_nz(wt4_actv_nz[62]),
.io_wt_actv_4_62_bits_data(wt4_actv_data[503:496]),

.io_wt_actv_4_63_valid(wt4_actv_pvld[63]),
.io_wt_actv_4_63_bits_nz(wt4_actv_nz[63]),
.io_wt_actv_4_63_bits_data(wt4_actv_data[511:504]),

.io_wt_actv_5_0_valid(wt5_actv_pvld[0]),
.io_wt_actv_5_0_bits_nz(wt5_actv_nz[0]),
.io_wt_actv_5_0_bits_data(wt5_actv_data[7:0]),

.io_wt_actv_5_1_valid(wt5_actv_pvld[1]),
.io_wt_actv_5_1_bits_nz(wt5_actv_nz[1]),
.io_wt_actv_5_1_bits_data(wt5_actv_data[15:8]),

.io_wt_actv_5_2_valid(wt5_actv_pvld[2]),
.io_wt_actv_5_2_bits_nz(wt5_actv_nz[2]),
.io_wt_actv_5_2_bits_data(wt5_actv_data[23:16]),

.io_wt_actv_5_3_valid(wt5_actv_pvld[3]),
.io_wt_actv_5_3_bits_nz(wt5_actv_nz[3]),
.io_wt_actv_5_3_bits_data(wt5_actv_data[31:24]),

.io_wt_actv_5_4_valid(wt5_actv_pvld[4]),
.io_wt_actv_5_4_bits_nz(wt5_actv_nz[4]),
.io_wt_actv_5_4_bits_data(wt5_actv_data[39:32]),

.io_wt_actv_5_5_valid(wt5_actv_pvld[5]),
.io_wt_actv_5_5_bits_nz(wt5_actv_nz[5]),
.io_wt_actv_5_5_bits_data(wt5_actv_data[47:40]),

.io_wt_actv_5_6_valid(wt5_actv_pvld[6]),
.io_wt_actv_5_6_bits_nz(wt5_actv_nz[6]),
.io_wt_actv_5_6_bits_data(wt5_actv_data[55:48]),

.io_wt_actv_5_7_valid(wt5_actv_pvld[7]),
.io_wt_actv_5_7_bits_nz(wt5_actv_nz[7]),
.io_wt_actv_5_7_bits_data(wt5_actv_data[63:56]),

.io_wt_actv_5_8_valid(wt5_actv_pvld[8]),
.io_wt_actv_5_8_bits_nz(wt5_actv_nz[8]),
.io_wt_actv_5_8_bits_data(wt5_actv_data[71:64]),

.io_wt_actv_5_9_valid(wt5_actv_pvld[9]),
.io_wt_actv_5_9_bits_nz(wt5_actv_nz[9]),
.io_wt_actv_5_9_bits_data(wt5_actv_data[79:72]),

.io_wt_actv_5_10_valid(wt5_actv_pvld[10]),
.io_wt_actv_5_10_bits_nz(wt5_actv_nz[10]),
.io_wt_actv_5_10_bits_data(wt5_actv_data[87:80]),

.io_wt_actv_5_11_valid(wt5_actv_pvld[11]),
.io_wt_actv_5_11_bits_nz(wt5_actv_nz[11]),
.io_wt_actv_5_11_bits_data(wt5_actv_data[95:88]),

.io_wt_actv_5_12_valid(wt5_actv_pvld[12]),
.io_wt_actv_5_12_bits_nz(wt5_actv_nz[12]),
.io_wt_actv_5_12_bits_data(wt5_actv_data[103:96]),

.io_wt_actv_5_13_valid(wt5_actv_pvld[13]),
.io_wt_actv_5_13_bits_nz(wt5_actv_nz[13]),
.io_wt_actv_5_13_bits_data(wt5_actv_data[111:104]),

.io_wt_actv_5_14_valid(wt5_actv_pvld[14]),
.io_wt_actv_5_14_bits_nz(wt5_actv_nz[14]),
.io_wt_actv_5_14_bits_data(wt5_actv_data[119:112]),

.io_wt_actv_5_15_valid(wt5_actv_pvld[15]),
.io_wt_actv_5_15_bits_nz(wt5_actv_nz[15]),
.io_wt_actv_5_15_bits_data(wt5_actv_data[127:120]),

.io_wt_actv_5_16_valid(wt5_actv_pvld[16]),
.io_wt_actv_5_16_bits_nz(wt5_actv_nz[16]),
.io_wt_actv_5_16_bits_data(wt5_actv_data[135:128]),

.io_wt_actv_5_17_valid(wt5_actv_pvld[17]),
.io_wt_actv_5_17_bits_nz(wt5_actv_nz[17]),
.io_wt_actv_5_17_bits_data(wt5_actv_data[143:136]),

.io_wt_actv_5_18_valid(wt5_actv_pvld[18]),
.io_wt_actv_5_18_bits_nz(wt5_actv_nz[18]),
.io_wt_actv_5_18_bits_data(wt5_actv_data[151:144]),

.io_wt_actv_5_19_valid(wt5_actv_pvld[19]),
.io_wt_actv_5_19_bits_nz(wt5_actv_nz[19]),
.io_wt_actv_5_19_bits_data(wt5_actv_data[159:152]),

.io_wt_actv_5_20_valid(wt5_actv_pvld[20]),
.io_wt_actv_5_20_bits_nz(wt5_actv_nz[20]),
.io_wt_actv_5_20_bits_data(wt5_actv_data[167:160]),

.io_wt_actv_5_21_valid(wt5_actv_pvld[21]),
.io_wt_actv_5_21_bits_nz(wt5_actv_nz[21]),
.io_wt_actv_5_21_bits_data(wt5_actv_data[175:168]),

.io_wt_actv_5_22_valid(wt5_actv_pvld[22]),
.io_wt_actv_5_22_bits_nz(wt5_actv_nz[22]),
.io_wt_actv_5_22_bits_data(wt5_actv_data[183:176]),

.io_wt_actv_5_23_valid(wt5_actv_pvld[23]),
.io_wt_actv_5_23_bits_nz(wt5_actv_nz[23]),
.io_wt_actv_5_23_bits_data(wt5_actv_data[191:184]),

.io_wt_actv_5_24_valid(wt5_actv_pvld[24]),
.io_wt_actv_5_24_bits_nz(wt5_actv_nz[24]),
.io_wt_actv_5_24_bits_data(wt5_actv_data[199:192]),

.io_wt_actv_5_25_valid(wt5_actv_pvld[25]),
.io_wt_actv_5_25_bits_nz(wt5_actv_nz[25]),
.io_wt_actv_5_25_bits_data(wt5_actv_data[207:200]),

.io_wt_actv_5_26_valid(wt5_actv_pvld[26]),
.io_wt_actv_5_26_bits_nz(wt5_actv_nz[26]),
.io_wt_actv_5_26_bits_data(wt5_actv_data[215:208]),

.io_wt_actv_5_27_valid(wt5_actv_pvld[27]),
.io_wt_actv_5_27_bits_nz(wt5_actv_nz[27]),
.io_wt_actv_5_27_bits_data(wt5_actv_data[223:216]),

.io_wt_actv_5_28_valid(wt5_actv_pvld[28]),
.io_wt_actv_5_28_bits_nz(wt5_actv_nz[28]),
.io_wt_actv_5_28_bits_data(wt5_actv_data[231:224]),

.io_wt_actv_5_29_valid(wt5_actv_pvld[29]),
.io_wt_actv_5_29_bits_nz(wt5_actv_nz[29]),
.io_wt_actv_5_29_bits_data(wt5_actv_data[239:232]),

.io_wt_actv_5_30_valid(wt5_actv_pvld[30]),
.io_wt_actv_5_30_bits_nz(wt5_actv_nz[30]),
.io_wt_actv_5_30_bits_data(wt5_actv_data[247:240]),

.io_wt_actv_5_31_valid(wt5_actv_pvld[31]),
.io_wt_actv_5_31_bits_nz(wt5_actv_nz[31]),
.io_wt_actv_5_31_bits_data(wt5_actv_data[255:248]),

.io_wt_actv_5_32_valid(wt5_actv_pvld[32]),
.io_wt_actv_5_32_bits_nz(wt5_actv_nz[32]),
.io_wt_actv_5_32_bits_data(wt5_actv_data[263:256]),

.io_wt_actv_5_33_valid(wt5_actv_pvld[33]),
.io_wt_actv_5_33_bits_nz(wt5_actv_nz[33]),
.io_wt_actv_5_33_bits_data(wt5_actv_data[271:264]),

.io_wt_actv_5_34_valid(wt5_actv_pvld[34]),
.io_wt_actv_5_34_bits_nz(wt5_actv_nz[34]),
.io_wt_actv_5_34_bits_data(wt5_actv_data[279:272]),

.io_wt_actv_5_35_valid(wt5_actv_pvld[35]),
.io_wt_actv_5_35_bits_nz(wt5_actv_nz[35]),
.io_wt_actv_5_35_bits_data(wt5_actv_data[287:280]),

.io_wt_actv_5_36_valid(wt5_actv_pvld[36]),
.io_wt_actv_5_36_bits_nz(wt5_actv_nz[36]),
.io_wt_actv_5_36_bits_data(wt5_actv_data[295:288]),

.io_wt_actv_5_37_valid(wt5_actv_pvld[37]),
.io_wt_actv_5_37_bits_nz(wt5_actv_nz[37]),
.io_wt_actv_5_37_bits_data(wt5_actv_data[303:296]),

.io_wt_actv_5_38_valid(wt5_actv_pvld[38]),
.io_wt_actv_5_38_bits_nz(wt5_actv_nz[38]),
.io_wt_actv_5_38_bits_data(wt5_actv_data[311:304]),

.io_wt_actv_5_39_valid(wt5_actv_pvld[39]),
.io_wt_actv_5_39_bits_nz(wt5_actv_nz[39]),
.io_wt_actv_5_39_bits_data(wt5_actv_data[319:312]),

.io_wt_actv_5_40_valid(wt5_actv_pvld[40]),
.io_wt_actv_5_40_bits_nz(wt5_actv_nz[40]),
.io_wt_actv_5_40_bits_data(wt5_actv_data[327:320]),

.io_wt_actv_5_41_valid(wt5_actv_pvld[41]),
.io_wt_actv_5_41_bits_nz(wt5_actv_nz[41]),
.io_wt_actv_5_41_bits_data(wt5_actv_data[335:328]),

.io_wt_actv_5_42_valid(wt5_actv_pvld[42]),
.io_wt_actv_5_42_bits_nz(wt5_actv_nz[42]),
.io_wt_actv_5_42_bits_data(wt5_actv_data[343:336]),

.io_wt_actv_5_43_valid(wt5_actv_pvld[43]),
.io_wt_actv_5_43_bits_nz(wt5_actv_nz[43]),
.io_wt_actv_5_43_bits_data(wt5_actv_data[351:344]),

.io_wt_actv_5_44_valid(wt5_actv_pvld[44]),
.io_wt_actv_5_44_bits_nz(wt5_actv_nz[44]),
.io_wt_actv_5_44_bits_data(wt5_actv_data[359:352]),

.io_wt_actv_5_45_valid(wt5_actv_pvld[45]),
.io_wt_actv_5_45_bits_nz(wt5_actv_nz[45]),
.io_wt_actv_5_45_bits_data(wt5_actv_data[367:360]),

.io_wt_actv_5_46_valid(wt5_actv_pvld[46]),
.io_wt_actv_5_46_bits_nz(wt5_actv_nz[46]),
.io_wt_actv_5_46_bits_data(wt5_actv_data[375:368]),

.io_wt_actv_5_47_valid(wt5_actv_pvld[47]),
.io_wt_actv_5_47_bits_nz(wt5_actv_nz[47]),
.io_wt_actv_5_47_bits_data(wt5_actv_data[383:376]),

.io_wt_actv_5_48_valid(wt5_actv_pvld[48]),
.io_wt_actv_5_48_bits_nz(wt5_actv_nz[48]),
.io_wt_actv_5_48_bits_data(wt5_actv_data[391:384]),

.io_wt_actv_5_49_valid(wt5_actv_pvld[49]),
.io_wt_actv_5_49_bits_nz(wt5_actv_nz[49]),
.io_wt_actv_5_49_bits_data(wt5_actv_data[399:392]),

.io_wt_actv_5_50_valid(wt5_actv_pvld[50]),
.io_wt_actv_5_50_bits_nz(wt5_actv_nz[50]),
.io_wt_actv_5_50_bits_data(wt5_actv_data[407:400]),

.io_wt_actv_5_51_valid(wt5_actv_pvld[51]),
.io_wt_actv_5_51_bits_nz(wt5_actv_nz[51]),
.io_wt_actv_5_51_bits_data(wt5_actv_data[415:408]),

.io_wt_actv_5_52_valid(wt5_actv_pvld[52]),
.io_wt_actv_5_52_bits_nz(wt5_actv_nz[52]),
.io_wt_actv_5_52_bits_data(wt5_actv_data[423:416]),

.io_wt_actv_5_53_valid(wt5_actv_pvld[53]),
.io_wt_actv_5_53_bits_nz(wt5_actv_nz[53]),
.io_wt_actv_5_53_bits_data(wt5_actv_data[431:424]),

.io_wt_actv_5_54_valid(wt5_actv_pvld[54]),
.io_wt_actv_5_54_bits_nz(wt5_actv_nz[54]),
.io_wt_actv_5_54_bits_data(wt5_actv_data[439:432]),

.io_wt_actv_5_55_valid(wt5_actv_pvld[55]),
.io_wt_actv_5_55_bits_nz(wt5_actv_nz[55]),
.io_wt_actv_5_55_bits_data(wt5_actv_data[447:440]),

.io_wt_actv_5_56_valid(wt5_actv_pvld[56]),
.io_wt_actv_5_56_bits_nz(wt5_actv_nz[56]),
.io_wt_actv_5_56_bits_data(wt5_actv_data[455:448]),

.io_wt_actv_5_57_valid(wt5_actv_pvld[57]),
.io_wt_actv_5_57_bits_nz(wt5_actv_nz[57]),
.io_wt_actv_5_57_bits_data(wt5_actv_data[463:456]),

.io_wt_actv_5_58_valid(wt5_actv_pvld[58]),
.io_wt_actv_5_58_bits_nz(wt5_actv_nz[58]),
.io_wt_actv_5_58_bits_data(wt5_actv_data[471:464]),

.io_wt_actv_5_59_valid(wt5_actv_pvld[59]),
.io_wt_actv_5_59_bits_nz(wt5_actv_nz[59]),
.io_wt_actv_5_59_bits_data(wt5_actv_data[479:472]),

.io_wt_actv_5_60_valid(wt5_actv_pvld[60]),
.io_wt_actv_5_60_bits_nz(wt5_actv_nz[60]),
.io_wt_actv_5_60_bits_data(wt5_actv_data[487:480]),

.io_wt_actv_5_61_valid(wt5_actv_pvld[61]),
.io_wt_actv_5_61_bits_nz(wt5_actv_nz[61]),
.io_wt_actv_5_61_bits_data(wt5_actv_data[495:488]),

.io_wt_actv_5_62_valid(wt5_actv_pvld[62]),
.io_wt_actv_5_62_bits_nz(wt5_actv_nz[62]),
.io_wt_actv_5_62_bits_data(wt5_actv_data[503:496]),

.io_wt_actv_5_63_valid(wt5_actv_pvld[63]),
.io_wt_actv_5_63_bits_nz(wt5_actv_nz[63]),
.io_wt_actv_5_63_bits_data(wt5_actv_data[511:504]),

.io_wt_actv_6_0_valid(wt6_actv_pvld[0]),
.io_wt_actv_6_0_bits_nz(wt6_actv_nz[0]),
.io_wt_actv_6_0_bits_data(wt6_actv_data[7:0]),

.io_wt_actv_6_1_valid(wt6_actv_pvld[1]),
.io_wt_actv_6_1_bits_nz(wt6_actv_nz[1]),
.io_wt_actv_6_1_bits_data(wt6_actv_data[15:8]),

.io_wt_actv_6_2_valid(wt6_actv_pvld[2]),
.io_wt_actv_6_2_bits_nz(wt6_actv_nz[2]),
.io_wt_actv_6_2_bits_data(wt6_actv_data[23:16]),

.io_wt_actv_6_3_valid(wt6_actv_pvld[3]),
.io_wt_actv_6_3_bits_nz(wt6_actv_nz[3]),
.io_wt_actv_6_3_bits_data(wt6_actv_data[31:24]),

.io_wt_actv_6_4_valid(wt6_actv_pvld[4]),
.io_wt_actv_6_4_bits_nz(wt6_actv_nz[4]),
.io_wt_actv_6_4_bits_data(wt6_actv_data[39:32]),

.io_wt_actv_6_5_valid(wt6_actv_pvld[5]),
.io_wt_actv_6_5_bits_nz(wt6_actv_nz[5]),
.io_wt_actv_6_5_bits_data(wt6_actv_data[47:40]),

.io_wt_actv_6_6_valid(wt6_actv_pvld[6]),
.io_wt_actv_6_6_bits_nz(wt6_actv_nz[6]),
.io_wt_actv_6_6_bits_data(wt6_actv_data[55:48]),

.io_wt_actv_6_7_valid(wt6_actv_pvld[7]),
.io_wt_actv_6_7_bits_nz(wt6_actv_nz[7]),
.io_wt_actv_6_7_bits_data(wt6_actv_data[63:56]),

.io_wt_actv_6_8_valid(wt6_actv_pvld[8]),
.io_wt_actv_6_8_bits_nz(wt6_actv_nz[8]),
.io_wt_actv_6_8_bits_data(wt6_actv_data[71:64]),

.io_wt_actv_6_9_valid(wt6_actv_pvld[9]),
.io_wt_actv_6_9_bits_nz(wt6_actv_nz[9]),
.io_wt_actv_6_9_bits_data(wt6_actv_data[79:72]),

.io_wt_actv_6_10_valid(wt6_actv_pvld[10]),
.io_wt_actv_6_10_bits_nz(wt6_actv_nz[10]),
.io_wt_actv_6_10_bits_data(wt6_actv_data[87:80]),

.io_wt_actv_6_11_valid(wt6_actv_pvld[11]),
.io_wt_actv_6_11_bits_nz(wt6_actv_nz[11]),
.io_wt_actv_6_11_bits_data(wt6_actv_data[95:88]),

.io_wt_actv_6_12_valid(wt6_actv_pvld[12]),
.io_wt_actv_6_12_bits_nz(wt6_actv_nz[12]),
.io_wt_actv_6_12_bits_data(wt6_actv_data[103:96]),

.io_wt_actv_6_13_valid(wt6_actv_pvld[13]),
.io_wt_actv_6_13_bits_nz(wt6_actv_nz[13]),
.io_wt_actv_6_13_bits_data(wt6_actv_data[111:104]),

.io_wt_actv_6_14_valid(wt6_actv_pvld[14]),
.io_wt_actv_6_14_bits_nz(wt6_actv_nz[14]),
.io_wt_actv_6_14_bits_data(wt6_actv_data[119:112]),

.io_wt_actv_6_15_valid(wt6_actv_pvld[15]),
.io_wt_actv_6_15_bits_nz(wt6_actv_nz[15]),
.io_wt_actv_6_15_bits_data(wt6_actv_data[127:120]),

.io_wt_actv_6_16_valid(wt6_actv_pvld[16]),
.io_wt_actv_6_16_bits_nz(wt6_actv_nz[16]),
.io_wt_actv_6_16_bits_data(wt6_actv_data[135:128]),

.io_wt_actv_6_17_valid(wt6_actv_pvld[17]),
.io_wt_actv_6_17_bits_nz(wt6_actv_nz[17]),
.io_wt_actv_6_17_bits_data(wt6_actv_data[143:136]),

.io_wt_actv_6_18_valid(wt6_actv_pvld[18]),
.io_wt_actv_6_18_bits_nz(wt6_actv_nz[18]),
.io_wt_actv_6_18_bits_data(wt6_actv_data[151:144]),

.io_wt_actv_6_19_valid(wt6_actv_pvld[19]),
.io_wt_actv_6_19_bits_nz(wt6_actv_nz[19]),
.io_wt_actv_6_19_bits_data(wt6_actv_data[159:152]),

.io_wt_actv_6_20_valid(wt6_actv_pvld[20]),
.io_wt_actv_6_20_bits_nz(wt6_actv_nz[20]),
.io_wt_actv_6_20_bits_data(wt6_actv_data[167:160]),

.io_wt_actv_6_21_valid(wt6_actv_pvld[21]),
.io_wt_actv_6_21_bits_nz(wt6_actv_nz[21]),
.io_wt_actv_6_21_bits_data(wt6_actv_data[175:168]),

.io_wt_actv_6_22_valid(wt6_actv_pvld[22]),
.io_wt_actv_6_22_bits_nz(wt6_actv_nz[22]),
.io_wt_actv_6_22_bits_data(wt6_actv_data[183:176]),

.io_wt_actv_6_23_valid(wt6_actv_pvld[23]),
.io_wt_actv_6_23_bits_nz(wt6_actv_nz[23]),
.io_wt_actv_6_23_bits_data(wt6_actv_data[191:184]),

.io_wt_actv_6_24_valid(wt6_actv_pvld[24]),
.io_wt_actv_6_24_bits_nz(wt6_actv_nz[24]),
.io_wt_actv_6_24_bits_data(wt6_actv_data[199:192]),

.io_wt_actv_6_25_valid(wt6_actv_pvld[25]),
.io_wt_actv_6_25_bits_nz(wt6_actv_nz[25]),
.io_wt_actv_6_25_bits_data(wt6_actv_data[207:200]),

.io_wt_actv_6_26_valid(wt6_actv_pvld[26]),
.io_wt_actv_6_26_bits_nz(wt6_actv_nz[26]),
.io_wt_actv_6_26_bits_data(wt6_actv_data[215:208]),

.io_wt_actv_6_27_valid(wt6_actv_pvld[27]),
.io_wt_actv_6_27_bits_nz(wt6_actv_nz[27]),
.io_wt_actv_6_27_bits_data(wt6_actv_data[223:216]),

.io_wt_actv_6_28_valid(wt6_actv_pvld[28]),
.io_wt_actv_6_28_bits_nz(wt6_actv_nz[28]),
.io_wt_actv_6_28_bits_data(wt6_actv_data[231:224]),

.io_wt_actv_6_29_valid(wt6_actv_pvld[29]),
.io_wt_actv_6_29_bits_nz(wt6_actv_nz[29]),
.io_wt_actv_6_29_bits_data(wt6_actv_data[239:232]),

.io_wt_actv_6_30_valid(wt6_actv_pvld[30]),
.io_wt_actv_6_30_bits_nz(wt6_actv_nz[30]),
.io_wt_actv_6_30_bits_data(wt6_actv_data[247:240]),

.io_wt_actv_6_31_valid(wt6_actv_pvld[31]),
.io_wt_actv_6_31_bits_nz(wt6_actv_nz[31]),
.io_wt_actv_6_31_bits_data(wt6_actv_data[255:248]),

.io_wt_actv_6_32_valid(wt6_actv_pvld[32]),
.io_wt_actv_6_32_bits_nz(wt6_actv_nz[32]),
.io_wt_actv_6_32_bits_data(wt6_actv_data[263:256]),

.io_wt_actv_6_33_valid(wt6_actv_pvld[33]),
.io_wt_actv_6_33_bits_nz(wt6_actv_nz[33]),
.io_wt_actv_6_33_bits_data(wt6_actv_data[271:264]),

.io_wt_actv_6_34_valid(wt6_actv_pvld[34]),
.io_wt_actv_6_34_bits_nz(wt6_actv_nz[34]),
.io_wt_actv_6_34_bits_data(wt6_actv_data[279:272]),

.io_wt_actv_6_35_valid(wt6_actv_pvld[35]),
.io_wt_actv_6_35_bits_nz(wt6_actv_nz[35]),
.io_wt_actv_6_35_bits_data(wt6_actv_data[287:280]),

.io_wt_actv_6_36_valid(wt6_actv_pvld[36]),
.io_wt_actv_6_36_bits_nz(wt6_actv_nz[36]),
.io_wt_actv_6_36_bits_data(wt6_actv_data[295:288]),

.io_wt_actv_6_37_valid(wt6_actv_pvld[37]),
.io_wt_actv_6_37_bits_nz(wt6_actv_nz[37]),
.io_wt_actv_6_37_bits_data(wt6_actv_data[303:296]),

.io_wt_actv_6_38_valid(wt6_actv_pvld[38]),
.io_wt_actv_6_38_bits_nz(wt6_actv_nz[38]),
.io_wt_actv_6_38_bits_data(wt6_actv_data[311:304]),

.io_wt_actv_6_39_valid(wt6_actv_pvld[39]),
.io_wt_actv_6_39_bits_nz(wt6_actv_nz[39]),
.io_wt_actv_6_39_bits_data(wt6_actv_data[319:312]),

.io_wt_actv_6_40_valid(wt6_actv_pvld[40]),
.io_wt_actv_6_40_bits_nz(wt6_actv_nz[40]),
.io_wt_actv_6_40_bits_data(wt6_actv_data[327:320]),

.io_wt_actv_6_41_valid(wt6_actv_pvld[41]),
.io_wt_actv_6_41_bits_nz(wt6_actv_nz[41]),
.io_wt_actv_6_41_bits_data(wt6_actv_data[335:328]),

.io_wt_actv_6_42_valid(wt6_actv_pvld[42]),
.io_wt_actv_6_42_bits_nz(wt6_actv_nz[42]),
.io_wt_actv_6_42_bits_data(wt6_actv_data[343:336]),

.io_wt_actv_6_43_valid(wt6_actv_pvld[43]),
.io_wt_actv_6_43_bits_nz(wt6_actv_nz[43]),
.io_wt_actv_6_43_bits_data(wt6_actv_data[351:344]),

.io_wt_actv_6_44_valid(wt6_actv_pvld[44]),
.io_wt_actv_6_44_bits_nz(wt6_actv_nz[44]),
.io_wt_actv_6_44_bits_data(wt6_actv_data[359:352]),

.io_wt_actv_6_45_valid(wt6_actv_pvld[45]),
.io_wt_actv_6_45_bits_nz(wt6_actv_nz[45]),
.io_wt_actv_6_45_bits_data(wt6_actv_data[367:360]),

.io_wt_actv_6_46_valid(wt6_actv_pvld[46]),
.io_wt_actv_6_46_bits_nz(wt6_actv_nz[46]),
.io_wt_actv_6_46_bits_data(wt6_actv_data[375:368]),

.io_wt_actv_6_47_valid(wt6_actv_pvld[47]),
.io_wt_actv_6_47_bits_nz(wt6_actv_nz[47]),
.io_wt_actv_6_47_bits_data(wt6_actv_data[383:376]),

.io_wt_actv_6_48_valid(wt6_actv_pvld[48]),
.io_wt_actv_6_48_bits_nz(wt6_actv_nz[48]),
.io_wt_actv_6_48_bits_data(wt6_actv_data[391:384]),

.io_wt_actv_6_49_valid(wt6_actv_pvld[49]),
.io_wt_actv_6_49_bits_nz(wt6_actv_nz[49]),
.io_wt_actv_6_49_bits_data(wt6_actv_data[399:392]),

.io_wt_actv_6_50_valid(wt6_actv_pvld[50]),
.io_wt_actv_6_50_bits_nz(wt6_actv_nz[50]),
.io_wt_actv_6_50_bits_data(wt6_actv_data[407:400]),

.io_wt_actv_6_51_valid(wt6_actv_pvld[51]),
.io_wt_actv_6_51_bits_nz(wt6_actv_nz[51]),
.io_wt_actv_6_51_bits_data(wt6_actv_data[415:408]),

.io_wt_actv_6_52_valid(wt6_actv_pvld[52]),
.io_wt_actv_6_52_bits_nz(wt6_actv_nz[52]),
.io_wt_actv_6_52_bits_data(wt6_actv_data[423:416]),

.io_wt_actv_6_53_valid(wt6_actv_pvld[53]),
.io_wt_actv_6_53_bits_nz(wt6_actv_nz[53]),
.io_wt_actv_6_53_bits_data(wt6_actv_data[431:424]),

.io_wt_actv_6_54_valid(wt6_actv_pvld[54]),
.io_wt_actv_6_54_bits_nz(wt6_actv_nz[54]),
.io_wt_actv_6_54_bits_data(wt6_actv_data[439:432]),

.io_wt_actv_6_55_valid(wt6_actv_pvld[55]),
.io_wt_actv_6_55_bits_nz(wt6_actv_nz[55]),
.io_wt_actv_6_55_bits_data(wt6_actv_data[447:440]),

.io_wt_actv_6_56_valid(wt6_actv_pvld[56]),
.io_wt_actv_6_56_bits_nz(wt6_actv_nz[56]),
.io_wt_actv_6_56_bits_data(wt6_actv_data[455:448]),

.io_wt_actv_6_57_valid(wt6_actv_pvld[57]),
.io_wt_actv_6_57_bits_nz(wt6_actv_nz[57]),
.io_wt_actv_6_57_bits_data(wt6_actv_data[463:456]),

.io_wt_actv_6_58_valid(wt6_actv_pvld[58]),
.io_wt_actv_6_58_bits_nz(wt6_actv_nz[58]),
.io_wt_actv_6_58_bits_data(wt6_actv_data[471:464]),

.io_wt_actv_6_59_valid(wt6_actv_pvld[59]),
.io_wt_actv_6_59_bits_nz(wt6_actv_nz[59]),
.io_wt_actv_6_59_bits_data(wt6_actv_data[479:472]),

.io_wt_actv_6_60_valid(wt6_actv_pvld[60]),
.io_wt_actv_6_60_bits_nz(wt6_actv_nz[60]),
.io_wt_actv_6_60_bits_data(wt6_actv_data[487:480]),

.io_wt_actv_6_61_valid(wt6_actv_pvld[61]),
.io_wt_actv_6_61_bits_nz(wt6_actv_nz[61]),
.io_wt_actv_6_61_bits_data(wt6_actv_data[495:488]),

.io_wt_actv_6_62_valid(wt6_actv_pvld[62]),
.io_wt_actv_6_62_bits_nz(wt6_actv_nz[62]),
.io_wt_actv_6_62_bits_data(wt6_actv_data[503:496]),

.io_wt_actv_6_63_valid(wt6_actv_pvld[63]),
.io_wt_actv_6_63_bits_nz(wt6_actv_nz[63]),
.io_wt_actv_6_63_bits_data(wt6_actv_data[511:504]),

.io_wt_actv_7_0_valid(wt7_actv_pvld[0]),
.io_wt_actv_7_0_bits_nz(wt7_actv_nz[0]),
.io_wt_actv_7_0_bits_data(wt7_actv_data[7:0]),

.io_wt_actv_7_1_valid(wt7_actv_pvld[1]),
.io_wt_actv_7_1_bits_nz(wt7_actv_nz[1]),
.io_wt_actv_7_1_bits_data(wt7_actv_data[15:8]),

.io_wt_actv_7_2_valid(wt7_actv_pvld[2]),
.io_wt_actv_7_2_bits_nz(wt7_actv_nz[2]),
.io_wt_actv_7_2_bits_data(wt7_actv_data[23:16]),

.io_wt_actv_7_3_valid(wt7_actv_pvld[3]),
.io_wt_actv_7_3_bits_nz(wt7_actv_nz[3]),
.io_wt_actv_7_3_bits_data(wt7_actv_data[31:24]),

.io_wt_actv_7_4_valid(wt7_actv_pvld[4]),
.io_wt_actv_7_4_bits_nz(wt7_actv_nz[4]),
.io_wt_actv_7_4_bits_data(wt7_actv_data[39:32]),

.io_wt_actv_7_5_valid(wt7_actv_pvld[5]),
.io_wt_actv_7_5_bits_nz(wt7_actv_nz[5]),
.io_wt_actv_7_5_bits_data(wt7_actv_data[47:40]),

.io_wt_actv_7_6_valid(wt7_actv_pvld[6]),
.io_wt_actv_7_6_bits_nz(wt7_actv_nz[6]),
.io_wt_actv_7_6_bits_data(wt7_actv_data[55:48]),

.io_wt_actv_7_7_valid(wt7_actv_pvld[7]),
.io_wt_actv_7_7_bits_nz(wt7_actv_nz[7]),
.io_wt_actv_7_7_bits_data(wt7_actv_data[63:56]),

.io_wt_actv_7_8_valid(wt7_actv_pvld[8]),
.io_wt_actv_7_8_bits_nz(wt7_actv_nz[8]),
.io_wt_actv_7_8_bits_data(wt7_actv_data[71:64]),

.io_wt_actv_7_9_valid(wt7_actv_pvld[9]),
.io_wt_actv_7_9_bits_nz(wt7_actv_nz[9]),
.io_wt_actv_7_9_bits_data(wt7_actv_data[79:72]),

.io_wt_actv_7_10_valid(wt7_actv_pvld[10]),
.io_wt_actv_7_10_bits_nz(wt7_actv_nz[10]),
.io_wt_actv_7_10_bits_data(wt7_actv_data[87:80]),

.io_wt_actv_7_11_valid(wt7_actv_pvld[11]),
.io_wt_actv_7_11_bits_nz(wt7_actv_nz[11]),
.io_wt_actv_7_11_bits_data(wt7_actv_data[95:88]),

.io_wt_actv_7_12_valid(wt7_actv_pvld[12]),
.io_wt_actv_7_12_bits_nz(wt7_actv_nz[12]),
.io_wt_actv_7_12_bits_data(wt7_actv_data[103:96]),

.io_wt_actv_7_13_valid(wt7_actv_pvld[13]),
.io_wt_actv_7_13_bits_nz(wt7_actv_nz[13]),
.io_wt_actv_7_13_bits_data(wt7_actv_data[111:104]),

.io_wt_actv_7_14_valid(wt7_actv_pvld[14]),
.io_wt_actv_7_14_bits_nz(wt7_actv_nz[14]),
.io_wt_actv_7_14_bits_data(wt7_actv_data[119:112]),

.io_wt_actv_7_15_valid(wt7_actv_pvld[15]),
.io_wt_actv_7_15_bits_nz(wt7_actv_nz[15]),
.io_wt_actv_7_15_bits_data(wt7_actv_data[127:120]),

.io_wt_actv_7_16_valid(wt7_actv_pvld[16]),
.io_wt_actv_7_16_bits_nz(wt7_actv_nz[16]),
.io_wt_actv_7_16_bits_data(wt7_actv_data[135:128]),

.io_wt_actv_7_17_valid(wt7_actv_pvld[17]),
.io_wt_actv_7_17_bits_nz(wt7_actv_nz[17]),
.io_wt_actv_7_17_bits_data(wt7_actv_data[143:136]),

.io_wt_actv_7_18_valid(wt7_actv_pvld[18]),
.io_wt_actv_7_18_bits_nz(wt7_actv_nz[18]),
.io_wt_actv_7_18_bits_data(wt7_actv_data[151:144]),

.io_wt_actv_7_19_valid(wt7_actv_pvld[19]),
.io_wt_actv_7_19_bits_nz(wt7_actv_nz[19]),
.io_wt_actv_7_19_bits_data(wt7_actv_data[159:152]),

.io_wt_actv_7_20_valid(wt7_actv_pvld[20]),
.io_wt_actv_7_20_bits_nz(wt7_actv_nz[20]),
.io_wt_actv_7_20_bits_data(wt7_actv_data[167:160]),

.io_wt_actv_7_21_valid(wt7_actv_pvld[21]),
.io_wt_actv_7_21_bits_nz(wt7_actv_nz[21]),
.io_wt_actv_7_21_bits_data(wt7_actv_data[175:168]),

.io_wt_actv_7_22_valid(wt7_actv_pvld[22]),
.io_wt_actv_7_22_bits_nz(wt7_actv_nz[22]),
.io_wt_actv_7_22_bits_data(wt7_actv_data[183:176]),

.io_wt_actv_7_23_valid(wt7_actv_pvld[23]),
.io_wt_actv_7_23_bits_nz(wt7_actv_nz[23]),
.io_wt_actv_7_23_bits_data(wt7_actv_data[191:184]),

.io_wt_actv_7_24_valid(wt7_actv_pvld[24]),
.io_wt_actv_7_24_bits_nz(wt7_actv_nz[24]),
.io_wt_actv_7_24_bits_data(wt7_actv_data[199:192]),

.io_wt_actv_7_25_valid(wt7_actv_pvld[25]),
.io_wt_actv_7_25_bits_nz(wt7_actv_nz[25]),
.io_wt_actv_7_25_bits_data(wt7_actv_data[207:200]),

.io_wt_actv_7_26_valid(wt7_actv_pvld[26]),
.io_wt_actv_7_26_bits_nz(wt7_actv_nz[26]),
.io_wt_actv_7_26_bits_data(wt7_actv_data[215:208]),

.io_wt_actv_7_27_valid(wt7_actv_pvld[27]),
.io_wt_actv_7_27_bits_nz(wt7_actv_nz[27]),
.io_wt_actv_7_27_bits_data(wt7_actv_data[223:216]),

.io_wt_actv_7_28_valid(wt7_actv_pvld[28]),
.io_wt_actv_7_28_bits_nz(wt7_actv_nz[28]),
.io_wt_actv_7_28_bits_data(wt7_actv_data[231:224]),

.io_wt_actv_7_29_valid(wt7_actv_pvld[29]),
.io_wt_actv_7_29_bits_nz(wt7_actv_nz[29]),
.io_wt_actv_7_29_bits_data(wt7_actv_data[239:232]),

.io_wt_actv_7_30_valid(wt7_actv_pvld[30]),
.io_wt_actv_7_30_bits_nz(wt7_actv_nz[30]),
.io_wt_actv_7_30_bits_data(wt7_actv_data[247:240]),

.io_wt_actv_7_31_valid(wt7_actv_pvld[31]),
.io_wt_actv_7_31_bits_nz(wt7_actv_nz[31]),
.io_wt_actv_7_31_bits_data(wt7_actv_data[255:248]),

.io_wt_actv_7_32_valid(wt7_actv_pvld[32]),
.io_wt_actv_7_32_bits_nz(wt7_actv_nz[32]),
.io_wt_actv_7_32_bits_data(wt7_actv_data[263:256]),

.io_wt_actv_7_33_valid(wt7_actv_pvld[33]),
.io_wt_actv_7_33_bits_nz(wt7_actv_nz[33]),
.io_wt_actv_7_33_bits_data(wt7_actv_data[271:264]),

.io_wt_actv_7_34_valid(wt7_actv_pvld[34]),
.io_wt_actv_7_34_bits_nz(wt7_actv_nz[34]),
.io_wt_actv_7_34_bits_data(wt7_actv_data[279:272]),

.io_wt_actv_7_35_valid(wt7_actv_pvld[35]),
.io_wt_actv_7_35_bits_nz(wt7_actv_nz[35]),
.io_wt_actv_7_35_bits_data(wt7_actv_data[287:280]),

.io_wt_actv_7_36_valid(wt7_actv_pvld[36]),
.io_wt_actv_7_36_bits_nz(wt7_actv_nz[36]),
.io_wt_actv_7_36_bits_data(wt7_actv_data[295:288]),

.io_wt_actv_7_37_valid(wt7_actv_pvld[37]),
.io_wt_actv_7_37_bits_nz(wt7_actv_nz[37]),
.io_wt_actv_7_37_bits_data(wt7_actv_data[303:296]),

.io_wt_actv_7_38_valid(wt7_actv_pvld[38]),
.io_wt_actv_7_38_bits_nz(wt7_actv_nz[38]),
.io_wt_actv_7_38_bits_data(wt7_actv_data[311:304]),

.io_wt_actv_7_39_valid(wt7_actv_pvld[39]),
.io_wt_actv_7_39_bits_nz(wt7_actv_nz[39]),
.io_wt_actv_7_39_bits_data(wt7_actv_data[319:312]),

.io_wt_actv_7_40_valid(wt7_actv_pvld[40]),
.io_wt_actv_7_40_bits_nz(wt7_actv_nz[40]),
.io_wt_actv_7_40_bits_data(wt7_actv_data[327:320]),

.io_wt_actv_7_41_valid(wt7_actv_pvld[41]),
.io_wt_actv_7_41_bits_nz(wt7_actv_nz[41]),
.io_wt_actv_7_41_bits_data(wt7_actv_data[335:328]),

.io_wt_actv_7_42_valid(wt7_actv_pvld[42]),
.io_wt_actv_7_42_bits_nz(wt7_actv_nz[42]),
.io_wt_actv_7_42_bits_data(wt7_actv_data[343:336]),

.io_wt_actv_7_43_valid(wt7_actv_pvld[43]),
.io_wt_actv_7_43_bits_nz(wt7_actv_nz[43]),
.io_wt_actv_7_43_bits_data(wt7_actv_data[351:344]),

.io_wt_actv_7_44_valid(wt7_actv_pvld[44]),
.io_wt_actv_7_44_bits_nz(wt7_actv_nz[44]),
.io_wt_actv_7_44_bits_data(wt7_actv_data[359:352]),

.io_wt_actv_7_45_valid(wt7_actv_pvld[45]),
.io_wt_actv_7_45_bits_nz(wt7_actv_nz[45]),
.io_wt_actv_7_45_bits_data(wt7_actv_data[367:360]),

.io_wt_actv_7_46_valid(wt7_actv_pvld[46]),
.io_wt_actv_7_46_bits_nz(wt7_actv_nz[46]),
.io_wt_actv_7_46_bits_data(wt7_actv_data[375:368]),

.io_wt_actv_7_47_valid(wt7_actv_pvld[47]),
.io_wt_actv_7_47_bits_nz(wt7_actv_nz[47]),
.io_wt_actv_7_47_bits_data(wt7_actv_data[383:376]),

.io_wt_actv_7_48_valid(wt7_actv_pvld[48]),
.io_wt_actv_7_48_bits_nz(wt7_actv_nz[48]),
.io_wt_actv_7_48_bits_data(wt7_actv_data[391:384]),

.io_wt_actv_7_49_valid(wt7_actv_pvld[49]),
.io_wt_actv_7_49_bits_nz(wt7_actv_nz[49]),
.io_wt_actv_7_49_bits_data(wt7_actv_data[399:392]),

.io_wt_actv_7_50_valid(wt7_actv_pvld[50]),
.io_wt_actv_7_50_bits_nz(wt7_actv_nz[50]),
.io_wt_actv_7_50_bits_data(wt7_actv_data[407:400]),

.io_wt_actv_7_51_valid(wt7_actv_pvld[51]),
.io_wt_actv_7_51_bits_nz(wt7_actv_nz[51]),
.io_wt_actv_7_51_bits_data(wt7_actv_data[415:408]),

.io_wt_actv_7_52_valid(wt7_actv_pvld[52]),
.io_wt_actv_7_52_bits_nz(wt7_actv_nz[52]),
.io_wt_actv_7_52_bits_data(wt7_actv_data[423:416]),

.io_wt_actv_7_53_valid(wt7_actv_pvld[53]),
.io_wt_actv_7_53_bits_nz(wt7_actv_nz[53]),
.io_wt_actv_7_53_bits_data(wt7_actv_data[431:424]),

.io_wt_actv_7_54_valid(wt7_actv_pvld[54]),
.io_wt_actv_7_54_bits_nz(wt7_actv_nz[54]),
.io_wt_actv_7_54_bits_data(wt7_actv_data[439:432]),

.io_wt_actv_7_55_valid(wt7_actv_pvld[55]),
.io_wt_actv_7_55_bits_nz(wt7_actv_nz[55]),
.io_wt_actv_7_55_bits_data(wt7_actv_data[447:440]),

.io_wt_actv_7_56_valid(wt7_actv_pvld[56]),
.io_wt_actv_7_56_bits_nz(wt7_actv_nz[56]),
.io_wt_actv_7_56_bits_data(wt7_actv_data[455:448]),

.io_wt_actv_7_57_valid(wt7_actv_pvld[57]),
.io_wt_actv_7_57_bits_nz(wt7_actv_nz[57]),
.io_wt_actv_7_57_bits_data(wt7_actv_data[463:456]),

.io_wt_actv_7_58_valid(wt7_actv_pvld[58]),
.io_wt_actv_7_58_bits_nz(wt7_actv_nz[58]),
.io_wt_actv_7_58_bits_data(wt7_actv_data[471:464]),

.io_wt_actv_7_59_valid(wt7_actv_pvld[59]),
.io_wt_actv_7_59_bits_nz(wt7_actv_nz[59]),
.io_wt_actv_7_59_bits_data(wt7_actv_data[479:472]),

.io_wt_actv_7_60_valid(wt7_actv_pvld[60]),
.io_wt_actv_7_60_bits_nz(wt7_actv_nz[60]),
.io_wt_actv_7_60_bits_data(wt7_actv_data[487:480]),

.io_wt_actv_7_61_valid(wt7_actv_pvld[61]),
.io_wt_actv_7_61_bits_nz(wt7_actv_nz[61]),
.io_wt_actv_7_61_bits_data(wt7_actv_data[495:488]),

.io_wt_actv_7_62_valid(wt7_actv_pvld[62]),
.io_wt_actv_7_62_bits_nz(wt7_actv_nz[62]),
.io_wt_actv_7_62_bits_data(wt7_actv_data[503:496]),

.io_wt_actv_7_63_valid(wt7_actv_pvld[63]),
.io_wt_actv_7_63_bits_nz(wt7_actv_nz[63]),
.io_wt_actv_7_63_bits_data(wt7_actv_data[511:504]),

.io_wt_actv_8_0_valid(wt8_actv_pvld[0]),
.io_wt_actv_8_0_bits_nz(wt8_actv_nz[0]),
.io_wt_actv_8_0_bits_data(wt8_actv_data[7:0]),

.io_wt_actv_8_1_valid(wt8_actv_pvld[1]),
.io_wt_actv_8_1_bits_nz(wt8_actv_nz[1]),
.io_wt_actv_8_1_bits_data(wt8_actv_data[15:8]),

.io_wt_actv_8_2_valid(wt8_actv_pvld[2]),
.io_wt_actv_8_2_bits_nz(wt8_actv_nz[2]),
.io_wt_actv_8_2_bits_data(wt8_actv_data[23:16]),

.io_wt_actv_8_3_valid(wt8_actv_pvld[3]),
.io_wt_actv_8_3_bits_nz(wt8_actv_nz[3]),
.io_wt_actv_8_3_bits_data(wt8_actv_data[31:24]),

.io_wt_actv_8_4_valid(wt8_actv_pvld[4]),
.io_wt_actv_8_4_bits_nz(wt8_actv_nz[4]),
.io_wt_actv_8_4_bits_data(wt8_actv_data[39:32]),

.io_wt_actv_8_5_valid(wt8_actv_pvld[5]),
.io_wt_actv_8_5_bits_nz(wt8_actv_nz[5]),
.io_wt_actv_8_5_bits_data(wt8_actv_data[47:40]),

.io_wt_actv_8_6_valid(wt8_actv_pvld[6]),
.io_wt_actv_8_6_bits_nz(wt8_actv_nz[6]),
.io_wt_actv_8_6_bits_data(wt8_actv_data[55:48]),

.io_wt_actv_8_7_valid(wt8_actv_pvld[7]),
.io_wt_actv_8_7_bits_nz(wt8_actv_nz[7]),
.io_wt_actv_8_7_bits_data(wt8_actv_data[63:56]),

.io_wt_actv_8_8_valid(wt8_actv_pvld[8]),
.io_wt_actv_8_8_bits_nz(wt8_actv_nz[8]),
.io_wt_actv_8_8_bits_data(wt8_actv_data[71:64]),

.io_wt_actv_8_9_valid(wt8_actv_pvld[9]),
.io_wt_actv_8_9_bits_nz(wt8_actv_nz[9]),
.io_wt_actv_8_9_bits_data(wt8_actv_data[79:72]),

.io_wt_actv_8_10_valid(wt8_actv_pvld[10]),
.io_wt_actv_8_10_bits_nz(wt8_actv_nz[10]),
.io_wt_actv_8_10_bits_data(wt8_actv_data[87:80]),

.io_wt_actv_8_11_valid(wt8_actv_pvld[11]),
.io_wt_actv_8_11_bits_nz(wt8_actv_nz[11]),
.io_wt_actv_8_11_bits_data(wt8_actv_data[95:88]),

.io_wt_actv_8_12_valid(wt8_actv_pvld[12]),
.io_wt_actv_8_12_bits_nz(wt8_actv_nz[12]),
.io_wt_actv_8_12_bits_data(wt8_actv_data[103:96]),

.io_wt_actv_8_13_valid(wt8_actv_pvld[13]),
.io_wt_actv_8_13_bits_nz(wt8_actv_nz[13]),
.io_wt_actv_8_13_bits_data(wt8_actv_data[111:104]),

.io_wt_actv_8_14_valid(wt8_actv_pvld[14]),
.io_wt_actv_8_14_bits_nz(wt8_actv_nz[14]),
.io_wt_actv_8_14_bits_data(wt8_actv_data[119:112]),

.io_wt_actv_8_15_valid(wt8_actv_pvld[15]),
.io_wt_actv_8_15_bits_nz(wt8_actv_nz[15]),
.io_wt_actv_8_15_bits_data(wt8_actv_data[127:120]),

.io_wt_actv_8_16_valid(wt8_actv_pvld[16]),
.io_wt_actv_8_16_bits_nz(wt8_actv_nz[16]),
.io_wt_actv_8_16_bits_data(wt8_actv_data[135:128]),

.io_wt_actv_8_17_valid(wt8_actv_pvld[17]),
.io_wt_actv_8_17_bits_nz(wt8_actv_nz[17]),
.io_wt_actv_8_17_bits_data(wt8_actv_data[143:136]),

.io_wt_actv_8_18_valid(wt8_actv_pvld[18]),
.io_wt_actv_8_18_bits_nz(wt8_actv_nz[18]),
.io_wt_actv_8_18_bits_data(wt8_actv_data[151:144]),

.io_wt_actv_8_19_valid(wt8_actv_pvld[19]),
.io_wt_actv_8_19_bits_nz(wt8_actv_nz[19]),
.io_wt_actv_8_19_bits_data(wt8_actv_data[159:152]),

.io_wt_actv_8_20_valid(wt8_actv_pvld[20]),
.io_wt_actv_8_20_bits_nz(wt8_actv_nz[20]),
.io_wt_actv_8_20_bits_data(wt8_actv_data[167:160]),

.io_wt_actv_8_21_valid(wt8_actv_pvld[21]),
.io_wt_actv_8_21_bits_nz(wt8_actv_nz[21]),
.io_wt_actv_8_21_bits_data(wt8_actv_data[175:168]),

.io_wt_actv_8_22_valid(wt8_actv_pvld[22]),
.io_wt_actv_8_22_bits_nz(wt8_actv_nz[22]),
.io_wt_actv_8_22_bits_data(wt8_actv_data[183:176]),

.io_wt_actv_8_23_valid(wt8_actv_pvld[23]),
.io_wt_actv_8_23_bits_nz(wt8_actv_nz[23]),
.io_wt_actv_8_23_bits_data(wt8_actv_data[191:184]),

.io_wt_actv_8_24_valid(wt8_actv_pvld[24]),
.io_wt_actv_8_24_bits_nz(wt8_actv_nz[24]),
.io_wt_actv_8_24_bits_data(wt8_actv_data[199:192]),

.io_wt_actv_8_25_valid(wt8_actv_pvld[25]),
.io_wt_actv_8_25_bits_nz(wt8_actv_nz[25]),
.io_wt_actv_8_25_bits_data(wt8_actv_data[207:200]),

.io_wt_actv_8_26_valid(wt8_actv_pvld[26]),
.io_wt_actv_8_26_bits_nz(wt8_actv_nz[26]),
.io_wt_actv_8_26_bits_data(wt8_actv_data[215:208]),

.io_wt_actv_8_27_valid(wt8_actv_pvld[27]),
.io_wt_actv_8_27_bits_nz(wt8_actv_nz[27]),
.io_wt_actv_8_27_bits_data(wt8_actv_data[223:216]),

.io_wt_actv_8_28_valid(wt8_actv_pvld[28]),
.io_wt_actv_8_28_bits_nz(wt8_actv_nz[28]),
.io_wt_actv_8_28_bits_data(wt8_actv_data[231:224]),

.io_wt_actv_8_29_valid(wt8_actv_pvld[29]),
.io_wt_actv_8_29_bits_nz(wt8_actv_nz[29]),
.io_wt_actv_8_29_bits_data(wt8_actv_data[239:232]),

.io_wt_actv_8_30_valid(wt8_actv_pvld[30]),
.io_wt_actv_8_30_bits_nz(wt8_actv_nz[30]),
.io_wt_actv_8_30_bits_data(wt8_actv_data[247:240]),

.io_wt_actv_8_31_valid(wt8_actv_pvld[31]),
.io_wt_actv_8_31_bits_nz(wt8_actv_nz[31]),
.io_wt_actv_8_31_bits_data(wt8_actv_data[255:248]),

.io_wt_actv_8_32_valid(wt8_actv_pvld[32]),
.io_wt_actv_8_32_bits_nz(wt8_actv_nz[32]),
.io_wt_actv_8_32_bits_data(wt8_actv_data[263:256]),

.io_wt_actv_8_33_valid(wt8_actv_pvld[33]),
.io_wt_actv_8_33_bits_nz(wt8_actv_nz[33]),
.io_wt_actv_8_33_bits_data(wt8_actv_data[271:264]),

.io_wt_actv_8_34_valid(wt8_actv_pvld[34]),
.io_wt_actv_8_34_bits_nz(wt8_actv_nz[34]),
.io_wt_actv_8_34_bits_data(wt8_actv_data[279:272]),

.io_wt_actv_8_35_valid(wt8_actv_pvld[35]),
.io_wt_actv_8_35_bits_nz(wt8_actv_nz[35]),
.io_wt_actv_8_35_bits_data(wt8_actv_data[287:280]),

.io_wt_actv_8_36_valid(wt8_actv_pvld[36]),
.io_wt_actv_8_36_bits_nz(wt8_actv_nz[36]),
.io_wt_actv_8_36_bits_data(wt8_actv_data[295:288]),

.io_wt_actv_8_37_valid(wt8_actv_pvld[37]),
.io_wt_actv_8_37_bits_nz(wt8_actv_nz[37]),
.io_wt_actv_8_37_bits_data(wt8_actv_data[303:296]),

.io_wt_actv_8_38_valid(wt8_actv_pvld[38]),
.io_wt_actv_8_38_bits_nz(wt8_actv_nz[38]),
.io_wt_actv_8_38_bits_data(wt8_actv_data[311:304]),

.io_wt_actv_8_39_valid(wt8_actv_pvld[39]),
.io_wt_actv_8_39_bits_nz(wt8_actv_nz[39]),
.io_wt_actv_8_39_bits_data(wt8_actv_data[319:312]),

.io_wt_actv_8_40_valid(wt8_actv_pvld[40]),
.io_wt_actv_8_40_bits_nz(wt8_actv_nz[40]),
.io_wt_actv_8_40_bits_data(wt8_actv_data[327:320]),

.io_wt_actv_8_41_valid(wt8_actv_pvld[41]),
.io_wt_actv_8_41_bits_nz(wt8_actv_nz[41]),
.io_wt_actv_8_41_bits_data(wt8_actv_data[335:328]),

.io_wt_actv_8_42_valid(wt8_actv_pvld[42]),
.io_wt_actv_8_42_bits_nz(wt8_actv_nz[42]),
.io_wt_actv_8_42_bits_data(wt8_actv_data[343:336]),

.io_wt_actv_8_43_valid(wt8_actv_pvld[43]),
.io_wt_actv_8_43_bits_nz(wt8_actv_nz[43]),
.io_wt_actv_8_43_bits_data(wt8_actv_data[351:344]),

.io_wt_actv_8_44_valid(wt8_actv_pvld[44]),
.io_wt_actv_8_44_bits_nz(wt8_actv_nz[44]),
.io_wt_actv_8_44_bits_data(wt8_actv_data[359:352]),

.io_wt_actv_8_45_valid(wt8_actv_pvld[45]),
.io_wt_actv_8_45_bits_nz(wt8_actv_nz[45]),
.io_wt_actv_8_45_bits_data(wt8_actv_data[367:360]),

.io_wt_actv_8_46_valid(wt8_actv_pvld[46]),
.io_wt_actv_8_46_bits_nz(wt8_actv_nz[46]),
.io_wt_actv_8_46_bits_data(wt8_actv_data[375:368]),

.io_wt_actv_8_47_valid(wt8_actv_pvld[47]),
.io_wt_actv_8_47_bits_nz(wt8_actv_nz[47]),
.io_wt_actv_8_47_bits_data(wt8_actv_data[383:376]),

.io_wt_actv_8_48_valid(wt8_actv_pvld[48]),
.io_wt_actv_8_48_bits_nz(wt8_actv_nz[48]),
.io_wt_actv_8_48_bits_data(wt8_actv_data[391:384]),

.io_wt_actv_8_49_valid(wt8_actv_pvld[49]),
.io_wt_actv_8_49_bits_nz(wt8_actv_nz[49]),
.io_wt_actv_8_49_bits_data(wt8_actv_data[399:392]),

.io_wt_actv_8_50_valid(wt8_actv_pvld[50]),
.io_wt_actv_8_50_bits_nz(wt8_actv_nz[50]),
.io_wt_actv_8_50_bits_data(wt8_actv_data[407:400]),

.io_wt_actv_8_51_valid(wt8_actv_pvld[51]),
.io_wt_actv_8_51_bits_nz(wt8_actv_nz[51]),
.io_wt_actv_8_51_bits_data(wt8_actv_data[415:408]),

.io_wt_actv_8_52_valid(wt8_actv_pvld[52]),
.io_wt_actv_8_52_bits_nz(wt8_actv_nz[52]),
.io_wt_actv_8_52_bits_data(wt8_actv_data[423:416]),

.io_wt_actv_8_53_valid(wt8_actv_pvld[53]),
.io_wt_actv_8_53_bits_nz(wt8_actv_nz[53]),
.io_wt_actv_8_53_bits_data(wt8_actv_data[431:424]),

.io_wt_actv_8_54_valid(wt8_actv_pvld[54]),
.io_wt_actv_8_54_bits_nz(wt8_actv_nz[54]),
.io_wt_actv_8_54_bits_data(wt8_actv_data[439:432]),

.io_wt_actv_8_55_valid(wt8_actv_pvld[55]),
.io_wt_actv_8_55_bits_nz(wt8_actv_nz[55]),
.io_wt_actv_8_55_bits_data(wt8_actv_data[447:440]),

.io_wt_actv_8_56_valid(wt8_actv_pvld[56]),
.io_wt_actv_8_56_bits_nz(wt8_actv_nz[56]),
.io_wt_actv_8_56_bits_data(wt8_actv_data[455:448]),

.io_wt_actv_8_57_valid(wt8_actv_pvld[57]),
.io_wt_actv_8_57_bits_nz(wt8_actv_nz[57]),
.io_wt_actv_8_57_bits_data(wt8_actv_data[463:456]),

.io_wt_actv_8_58_valid(wt8_actv_pvld[58]),
.io_wt_actv_8_58_bits_nz(wt8_actv_nz[58]),
.io_wt_actv_8_58_bits_data(wt8_actv_data[471:464]),

.io_wt_actv_8_59_valid(wt8_actv_pvld[59]),
.io_wt_actv_8_59_bits_nz(wt8_actv_nz[59]),
.io_wt_actv_8_59_bits_data(wt8_actv_data[479:472]),

.io_wt_actv_8_60_valid(wt8_actv_pvld[60]),
.io_wt_actv_8_60_bits_nz(wt8_actv_nz[60]),
.io_wt_actv_8_60_bits_data(wt8_actv_data[487:480]),

.io_wt_actv_8_61_valid(wt8_actv_pvld[61]),
.io_wt_actv_8_61_bits_nz(wt8_actv_nz[61]),
.io_wt_actv_8_61_bits_data(wt8_actv_data[495:488]),

.io_wt_actv_8_62_valid(wt8_actv_pvld[62]),
.io_wt_actv_8_62_bits_nz(wt8_actv_nz[62]),
.io_wt_actv_8_62_bits_data(wt8_actv_data[503:496]),

.io_wt_actv_8_63_valid(wt8_actv_pvld[63]),
.io_wt_actv_8_63_bits_nz(wt8_actv_nz[63]),
.io_wt_actv_8_63_bits_data(wt8_actv_data[511:504]),

.io_wt_actv_9_0_valid(wt9_actv_pvld[0]),
.io_wt_actv_9_0_bits_nz(wt9_actv_nz[0]),
.io_wt_actv_9_0_bits_data(wt9_actv_data[7:0]),

.io_wt_actv_9_1_valid(wt9_actv_pvld[1]),
.io_wt_actv_9_1_bits_nz(wt9_actv_nz[1]),
.io_wt_actv_9_1_bits_data(wt9_actv_data[15:8]),

.io_wt_actv_9_2_valid(wt9_actv_pvld[2]),
.io_wt_actv_9_2_bits_nz(wt9_actv_nz[2]),
.io_wt_actv_9_2_bits_data(wt9_actv_data[23:16]),

.io_wt_actv_9_3_valid(wt9_actv_pvld[3]),
.io_wt_actv_9_3_bits_nz(wt9_actv_nz[3]),
.io_wt_actv_9_3_bits_data(wt9_actv_data[31:24]),

.io_wt_actv_9_4_valid(wt9_actv_pvld[4]),
.io_wt_actv_9_4_bits_nz(wt9_actv_nz[4]),
.io_wt_actv_9_4_bits_data(wt9_actv_data[39:32]),

.io_wt_actv_9_5_valid(wt9_actv_pvld[5]),
.io_wt_actv_9_5_bits_nz(wt9_actv_nz[5]),
.io_wt_actv_9_5_bits_data(wt9_actv_data[47:40]),

.io_wt_actv_9_6_valid(wt9_actv_pvld[6]),
.io_wt_actv_9_6_bits_nz(wt9_actv_nz[6]),
.io_wt_actv_9_6_bits_data(wt9_actv_data[55:48]),

.io_wt_actv_9_7_valid(wt9_actv_pvld[7]),
.io_wt_actv_9_7_bits_nz(wt9_actv_nz[7]),
.io_wt_actv_9_7_bits_data(wt9_actv_data[63:56]),

.io_wt_actv_9_8_valid(wt9_actv_pvld[8]),
.io_wt_actv_9_8_bits_nz(wt9_actv_nz[8]),
.io_wt_actv_9_8_bits_data(wt9_actv_data[71:64]),

.io_wt_actv_9_9_valid(wt9_actv_pvld[9]),
.io_wt_actv_9_9_bits_nz(wt9_actv_nz[9]),
.io_wt_actv_9_9_bits_data(wt9_actv_data[79:72]),

.io_wt_actv_9_10_valid(wt9_actv_pvld[10]),
.io_wt_actv_9_10_bits_nz(wt9_actv_nz[10]),
.io_wt_actv_9_10_bits_data(wt9_actv_data[87:80]),

.io_wt_actv_9_11_valid(wt9_actv_pvld[11]),
.io_wt_actv_9_11_bits_nz(wt9_actv_nz[11]),
.io_wt_actv_9_11_bits_data(wt9_actv_data[95:88]),

.io_wt_actv_9_12_valid(wt9_actv_pvld[12]),
.io_wt_actv_9_12_bits_nz(wt9_actv_nz[12]),
.io_wt_actv_9_12_bits_data(wt9_actv_data[103:96]),

.io_wt_actv_9_13_valid(wt9_actv_pvld[13]),
.io_wt_actv_9_13_bits_nz(wt9_actv_nz[13]),
.io_wt_actv_9_13_bits_data(wt9_actv_data[111:104]),

.io_wt_actv_9_14_valid(wt9_actv_pvld[14]),
.io_wt_actv_9_14_bits_nz(wt9_actv_nz[14]),
.io_wt_actv_9_14_bits_data(wt9_actv_data[119:112]),

.io_wt_actv_9_15_valid(wt9_actv_pvld[15]),
.io_wt_actv_9_15_bits_nz(wt9_actv_nz[15]),
.io_wt_actv_9_15_bits_data(wt9_actv_data[127:120]),

.io_wt_actv_9_16_valid(wt9_actv_pvld[16]),
.io_wt_actv_9_16_bits_nz(wt9_actv_nz[16]),
.io_wt_actv_9_16_bits_data(wt9_actv_data[135:128]),

.io_wt_actv_9_17_valid(wt9_actv_pvld[17]),
.io_wt_actv_9_17_bits_nz(wt9_actv_nz[17]),
.io_wt_actv_9_17_bits_data(wt9_actv_data[143:136]),

.io_wt_actv_9_18_valid(wt9_actv_pvld[18]),
.io_wt_actv_9_18_bits_nz(wt9_actv_nz[18]),
.io_wt_actv_9_18_bits_data(wt9_actv_data[151:144]),

.io_wt_actv_9_19_valid(wt9_actv_pvld[19]),
.io_wt_actv_9_19_bits_nz(wt9_actv_nz[19]),
.io_wt_actv_9_19_bits_data(wt9_actv_data[159:152]),

.io_wt_actv_9_20_valid(wt9_actv_pvld[20]),
.io_wt_actv_9_20_bits_nz(wt9_actv_nz[20]),
.io_wt_actv_9_20_bits_data(wt9_actv_data[167:160]),

.io_wt_actv_9_21_valid(wt9_actv_pvld[21]),
.io_wt_actv_9_21_bits_nz(wt9_actv_nz[21]),
.io_wt_actv_9_21_bits_data(wt9_actv_data[175:168]),

.io_wt_actv_9_22_valid(wt9_actv_pvld[22]),
.io_wt_actv_9_22_bits_nz(wt9_actv_nz[22]),
.io_wt_actv_9_22_bits_data(wt9_actv_data[183:176]),

.io_wt_actv_9_23_valid(wt9_actv_pvld[23]),
.io_wt_actv_9_23_bits_nz(wt9_actv_nz[23]),
.io_wt_actv_9_23_bits_data(wt9_actv_data[191:184]),

.io_wt_actv_9_24_valid(wt9_actv_pvld[24]),
.io_wt_actv_9_24_bits_nz(wt9_actv_nz[24]),
.io_wt_actv_9_24_bits_data(wt9_actv_data[199:192]),

.io_wt_actv_9_25_valid(wt9_actv_pvld[25]),
.io_wt_actv_9_25_bits_nz(wt9_actv_nz[25]),
.io_wt_actv_9_25_bits_data(wt9_actv_data[207:200]),

.io_wt_actv_9_26_valid(wt9_actv_pvld[26]),
.io_wt_actv_9_26_bits_nz(wt9_actv_nz[26]),
.io_wt_actv_9_26_bits_data(wt9_actv_data[215:208]),

.io_wt_actv_9_27_valid(wt9_actv_pvld[27]),
.io_wt_actv_9_27_bits_nz(wt9_actv_nz[27]),
.io_wt_actv_9_27_bits_data(wt9_actv_data[223:216]),

.io_wt_actv_9_28_valid(wt9_actv_pvld[28]),
.io_wt_actv_9_28_bits_nz(wt9_actv_nz[28]),
.io_wt_actv_9_28_bits_data(wt9_actv_data[231:224]),

.io_wt_actv_9_29_valid(wt9_actv_pvld[29]),
.io_wt_actv_9_29_bits_nz(wt9_actv_nz[29]),
.io_wt_actv_9_29_bits_data(wt9_actv_data[239:232]),

.io_wt_actv_9_30_valid(wt9_actv_pvld[30]),
.io_wt_actv_9_30_bits_nz(wt9_actv_nz[30]),
.io_wt_actv_9_30_bits_data(wt9_actv_data[247:240]),

.io_wt_actv_9_31_valid(wt9_actv_pvld[31]),
.io_wt_actv_9_31_bits_nz(wt9_actv_nz[31]),
.io_wt_actv_9_31_bits_data(wt9_actv_data[255:248]),

.io_wt_actv_9_32_valid(wt9_actv_pvld[32]),
.io_wt_actv_9_32_bits_nz(wt9_actv_nz[32]),
.io_wt_actv_9_32_bits_data(wt9_actv_data[263:256]),

.io_wt_actv_9_33_valid(wt9_actv_pvld[33]),
.io_wt_actv_9_33_bits_nz(wt9_actv_nz[33]),
.io_wt_actv_9_33_bits_data(wt9_actv_data[271:264]),

.io_wt_actv_9_34_valid(wt9_actv_pvld[34]),
.io_wt_actv_9_34_bits_nz(wt9_actv_nz[34]),
.io_wt_actv_9_34_bits_data(wt9_actv_data[279:272]),

.io_wt_actv_9_35_valid(wt9_actv_pvld[35]),
.io_wt_actv_9_35_bits_nz(wt9_actv_nz[35]),
.io_wt_actv_9_35_bits_data(wt9_actv_data[287:280]),

.io_wt_actv_9_36_valid(wt9_actv_pvld[36]),
.io_wt_actv_9_36_bits_nz(wt9_actv_nz[36]),
.io_wt_actv_9_36_bits_data(wt9_actv_data[295:288]),

.io_wt_actv_9_37_valid(wt9_actv_pvld[37]),
.io_wt_actv_9_37_bits_nz(wt9_actv_nz[37]),
.io_wt_actv_9_37_bits_data(wt9_actv_data[303:296]),

.io_wt_actv_9_38_valid(wt9_actv_pvld[38]),
.io_wt_actv_9_38_bits_nz(wt9_actv_nz[38]),
.io_wt_actv_9_38_bits_data(wt9_actv_data[311:304]),

.io_wt_actv_9_39_valid(wt9_actv_pvld[39]),
.io_wt_actv_9_39_bits_nz(wt9_actv_nz[39]),
.io_wt_actv_9_39_bits_data(wt9_actv_data[319:312]),

.io_wt_actv_9_40_valid(wt9_actv_pvld[40]),
.io_wt_actv_9_40_bits_nz(wt9_actv_nz[40]),
.io_wt_actv_9_40_bits_data(wt9_actv_data[327:320]),

.io_wt_actv_9_41_valid(wt9_actv_pvld[41]),
.io_wt_actv_9_41_bits_nz(wt9_actv_nz[41]),
.io_wt_actv_9_41_bits_data(wt9_actv_data[335:328]),

.io_wt_actv_9_42_valid(wt9_actv_pvld[42]),
.io_wt_actv_9_42_bits_nz(wt9_actv_nz[42]),
.io_wt_actv_9_42_bits_data(wt9_actv_data[343:336]),

.io_wt_actv_9_43_valid(wt9_actv_pvld[43]),
.io_wt_actv_9_43_bits_nz(wt9_actv_nz[43]),
.io_wt_actv_9_43_bits_data(wt9_actv_data[351:344]),

.io_wt_actv_9_44_valid(wt9_actv_pvld[44]),
.io_wt_actv_9_44_bits_nz(wt9_actv_nz[44]),
.io_wt_actv_9_44_bits_data(wt9_actv_data[359:352]),

.io_wt_actv_9_45_valid(wt9_actv_pvld[45]),
.io_wt_actv_9_45_bits_nz(wt9_actv_nz[45]),
.io_wt_actv_9_45_bits_data(wt9_actv_data[367:360]),

.io_wt_actv_9_46_valid(wt9_actv_pvld[46]),
.io_wt_actv_9_46_bits_nz(wt9_actv_nz[46]),
.io_wt_actv_9_46_bits_data(wt9_actv_data[375:368]),

.io_wt_actv_9_47_valid(wt9_actv_pvld[47]),
.io_wt_actv_9_47_bits_nz(wt9_actv_nz[47]),
.io_wt_actv_9_47_bits_data(wt9_actv_data[383:376]),

.io_wt_actv_9_48_valid(wt9_actv_pvld[48]),
.io_wt_actv_9_48_bits_nz(wt9_actv_nz[48]),
.io_wt_actv_9_48_bits_data(wt9_actv_data[391:384]),

.io_wt_actv_9_49_valid(wt9_actv_pvld[49]),
.io_wt_actv_9_49_bits_nz(wt9_actv_nz[49]),
.io_wt_actv_9_49_bits_data(wt9_actv_data[399:392]),

.io_wt_actv_9_50_valid(wt9_actv_pvld[50]),
.io_wt_actv_9_50_bits_nz(wt9_actv_nz[50]),
.io_wt_actv_9_50_bits_data(wt9_actv_data[407:400]),

.io_wt_actv_9_51_valid(wt9_actv_pvld[51]),
.io_wt_actv_9_51_bits_nz(wt9_actv_nz[51]),
.io_wt_actv_9_51_bits_data(wt9_actv_data[415:408]),

.io_wt_actv_9_52_valid(wt9_actv_pvld[52]),
.io_wt_actv_9_52_bits_nz(wt9_actv_nz[52]),
.io_wt_actv_9_52_bits_data(wt9_actv_data[423:416]),

.io_wt_actv_9_53_valid(wt9_actv_pvld[53]),
.io_wt_actv_9_53_bits_nz(wt9_actv_nz[53]),
.io_wt_actv_9_53_bits_data(wt9_actv_data[431:424]),

.io_wt_actv_9_54_valid(wt9_actv_pvld[54]),
.io_wt_actv_9_54_bits_nz(wt9_actv_nz[54]),
.io_wt_actv_9_54_bits_data(wt9_actv_data[439:432]),

.io_wt_actv_9_55_valid(wt9_actv_pvld[55]),
.io_wt_actv_9_55_bits_nz(wt9_actv_nz[55]),
.io_wt_actv_9_55_bits_data(wt9_actv_data[447:440]),

.io_wt_actv_9_56_valid(wt9_actv_pvld[56]),
.io_wt_actv_9_56_bits_nz(wt9_actv_nz[56]),
.io_wt_actv_9_56_bits_data(wt9_actv_data[455:448]),

.io_wt_actv_9_57_valid(wt9_actv_pvld[57]),
.io_wt_actv_9_57_bits_nz(wt9_actv_nz[57]),
.io_wt_actv_9_57_bits_data(wt9_actv_data[463:456]),

.io_wt_actv_9_58_valid(wt9_actv_pvld[58]),
.io_wt_actv_9_58_bits_nz(wt9_actv_nz[58]),
.io_wt_actv_9_58_bits_data(wt9_actv_data[471:464]),

.io_wt_actv_9_59_valid(wt9_actv_pvld[59]),
.io_wt_actv_9_59_bits_nz(wt9_actv_nz[59]),
.io_wt_actv_9_59_bits_data(wt9_actv_data[479:472]),

.io_wt_actv_9_60_valid(wt9_actv_pvld[60]),
.io_wt_actv_9_60_bits_nz(wt9_actv_nz[60]),
.io_wt_actv_9_60_bits_data(wt9_actv_data[487:480]),

.io_wt_actv_9_61_valid(wt9_actv_pvld[61]),
.io_wt_actv_9_61_bits_nz(wt9_actv_nz[61]),
.io_wt_actv_9_61_bits_data(wt9_actv_data[495:488]),

.io_wt_actv_9_62_valid(wt9_actv_pvld[62]),
.io_wt_actv_9_62_bits_nz(wt9_actv_nz[62]),
.io_wt_actv_9_62_bits_data(wt9_actv_data[503:496]),

.io_wt_actv_9_63_valid(wt9_actv_pvld[63]),
.io_wt_actv_9_63_bits_nz(wt9_actv_nz[63]),
.io_wt_actv_9_63_bits_data(wt9_actv_data[511:504]),

.io_wt_actv_10_0_valid(wt10_actv_pvld[0]),
.io_wt_actv_10_0_bits_nz(wt10_actv_nz[0]),
.io_wt_actv_10_0_bits_data(wt10_actv_data[7:0]),

.io_wt_actv_10_1_valid(wt10_actv_pvld[1]),
.io_wt_actv_10_1_bits_nz(wt10_actv_nz[1]),
.io_wt_actv_10_1_bits_data(wt10_actv_data[15:8]),

.io_wt_actv_10_2_valid(wt10_actv_pvld[2]),
.io_wt_actv_10_2_bits_nz(wt10_actv_nz[2]),
.io_wt_actv_10_2_bits_data(wt10_actv_data[23:16]),

.io_wt_actv_10_3_valid(wt10_actv_pvld[3]),
.io_wt_actv_10_3_bits_nz(wt10_actv_nz[3]),
.io_wt_actv_10_3_bits_data(wt10_actv_data[31:24]),

.io_wt_actv_10_4_valid(wt10_actv_pvld[4]),
.io_wt_actv_10_4_bits_nz(wt10_actv_nz[4]),
.io_wt_actv_10_4_bits_data(wt10_actv_data[39:32]),

.io_wt_actv_10_5_valid(wt10_actv_pvld[5]),
.io_wt_actv_10_5_bits_nz(wt10_actv_nz[5]),
.io_wt_actv_10_5_bits_data(wt10_actv_data[47:40]),

.io_wt_actv_10_6_valid(wt10_actv_pvld[6]),
.io_wt_actv_10_6_bits_nz(wt10_actv_nz[6]),
.io_wt_actv_10_6_bits_data(wt10_actv_data[55:48]),

.io_wt_actv_10_7_valid(wt10_actv_pvld[7]),
.io_wt_actv_10_7_bits_nz(wt10_actv_nz[7]),
.io_wt_actv_10_7_bits_data(wt10_actv_data[63:56]),

.io_wt_actv_10_8_valid(wt10_actv_pvld[8]),
.io_wt_actv_10_8_bits_nz(wt10_actv_nz[8]),
.io_wt_actv_10_8_bits_data(wt10_actv_data[71:64]),

.io_wt_actv_10_9_valid(wt10_actv_pvld[9]),
.io_wt_actv_10_9_bits_nz(wt10_actv_nz[9]),
.io_wt_actv_10_9_bits_data(wt10_actv_data[79:72]),

.io_wt_actv_10_10_valid(wt10_actv_pvld[10]),
.io_wt_actv_10_10_bits_nz(wt10_actv_nz[10]),
.io_wt_actv_10_10_bits_data(wt10_actv_data[87:80]),

.io_wt_actv_10_11_valid(wt10_actv_pvld[11]),
.io_wt_actv_10_11_bits_nz(wt10_actv_nz[11]),
.io_wt_actv_10_11_bits_data(wt10_actv_data[95:88]),

.io_wt_actv_10_12_valid(wt10_actv_pvld[12]),
.io_wt_actv_10_12_bits_nz(wt10_actv_nz[12]),
.io_wt_actv_10_12_bits_data(wt10_actv_data[103:96]),

.io_wt_actv_10_13_valid(wt10_actv_pvld[13]),
.io_wt_actv_10_13_bits_nz(wt10_actv_nz[13]),
.io_wt_actv_10_13_bits_data(wt10_actv_data[111:104]),

.io_wt_actv_10_14_valid(wt10_actv_pvld[14]),
.io_wt_actv_10_14_bits_nz(wt10_actv_nz[14]),
.io_wt_actv_10_14_bits_data(wt10_actv_data[119:112]),

.io_wt_actv_10_15_valid(wt10_actv_pvld[15]),
.io_wt_actv_10_15_bits_nz(wt10_actv_nz[15]),
.io_wt_actv_10_15_bits_data(wt10_actv_data[127:120]),

.io_wt_actv_10_16_valid(wt10_actv_pvld[16]),
.io_wt_actv_10_16_bits_nz(wt10_actv_nz[16]),
.io_wt_actv_10_16_bits_data(wt10_actv_data[135:128]),

.io_wt_actv_10_17_valid(wt10_actv_pvld[17]),
.io_wt_actv_10_17_bits_nz(wt10_actv_nz[17]),
.io_wt_actv_10_17_bits_data(wt10_actv_data[143:136]),

.io_wt_actv_10_18_valid(wt10_actv_pvld[18]),
.io_wt_actv_10_18_bits_nz(wt10_actv_nz[18]),
.io_wt_actv_10_18_bits_data(wt10_actv_data[151:144]),

.io_wt_actv_10_19_valid(wt10_actv_pvld[19]),
.io_wt_actv_10_19_bits_nz(wt10_actv_nz[19]),
.io_wt_actv_10_19_bits_data(wt10_actv_data[159:152]),

.io_wt_actv_10_20_valid(wt10_actv_pvld[20]),
.io_wt_actv_10_20_bits_nz(wt10_actv_nz[20]),
.io_wt_actv_10_20_bits_data(wt10_actv_data[167:160]),

.io_wt_actv_10_21_valid(wt10_actv_pvld[21]),
.io_wt_actv_10_21_bits_nz(wt10_actv_nz[21]),
.io_wt_actv_10_21_bits_data(wt10_actv_data[175:168]),

.io_wt_actv_10_22_valid(wt10_actv_pvld[22]),
.io_wt_actv_10_22_bits_nz(wt10_actv_nz[22]),
.io_wt_actv_10_22_bits_data(wt10_actv_data[183:176]),

.io_wt_actv_10_23_valid(wt10_actv_pvld[23]),
.io_wt_actv_10_23_bits_nz(wt10_actv_nz[23]),
.io_wt_actv_10_23_bits_data(wt10_actv_data[191:184]),

.io_wt_actv_10_24_valid(wt10_actv_pvld[24]),
.io_wt_actv_10_24_bits_nz(wt10_actv_nz[24]),
.io_wt_actv_10_24_bits_data(wt10_actv_data[199:192]),

.io_wt_actv_10_25_valid(wt10_actv_pvld[25]),
.io_wt_actv_10_25_bits_nz(wt10_actv_nz[25]),
.io_wt_actv_10_25_bits_data(wt10_actv_data[207:200]),

.io_wt_actv_10_26_valid(wt10_actv_pvld[26]),
.io_wt_actv_10_26_bits_nz(wt10_actv_nz[26]),
.io_wt_actv_10_26_bits_data(wt10_actv_data[215:208]),

.io_wt_actv_10_27_valid(wt10_actv_pvld[27]),
.io_wt_actv_10_27_bits_nz(wt10_actv_nz[27]),
.io_wt_actv_10_27_bits_data(wt10_actv_data[223:216]),

.io_wt_actv_10_28_valid(wt10_actv_pvld[28]),
.io_wt_actv_10_28_bits_nz(wt10_actv_nz[28]),
.io_wt_actv_10_28_bits_data(wt10_actv_data[231:224]),

.io_wt_actv_10_29_valid(wt10_actv_pvld[29]),
.io_wt_actv_10_29_bits_nz(wt10_actv_nz[29]),
.io_wt_actv_10_29_bits_data(wt10_actv_data[239:232]),

.io_wt_actv_10_30_valid(wt10_actv_pvld[30]),
.io_wt_actv_10_30_bits_nz(wt10_actv_nz[30]),
.io_wt_actv_10_30_bits_data(wt10_actv_data[247:240]),

.io_wt_actv_10_31_valid(wt10_actv_pvld[31]),
.io_wt_actv_10_31_bits_nz(wt10_actv_nz[31]),
.io_wt_actv_10_31_bits_data(wt10_actv_data[255:248]),

.io_wt_actv_10_32_valid(wt10_actv_pvld[32]),
.io_wt_actv_10_32_bits_nz(wt10_actv_nz[32]),
.io_wt_actv_10_32_bits_data(wt10_actv_data[263:256]),

.io_wt_actv_10_33_valid(wt10_actv_pvld[33]),
.io_wt_actv_10_33_bits_nz(wt10_actv_nz[33]),
.io_wt_actv_10_33_bits_data(wt10_actv_data[271:264]),

.io_wt_actv_10_34_valid(wt10_actv_pvld[34]),
.io_wt_actv_10_34_bits_nz(wt10_actv_nz[34]),
.io_wt_actv_10_34_bits_data(wt10_actv_data[279:272]),

.io_wt_actv_10_35_valid(wt10_actv_pvld[35]),
.io_wt_actv_10_35_bits_nz(wt10_actv_nz[35]),
.io_wt_actv_10_35_bits_data(wt10_actv_data[287:280]),

.io_wt_actv_10_36_valid(wt10_actv_pvld[36]),
.io_wt_actv_10_36_bits_nz(wt10_actv_nz[36]),
.io_wt_actv_10_36_bits_data(wt10_actv_data[295:288]),

.io_wt_actv_10_37_valid(wt10_actv_pvld[37]),
.io_wt_actv_10_37_bits_nz(wt10_actv_nz[37]),
.io_wt_actv_10_37_bits_data(wt10_actv_data[303:296]),

.io_wt_actv_10_38_valid(wt10_actv_pvld[38]),
.io_wt_actv_10_38_bits_nz(wt10_actv_nz[38]),
.io_wt_actv_10_38_bits_data(wt10_actv_data[311:304]),

.io_wt_actv_10_39_valid(wt10_actv_pvld[39]),
.io_wt_actv_10_39_bits_nz(wt10_actv_nz[39]),
.io_wt_actv_10_39_bits_data(wt10_actv_data[319:312]),

.io_wt_actv_10_40_valid(wt10_actv_pvld[40]),
.io_wt_actv_10_40_bits_nz(wt10_actv_nz[40]),
.io_wt_actv_10_40_bits_data(wt10_actv_data[327:320]),

.io_wt_actv_10_41_valid(wt10_actv_pvld[41]),
.io_wt_actv_10_41_bits_nz(wt10_actv_nz[41]),
.io_wt_actv_10_41_bits_data(wt10_actv_data[335:328]),

.io_wt_actv_10_42_valid(wt10_actv_pvld[42]),
.io_wt_actv_10_42_bits_nz(wt10_actv_nz[42]),
.io_wt_actv_10_42_bits_data(wt10_actv_data[343:336]),

.io_wt_actv_10_43_valid(wt10_actv_pvld[43]),
.io_wt_actv_10_43_bits_nz(wt10_actv_nz[43]),
.io_wt_actv_10_43_bits_data(wt10_actv_data[351:344]),

.io_wt_actv_10_44_valid(wt10_actv_pvld[44]),
.io_wt_actv_10_44_bits_nz(wt10_actv_nz[44]),
.io_wt_actv_10_44_bits_data(wt10_actv_data[359:352]),

.io_wt_actv_10_45_valid(wt10_actv_pvld[45]),
.io_wt_actv_10_45_bits_nz(wt10_actv_nz[45]),
.io_wt_actv_10_45_bits_data(wt10_actv_data[367:360]),

.io_wt_actv_10_46_valid(wt10_actv_pvld[46]),
.io_wt_actv_10_46_bits_nz(wt10_actv_nz[46]),
.io_wt_actv_10_46_bits_data(wt10_actv_data[375:368]),

.io_wt_actv_10_47_valid(wt10_actv_pvld[47]),
.io_wt_actv_10_47_bits_nz(wt10_actv_nz[47]),
.io_wt_actv_10_47_bits_data(wt10_actv_data[383:376]),

.io_wt_actv_10_48_valid(wt10_actv_pvld[48]),
.io_wt_actv_10_48_bits_nz(wt10_actv_nz[48]),
.io_wt_actv_10_48_bits_data(wt10_actv_data[391:384]),

.io_wt_actv_10_49_valid(wt10_actv_pvld[49]),
.io_wt_actv_10_49_bits_nz(wt10_actv_nz[49]),
.io_wt_actv_10_49_bits_data(wt10_actv_data[399:392]),

.io_wt_actv_10_50_valid(wt10_actv_pvld[50]),
.io_wt_actv_10_50_bits_nz(wt10_actv_nz[50]),
.io_wt_actv_10_50_bits_data(wt10_actv_data[407:400]),

.io_wt_actv_10_51_valid(wt10_actv_pvld[51]),
.io_wt_actv_10_51_bits_nz(wt10_actv_nz[51]),
.io_wt_actv_10_51_bits_data(wt10_actv_data[415:408]),

.io_wt_actv_10_52_valid(wt10_actv_pvld[52]),
.io_wt_actv_10_52_bits_nz(wt10_actv_nz[52]),
.io_wt_actv_10_52_bits_data(wt10_actv_data[423:416]),

.io_wt_actv_10_53_valid(wt10_actv_pvld[53]),
.io_wt_actv_10_53_bits_nz(wt10_actv_nz[53]),
.io_wt_actv_10_53_bits_data(wt10_actv_data[431:424]),

.io_wt_actv_10_54_valid(wt10_actv_pvld[54]),
.io_wt_actv_10_54_bits_nz(wt10_actv_nz[54]),
.io_wt_actv_10_54_bits_data(wt10_actv_data[439:432]),

.io_wt_actv_10_55_valid(wt10_actv_pvld[55]),
.io_wt_actv_10_55_bits_nz(wt10_actv_nz[55]),
.io_wt_actv_10_55_bits_data(wt10_actv_data[447:440]),

.io_wt_actv_10_56_valid(wt10_actv_pvld[56]),
.io_wt_actv_10_56_bits_nz(wt10_actv_nz[56]),
.io_wt_actv_10_56_bits_data(wt10_actv_data[455:448]),

.io_wt_actv_10_57_valid(wt10_actv_pvld[57]),
.io_wt_actv_10_57_bits_nz(wt10_actv_nz[57]),
.io_wt_actv_10_57_bits_data(wt10_actv_data[463:456]),

.io_wt_actv_10_58_valid(wt10_actv_pvld[58]),
.io_wt_actv_10_58_bits_nz(wt10_actv_nz[58]),
.io_wt_actv_10_58_bits_data(wt10_actv_data[471:464]),

.io_wt_actv_10_59_valid(wt10_actv_pvld[59]),
.io_wt_actv_10_59_bits_nz(wt10_actv_nz[59]),
.io_wt_actv_10_59_bits_data(wt10_actv_data[479:472]),

.io_wt_actv_10_60_valid(wt10_actv_pvld[60]),
.io_wt_actv_10_60_bits_nz(wt10_actv_nz[60]),
.io_wt_actv_10_60_bits_data(wt10_actv_data[487:480]),

.io_wt_actv_10_61_valid(wt10_actv_pvld[61]),
.io_wt_actv_10_61_bits_nz(wt10_actv_nz[61]),
.io_wt_actv_10_61_bits_data(wt10_actv_data[495:488]),

.io_wt_actv_10_62_valid(wt10_actv_pvld[62]),
.io_wt_actv_10_62_bits_nz(wt10_actv_nz[62]),
.io_wt_actv_10_62_bits_data(wt10_actv_data[503:496]),

.io_wt_actv_10_63_valid(wt10_actv_pvld[63]),
.io_wt_actv_10_63_bits_nz(wt10_actv_nz[63]),
.io_wt_actv_10_63_bits_data(wt10_actv_data[511:504]),

.io_wt_actv_11_0_valid(wt11_actv_pvld[0]),
.io_wt_actv_11_0_bits_nz(wt11_actv_nz[0]),
.io_wt_actv_11_0_bits_data(wt11_actv_data[7:0]),

.io_wt_actv_11_1_valid(wt11_actv_pvld[1]),
.io_wt_actv_11_1_bits_nz(wt11_actv_nz[1]),
.io_wt_actv_11_1_bits_data(wt11_actv_data[15:8]),

.io_wt_actv_11_2_valid(wt11_actv_pvld[2]),
.io_wt_actv_11_2_bits_nz(wt11_actv_nz[2]),
.io_wt_actv_11_2_bits_data(wt11_actv_data[23:16]),

.io_wt_actv_11_3_valid(wt11_actv_pvld[3]),
.io_wt_actv_11_3_bits_nz(wt11_actv_nz[3]),
.io_wt_actv_11_3_bits_data(wt11_actv_data[31:24]),

.io_wt_actv_11_4_valid(wt11_actv_pvld[4]),
.io_wt_actv_11_4_bits_nz(wt11_actv_nz[4]),
.io_wt_actv_11_4_bits_data(wt11_actv_data[39:32]),

.io_wt_actv_11_5_valid(wt11_actv_pvld[5]),
.io_wt_actv_11_5_bits_nz(wt11_actv_nz[5]),
.io_wt_actv_11_5_bits_data(wt11_actv_data[47:40]),

.io_wt_actv_11_6_valid(wt11_actv_pvld[6]),
.io_wt_actv_11_6_bits_nz(wt11_actv_nz[6]),
.io_wt_actv_11_6_bits_data(wt11_actv_data[55:48]),

.io_wt_actv_11_7_valid(wt11_actv_pvld[7]),
.io_wt_actv_11_7_bits_nz(wt11_actv_nz[7]),
.io_wt_actv_11_7_bits_data(wt11_actv_data[63:56]),

.io_wt_actv_11_8_valid(wt11_actv_pvld[8]),
.io_wt_actv_11_8_bits_nz(wt11_actv_nz[8]),
.io_wt_actv_11_8_bits_data(wt11_actv_data[71:64]),

.io_wt_actv_11_9_valid(wt11_actv_pvld[9]),
.io_wt_actv_11_9_bits_nz(wt11_actv_nz[9]),
.io_wt_actv_11_9_bits_data(wt11_actv_data[79:72]),

.io_wt_actv_11_10_valid(wt11_actv_pvld[10]),
.io_wt_actv_11_10_bits_nz(wt11_actv_nz[10]),
.io_wt_actv_11_10_bits_data(wt11_actv_data[87:80]),

.io_wt_actv_11_11_valid(wt11_actv_pvld[11]),
.io_wt_actv_11_11_bits_nz(wt11_actv_nz[11]),
.io_wt_actv_11_11_bits_data(wt11_actv_data[95:88]),

.io_wt_actv_11_12_valid(wt11_actv_pvld[12]),
.io_wt_actv_11_12_bits_nz(wt11_actv_nz[12]),
.io_wt_actv_11_12_bits_data(wt11_actv_data[103:96]),

.io_wt_actv_11_13_valid(wt11_actv_pvld[13]),
.io_wt_actv_11_13_bits_nz(wt11_actv_nz[13]),
.io_wt_actv_11_13_bits_data(wt11_actv_data[111:104]),

.io_wt_actv_11_14_valid(wt11_actv_pvld[14]),
.io_wt_actv_11_14_bits_nz(wt11_actv_nz[14]),
.io_wt_actv_11_14_bits_data(wt11_actv_data[119:112]),

.io_wt_actv_11_15_valid(wt11_actv_pvld[15]),
.io_wt_actv_11_15_bits_nz(wt11_actv_nz[15]),
.io_wt_actv_11_15_bits_data(wt11_actv_data[127:120]),

.io_wt_actv_11_16_valid(wt11_actv_pvld[16]),
.io_wt_actv_11_16_bits_nz(wt11_actv_nz[16]),
.io_wt_actv_11_16_bits_data(wt11_actv_data[135:128]),

.io_wt_actv_11_17_valid(wt11_actv_pvld[17]),
.io_wt_actv_11_17_bits_nz(wt11_actv_nz[17]),
.io_wt_actv_11_17_bits_data(wt11_actv_data[143:136]),

.io_wt_actv_11_18_valid(wt11_actv_pvld[18]),
.io_wt_actv_11_18_bits_nz(wt11_actv_nz[18]),
.io_wt_actv_11_18_bits_data(wt11_actv_data[151:144]),

.io_wt_actv_11_19_valid(wt11_actv_pvld[19]),
.io_wt_actv_11_19_bits_nz(wt11_actv_nz[19]),
.io_wt_actv_11_19_bits_data(wt11_actv_data[159:152]),

.io_wt_actv_11_20_valid(wt11_actv_pvld[20]),
.io_wt_actv_11_20_bits_nz(wt11_actv_nz[20]),
.io_wt_actv_11_20_bits_data(wt11_actv_data[167:160]),

.io_wt_actv_11_21_valid(wt11_actv_pvld[21]),
.io_wt_actv_11_21_bits_nz(wt11_actv_nz[21]),
.io_wt_actv_11_21_bits_data(wt11_actv_data[175:168]),

.io_wt_actv_11_22_valid(wt11_actv_pvld[22]),
.io_wt_actv_11_22_bits_nz(wt11_actv_nz[22]),
.io_wt_actv_11_22_bits_data(wt11_actv_data[183:176]),

.io_wt_actv_11_23_valid(wt11_actv_pvld[23]),
.io_wt_actv_11_23_bits_nz(wt11_actv_nz[23]),
.io_wt_actv_11_23_bits_data(wt11_actv_data[191:184]),

.io_wt_actv_11_24_valid(wt11_actv_pvld[24]),
.io_wt_actv_11_24_bits_nz(wt11_actv_nz[24]),
.io_wt_actv_11_24_bits_data(wt11_actv_data[199:192]),

.io_wt_actv_11_25_valid(wt11_actv_pvld[25]),
.io_wt_actv_11_25_bits_nz(wt11_actv_nz[25]),
.io_wt_actv_11_25_bits_data(wt11_actv_data[207:200]),

.io_wt_actv_11_26_valid(wt11_actv_pvld[26]),
.io_wt_actv_11_26_bits_nz(wt11_actv_nz[26]),
.io_wt_actv_11_26_bits_data(wt11_actv_data[215:208]),

.io_wt_actv_11_27_valid(wt11_actv_pvld[27]),
.io_wt_actv_11_27_bits_nz(wt11_actv_nz[27]),
.io_wt_actv_11_27_bits_data(wt11_actv_data[223:216]),

.io_wt_actv_11_28_valid(wt11_actv_pvld[28]),
.io_wt_actv_11_28_bits_nz(wt11_actv_nz[28]),
.io_wt_actv_11_28_bits_data(wt11_actv_data[231:224]),

.io_wt_actv_11_29_valid(wt11_actv_pvld[29]),
.io_wt_actv_11_29_bits_nz(wt11_actv_nz[29]),
.io_wt_actv_11_29_bits_data(wt11_actv_data[239:232]),

.io_wt_actv_11_30_valid(wt11_actv_pvld[30]),
.io_wt_actv_11_30_bits_nz(wt11_actv_nz[30]),
.io_wt_actv_11_30_bits_data(wt11_actv_data[247:240]),

.io_wt_actv_11_31_valid(wt11_actv_pvld[31]),
.io_wt_actv_11_31_bits_nz(wt11_actv_nz[31]),
.io_wt_actv_11_31_bits_data(wt11_actv_data[255:248]),

.io_wt_actv_11_32_valid(wt11_actv_pvld[32]),
.io_wt_actv_11_32_bits_nz(wt11_actv_nz[32]),
.io_wt_actv_11_32_bits_data(wt11_actv_data[263:256]),

.io_wt_actv_11_33_valid(wt11_actv_pvld[33]),
.io_wt_actv_11_33_bits_nz(wt11_actv_nz[33]),
.io_wt_actv_11_33_bits_data(wt11_actv_data[271:264]),

.io_wt_actv_11_34_valid(wt11_actv_pvld[34]),
.io_wt_actv_11_34_bits_nz(wt11_actv_nz[34]),
.io_wt_actv_11_34_bits_data(wt11_actv_data[279:272]),

.io_wt_actv_11_35_valid(wt11_actv_pvld[35]),
.io_wt_actv_11_35_bits_nz(wt11_actv_nz[35]),
.io_wt_actv_11_35_bits_data(wt11_actv_data[287:280]),

.io_wt_actv_11_36_valid(wt11_actv_pvld[36]),
.io_wt_actv_11_36_bits_nz(wt11_actv_nz[36]),
.io_wt_actv_11_36_bits_data(wt11_actv_data[295:288]),

.io_wt_actv_11_37_valid(wt11_actv_pvld[37]),
.io_wt_actv_11_37_bits_nz(wt11_actv_nz[37]),
.io_wt_actv_11_37_bits_data(wt11_actv_data[303:296]),

.io_wt_actv_11_38_valid(wt11_actv_pvld[38]),
.io_wt_actv_11_38_bits_nz(wt11_actv_nz[38]),
.io_wt_actv_11_38_bits_data(wt11_actv_data[311:304]),

.io_wt_actv_11_39_valid(wt11_actv_pvld[39]),
.io_wt_actv_11_39_bits_nz(wt11_actv_nz[39]),
.io_wt_actv_11_39_bits_data(wt11_actv_data[319:312]),

.io_wt_actv_11_40_valid(wt11_actv_pvld[40]),
.io_wt_actv_11_40_bits_nz(wt11_actv_nz[40]),
.io_wt_actv_11_40_bits_data(wt11_actv_data[327:320]),

.io_wt_actv_11_41_valid(wt11_actv_pvld[41]),
.io_wt_actv_11_41_bits_nz(wt11_actv_nz[41]),
.io_wt_actv_11_41_bits_data(wt11_actv_data[335:328]),

.io_wt_actv_11_42_valid(wt11_actv_pvld[42]),
.io_wt_actv_11_42_bits_nz(wt11_actv_nz[42]),
.io_wt_actv_11_42_bits_data(wt11_actv_data[343:336]),

.io_wt_actv_11_43_valid(wt11_actv_pvld[43]),
.io_wt_actv_11_43_bits_nz(wt11_actv_nz[43]),
.io_wt_actv_11_43_bits_data(wt11_actv_data[351:344]),

.io_wt_actv_11_44_valid(wt11_actv_pvld[44]),
.io_wt_actv_11_44_bits_nz(wt11_actv_nz[44]),
.io_wt_actv_11_44_bits_data(wt11_actv_data[359:352]),

.io_wt_actv_11_45_valid(wt11_actv_pvld[45]),
.io_wt_actv_11_45_bits_nz(wt11_actv_nz[45]),
.io_wt_actv_11_45_bits_data(wt11_actv_data[367:360]),

.io_wt_actv_11_46_valid(wt11_actv_pvld[46]),
.io_wt_actv_11_46_bits_nz(wt11_actv_nz[46]),
.io_wt_actv_11_46_bits_data(wt11_actv_data[375:368]),

.io_wt_actv_11_47_valid(wt11_actv_pvld[47]),
.io_wt_actv_11_47_bits_nz(wt11_actv_nz[47]),
.io_wt_actv_11_47_bits_data(wt11_actv_data[383:376]),

.io_wt_actv_11_48_valid(wt11_actv_pvld[48]),
.io_wt_actv_11_48_bits_nz(wt11_actv_nz[48]),
.io_wt_actv_11_48_bits_data(wt11_actv_data[391:384]),

.io_wt_actv_11_49_valid(wt11_actv_pvld[49]),
.io_wt_actv_11_49_bits_nz(wt11_actv_nz[49]),
.io_wt_actv_11_49_bits_data(wt11_actv_data[399:392]),

.io_wt_actv_11_50_valid(wt11_actv_pvld[50]),
.io_wt_actv_11_50_bits_nz(wt11_actv_nz[50]),
.io_wt_actv_11_50_bits_data(wt11_actv_data[407:400]),

.io_wt_actv_11_51_valid(wt11_actv_pvld[51]),
.io_wt_actv_11_51_bits_nz(wt11_actv_nz[51]),
.io_wt_actv_11_51_bits_data(wt11_actv_data[415:408]),

.io_wt_actv_11_52_valid(wt11_actv_pvld[52]),
.io_wt_actv_11_52_bits_nz(wt11_actv_nz[52]),
.io_wt_actv_11_52_bits_data(wt11_actv_data[423:416]),

.io_wt_actv_11_53_valid(wt11_actv_pvld[53]),
.io_wt_actv_11_53_bits_nz(wt11_actv_nz[53]),
.io_wt_actv_11_53_bits_data(wt11_actv_data[431:424]),

.io_wt_actv_11_54_valid(wt11_actv_pvld[54]),
.io_wt_actv_11_54_bits_nz(wt11_actv_nz[54]),
.io_wt_actv_11_54_bits_data(wt11_actv_data[439:432]),

.io_wt_actv_11_55_valid(wt11_actv_pvld[55]),
.io_wt_actv_11_55_bits_nz(wt11_actv_nz[55]),
.io_wt_actv_11_55_bits_data(wt11_actv_data[447:440]),

.io_wt_actv_11_56_valid(wt11_actv_pvld[56]),
.io_wt_actv_11_56_bits_nz(wt11_actv_nz[56]),
.io_wt_actv_11_56_bits_data(wt11_actv_data[455:448]),

.io_wt_actv_11_57_valid(wt11_actv_pvld[57]),
.io_wt_actv_11_57_bits_nz(wt11_actv_nz[57]),
.io_wt_actv_11_57_bits_data(wt11_actv_data[463:456]),

.io_wt_actv_11_58_valid(wt11_actv_pvld[58]),
.io_wt_actv_11_58_bits_nz(wt11_actv_nz[58]),
.io_wt_actv_11_58_bits_data(wt11_actv_data[471:464]),

.io_wt_actv_11_59_valid(wt11_actv_pvld[59]),
.io_wt_actv_11_59_bits_nz(wt11_actv_nz[59]),
.io_wt_actv_11_59_bits_data(wt11_actv_data[479:472]),

.io_wt_actv_11_60_valid(wt11_actv_pvld[60]),
.io_wt_actv_11_60_bits_nz(wt11_actv_nz[60]),
.io_wt_actv_11_60_bits_data(wt11_actv_data[487:480]),

.io_wt_actv_11_61_valid(wt11_actv_pvld[61]),
.io_wt_actv_11_61_bits_nz(wt11_actv_nz[61]),
.io_wt_actv_11_61_bits_data(wt11_actv_data[495:488]),

.io_wt_actv_11_62_valid(wt11_actv_pvld[62]),
.io_wt_actv_11_62_bits_nz(wt11_actv_nz[62]),
.io_wt_actv_11_62_bits_data(wt11_actv_data[503:496]),

.io_wt_actv_11_63_valid(wt11_actv_pvld[63]),
.io_wt_actv_11_63_bits_nz(wt11_actv_nz[63]),
.io_wt_actv_11_63_bits_data(wt11_actv_data[511:504]),

.io_wt_actv_12_0_valid(wt12_actv_pvld[0]),
.io_wt_actv_12_0_bits_nz(wt12_actv_nz[0]),
.io_wt_actv_12_0_bits_data(wt12_actv_data[7:0]),

.io_wt_actv_12_1_valid(wt12_actv_pvld[1]),
.io_wt_actv_12_1_bits_nz(wt12_actv_nz[1]),
.io_wt_actv_12_1_bits_data(wt12_actv_data[15:8]),

.io_wt_actv_12_2_valid(wt12_actv_pvld[2]),
.io_wt_actv_12_2_bits_nz(wt12_actv_nz[2]),
.io_wt_actv_12_2_bits_data(wt12_actv_data[23:16]),

.io_wt_actv_12_3_valid(wt12_actv_pvld[3]),
.io_wt_actv_12_3_bits_nz(wt12_actv_nz[3]),
.io_wt_actv_12_3_bits_data(wt12_actv_data[31:24]),

.io_wt_actv_12_4_valid(wt12_actv_pvld[4]),
.io_wt_actv_12_4_bits_nz(wt12_actv_nz[4]),
.io_wt_actv_12_4_bits_data(wt12_actv_data[39:32]),

.io_wt_actv_12_5_valid(wt12_actv_pvld[5]),
.io_wt_actv_12_5_bits_nz(wt12_actv_nz[5]),
.io_wt_actv_12_5_bits_data(wt12_actv_data[47:40]),

.io_wt_actv_12_6_valid(wt12_actv_pvld[6]),
.io_wt_actv_12_6_bits_nz(wt12_actv_nz[6]),
.io_wt_actv_12_6_bits_data(wt12_actv_data[55:48]),

.io_wt_actv_12_7_valid(wt12_actv_pvld[7]),
.io_wt_actv_12_7_bits_nz(wt12_actv_nz[7]),
.io_wt_actv_12_7_bits_data(wt12_actv_data[63:56]),

.io_wt_actv_12_8_valid(wt12_actv_pvld[8]),
.io_wt_actv_12_8_bits_nz(wt12_actv_nz[8]),
.io_wt_actv_12_8_bits_data(wt12_actv_data[71:64]),

.io_wt_actv_12_9_valid(wt12_actv_pvld[9]),
.io_wt_actv_12_9_bits_nz(wt12_actv_nz[9]),
.io_wt_actv_12_9_bits_data(wt12_actv_data[79:72]),

.io_wt_actv_12_10_valid(wt12_actv_pvld[10]),
.io_wt_actv_12_10_bits_nz(wt12_actv_nz[10]),
.io_wt_actv_12_10_bits_data(wt12_actv_data[87:80]),

.io_wt_actv_12_11_valid(wt12_actv_pvld[11]),
.io_wt_actv_12_11_bits_nz(wt12_actv_nz[11]),
.io_wt_actv_12_11_bits_data(wt12_actv_data[95:88]),

.io_wt_actv_12_12_valid(wt12_actv_pvld[12]),
.io_wt_actv_12_12_bits_nz(wt12_actv_nz[12]),
.io_wt_actv_12_12_bits_data(wt12_actv_data[103:96]),

.io_wt_actv_12_13_valid(wt12_actv_pvld[13]),
.io_wt_actv_12_13_bits_nz(wt12_actv_nz[13]),
.io_wt_actv_12_13_bits_data(wt12_actv_data[111:104]),

.io_wt_actv_12_14_valid(wt12_actv_pvld[14]),
.io_wt_actv_12_14_bits_nz(wt12_actv_nz[14]),
.io_wt_actv_12_14_bits_data(wt12_actv_data[119:112]),

.io_wt_actv_12_15_valid(wt12_actv_pvld[15]),
.io_wt_actv_12_15_bits_nz(wt12_actv_nz[15]),
.io_wt_actv_12_15_bits_data(wt12_actv_data[127:120]),

.io_wt_actv_12_16_valid(wt12_actv_pvld[16]),
.io_wt_actv_12_16_bits_nz(wt12_actv_nz[16]),
.io_wt_actv_12_16_bits_data(wt12_actv_data[135:128]),

.io_wt_actv_12_17_valid(wt12_actv_pvld[17]),
.io_wt_actv_12_17_bits_nz(wt12_actv_nz[17]),
.io_wt_actv_12_17_bits_data(wt12_actv_data[143:136]),

.io_wt_actv_12_18_valid(wt12_actv_pvld[18]),
.io_wt_actv_12_18_bits_nz(wt12_actv_nz[18]),
.io_wt_actv_12_18_bits_data(wt12_actv_data[151:144]),

.io_wt_actv_12_19_valid(wt12_actv_pvld[19]),
.io_wt_actv_12_19_bits_nz(wt12_actv_nz[19]),
.io_wt_actv_12_19_bits_data(wt12_actv_data[159:152]),

.io_wt_actv_12_20_valid(wt12_actv_pvld[20]),
.io_wt_actv_12_20_bits_nz(wt12_actv_nz[20]),
.io_wt_actv_12_20_bits_data(wt12_actv_data[167:160]),

.io_wt_actv_12_21_valid(wt12_actv_pvld[21]),
.io_wt_actv_12_21_bits_nz(wt12_actv_nz[21]),
.io_wt_actv_12_21_bits_data(wt12_actv_data[175:168]),

.io_wt_actv_12_22_valid(wt12_actv_pvld[22]),
.io_wt_actv_12_22_bits_nz(wt12_actv_nz[22]),
.io_wt_actv_12_22_bits_data(wt12_actv_data[183:176]),

.io_wt_actv_12_23_valid(wt12_actv_pvld[23]),
.io_wt_actv_12_23_bits_nz(wt12_actv_nz[23]),
.io_wt_actv_12_23_bits_data(wt12_actv_data[191:184]),

.io_wt_actv_12_24_valid(wt12_actv_pvld[24]),
.io_wt_actv_12_24_bits_nz(wt12_actv_nz[24]),
.io_wt_actv_12_24_bits_data(wt12_actv_data[199:192]),

.io_wt_actv_12_25_valid(wt12_actv_pvld[25]),
.io_wt_actv_12_25_bits_nz(wt12_actv_nz[25]),
.io_wt_actv_12_25_bits_data(wt12_actv_data[207:200]),

.io_wt_actv_12_26_valid(wt12_actv_pvld[26]),
.io_wt_actv_12_26_bits_nz(wt12_actv_nz[26]),
.io_wt_actv_12_26_bits_data(wt12_actv_data[215:208]),

.io_wt_actv_12_27_valid(wt12_actv_pvld[27]),
.io_wt_actv_12_27_bits_nz(wt12_actv_nz[27]),
.io_wt_actv_12_27_bits_data(wt12_actv_data[223:216]),

.io_wt_actv_12_28_valid(wt12_actv_pvld[28]),
.io_wt_actv_12_28_bits_nz(wt12_actv_nz[28]),
.io_wt_actv_12_28_bits_data(wt12_actv_data[231:224]),

.io_wt_actv_12_29_valid(wt12_actv_pvld[29]),
.io_wt_actv_12_29_bits_nz(wt12_actv_nz[29]),
.io_wt_actv_12_29_bits_data(wt12_actv_data[239:232]),

.io_wt_actv_12_30_valid(wt12_actv_pvld[30]),
.io_wt_actv_12_30_bits_nz(wt12_actv_nz[30]),
.io_wt_actv_12_30_bits_data(wt12_actv_data[247:240]),

.io_wt_actv_12_31_valid(wt12_actv_pvld[31]),
.io_wt_actv_12_31_bits_nz(wt12_actv_nz[31]),
.io_wt_actv_12_31_bits_data(wt12_actv_data[255:248]),

.io_wt_actv_12_32_valid(wt12_actv_pvld[32]),
.io_wt_actv_12_32_bits_nz(wt12_actv_nz[32]),
.io_wt_actv_12_32_bits_data(wt12_actv_data[263:256]),

.io_wt_actv_12_33_valid(wt12_actv_pvld[33]),
.io_wt_actv_12_33_bits_nz(wt12_actv_nz[33]),
.io_wt_actv_12_33_bits_data(wt12_actv_data[271:264]),

.io_wt_actv_12_34_valid(wt12_actv_pvld[34]),
.io_wt_actv_12_34_bits_nz(wt12_actv_nz[34]),
.io_wt_actv_12_34_bits_data(wt12_actv_data[279:272]),

.io_wt_actv_12_35_valid(wt12_actv_pvld[35]),
.io_wt_actv_12_35_bits_nz(wt12_actv_nz[35]),
.io_wt_actv_12_35_bits_data(wt12_actv_data[287:280]),

.io_wt_actv_12_36_valid(wt12_actv_pvld[36]),
.io_wt_actv_12_36_bits_nz(wt12_actv_nz[36]),
.io_wt_actv_12_36_bits_data(wt12_actv_data[295:288]),

.io_wt_actv_12_37_valid(wt12_actv_pvld[37]),
.io_wt_actv_12_37_bits_nz(wt12_actv_nz[37]),
.io_wt_actv_12_37_bits_data(wt12_actv_data[303:296]),

.io_wt_actv_12_38_valid(wt12_actv_pvld[38]),
.io_wt_actv_12_38_bits_nz(wt12_actv_nz[38]),
.io_wt_actv_12_38_bits_data(wt12_actv_data[311:304]),

.io_wt_actv_12_39_valid(wt12_actv_pvld[39]),
.io_wt_actv_12_39_bits_nz(wt12_actv_nz[39]),
.io_wt_actv_12_39_bits_data(wt12_actv_data[319:312]),

.io_wt_actv_12_40_valid(wt12_actv_pvld[40]),
.io_wt_actv_12_40_bits_nz(wt12_actv_nz[40]),
.io_wt_actv_12_40_bits_data(wt12_actv_data[327:320]),

.io_wt_actv_12_41_valid(wt12_actv_pvld[41]),
.io_wt_actv_12_41_bits_nz(wt12_actv_nz[41]),
.io_wt_actv_12_41_bits_data(wt12_actv_data[335:328]),

.io_wt_actv_12_42_valid(wt12_actv_pvld[42]),
.io_wt_actv_12_42_bits_nz(wt12_actv_nz[42]),
.io_wt_actv_12_42_bits_data(wt12_actv_data[343:336]),

.io_wt_actv_12_43_valid(wt12_actv_pvld[43]),
.io_wt_actv_12_43_bits_nz(wt12_actv_nz[43]),
.io_wt_actv_12_43_bits_data(wt12_actv_data[351:344]),

.io_wt_actv_12_44_valid(wt12_actv_pvld[44]),
.io_wt_actv_12_44_bits_nz(wt12_actv_nz[44]),
.io_wt_actv_12_44_bits_data(wt12_actv_data[359:352]),

.io_wt_actv_12_45_valid(wt12_actv_pvld[45]),
.io_wt_actv_12_45_bits_nz(wt12_actv_nz[45]),
.io_wt_actv_12_45_bits_data(wt12_actv_data[367:360]),

.io_wt_actv_12_46_valid(wt12_actv_pvld[46]),
.io_wt_actv_12_46_bits_nz(wt12_actv_nz[46]),
.io_wt_actv_12_46_bits_data(wt12_actv_data[375:368]),

.io_wt_actv_12_47_valid(wt12_actv_pvld[47]),
.io_wt_actv_12_47_bits_nz(wt12_actv_nz[47]),
.io_wt_actv_12_47_bits_data(wt12_actv_data[383:376]),

.io_wt_actv_12_48_valid(wt12_actv_pvld[48]),
.io_wt_actv_12_48_bits_nz(wt12_actv_nz[48]),
.io_wt_actv_12_48_bits_data(wt12_actv_data[391:384]),

.io_wt_actv_12_49_valid(wt12_actv_pvld[49]),
.io_wt_actv_12_49_bits_nz(wt12_actv_nz[49]),
.io_wt_actv_12_49_bits_data(wt12_actv_data[399:392]),

.io_wt_actv_12_50_valid(wt12_actv_pvld[50]),
.io_wt_actv_12_50_bits_nz(wt12_actv_nz[50]),
.io_wt_actv_12_50_bits_data(wt12_actv_data[407:400]),

.io_wt_actv_12_51_valid(wt12_actv_pvld[51]),
.io_wt_actv_12_51_bits_nz(wt12_actv_nz[51]),
.io_wt_actv_12_51_bits_data(wt12_actv_data[415:408]),

.io_wt_actv_12_52_valid(wt12_actv_pvld[52]),
.io_wt_actv_12_52_bits_nz(wt12_actv_nz[52]),
.io_wt_actv_12_52_bits_data(wt12_actv_data[423:416]),

.io_wt_actv_12_53_valid(wt12_actv_pvld[53]),
.io_wt_actv_12_53_bits_nz(wt12_actv_nz[53]),
.io_wt_actv_12_53_bits_data(wt12_actv_data[431:424]),

.io_wt_actv_12_54_valid(wt12_actv_pvld[54]),
.io_wt_actv_12_54_bits_nz(wt12_actv_nz[54]),
.io_wt_actv_12_54_bits_data(wt12_actv_data[439:432]),

.io_wt_actv_12_55_valid(wt12_actv_pvld[55]),
.io_wt_actv_12_55_bits_nz(wt12_actv_nz[55]),
.io_wt_actv_12_55_bits_data(wt12_actv_data[447:440]),

.io_wt_actv_12_56_valid(wt12_actv_pvld[56]),
.io_wt_actv_12_56_bits_nz(wt12_actv_nz[56]),
.io_wt_actv_12_56_bits_data(wt12_actv_data[455:448]),

.io_wt_actv_12_57_valid(wt12_actv_pvld[57]),
.io_wt_actv_12_57_bits_nz(wt12_actv_nz[57]),
.io_wt_actv_12_57_bits_data(wt12_actv_data[463:456]),

.io_wt_actv_12_58_valid(wt12_actv_pvld[58]),
.io_wt_actv_12_58_bits_nz(wt12_actv_nz[58]),
.io_wt_actv_12_58_bits_data(wt12_actv_data[471:464]),

.io_wt_actv_12_59_valid(wt12_actv_pvld[59]),
.io_wt_actv_12_59_bits_nz(wt12_actv_nz[59]),
.io_wt_actv_12_59_bits_data(wt12_actv_data[479:472]),

.io_wt_actv_12_60_valid(wt12_actv_pvld[60]),
.io_wt_actv_12_60_bits_nz(wt12_actv_nz[60]),
.io_wt_actv_12_60_bits_data(wt12_actv_data[487:480]),

.io_wt_actv_12_61_valid(wt12_actv_pvld[61]),
.io_wt_actv_12_61_bits_nz(wt12_actv_nz[61]),
.io_wt_actv_12_61_bits_data(wt12_actv_data[495:488]),

.io_wt_actv_12_62_valid(wt12_actv_pvld[62]),
.io_wt_actv_12_62_bits_nz(wt12_actv_nz[62]),
.io_wt_actv_12_62_bits_data(wt12_actv_data[503:496]),

.io_wt_actv_12_63_valid(wt12_actv_pvld[63]),
.io_wt_actv_12_63_bits_nz(wt12_actv_nz[63]),
.io_wt_actv_12_63_bits_data(wt12_actv_data[511:504]),

.io_wt_actv_13_0_valid(wt13_actv_pvld[0]),
.io_wt_actv_13_0_bits_nz(wt13_actv_nz[0]),
.io_wt_actv_13_0_bits_data(wt13_actv_data[7:0]),

.io_wt_actv_13_1_valid(wt13_actv_pvld[1]),
.io_wt_actv_13_1_bits_nz(wt13_actv_nz[1]),
.io_wt_actv_13_1_bits_data(wt13_actv_data[15:8]),

.io_wt_actv_13_2_valid(wt13_actv_pvld[2]),
.io_wt_actv_13_2_bits_nz(wt13_actv_nz[2]),
.io_wt_actv_13_2_bits_data(wt13_actv_data[23:16]),

.io_wt_actv_13_3_valid(wt13_actv_pvld[3]),
.io_wt_actv_13_3_bits_nz(wt13_actv_nz[3]),
.io_wt_actv_13_3_bits_data(wt13_actv_data[31:24]),

.io_wt_actv_13_4_valid(wt13_actv_pvld[4]),
.io_wt_actv_13_4_bits_nz(wt13_actv_nz[4]),
.io_wt_actv_13_4_bits_data(wt13_actv_data[39:32]),

.io_wt_actv_13_5_valid(wt13_actv_pvld[5]),
.io_wt_actv_13_5_bits_nz(wt13_actv_nz[5]),
.io_wt_actv_13_5_bits_data(wt13_actv_data[47:40]),

.io_wt_actv_13_6_valid(wt13_actv_pvld[6]),
.io_wt_actv_13_6_bits_nz(wt13_actv_nz[6]),
.io_wt_actv_13_6_bits_data(wt13_actv_data[55:48]),

.io_wt_actv_13_7_valid(wt13_actv_pvld[7]),
.io_wt_actv_13_7_bits_nz(wt13_actv_nz[7]),
.io_wt_actv_13_7_bits_data(wt13_actv_data[63:56]),

.io_wt_actv_13_8_valid(wt13_actv_pvld[8]),
.io_wt_actv_13_8_bits_nz(wt13_actv_nz[8]),
.io_wt_actv_13_8_bits_data(wt13_actv_data[71:64]),

.io_wt_actv_13_9_valid(wt13_actv_pvld[9]),
.io_wt_actv_13_9_bits_nz(wt13_actv_nz[9]),
.io_wt_actv_13_9_bits_data(wt13_actv_data[79:72]),

.io_wt_actv_13_10_valid(wt13_actv_pvld[10]),
.io_wt_actv_13_10_bits_nz(wt13_actv_nz[10]),
.io_wt_actv_13_10_bits_data(wt13_actv_data[87:80]),

.io_wt_actv_13_11_valid(wt13_actv_pvld[11]),
.io_wt_actv_13_11_bits_nz(wt13_actv_nz[11]),
.io_wt_actv_13_11_bits_data(wt13_actv_data[95:88]),

.io_wt_actv_13_12_valid(wt13_actv_pvld[12]),
.io_wt_actv_13_12_bits_nz(wt13_actv_nz[12]),
.io_wt_actv_13_12_bits_data(wt13_actv_data[103:96]),

.io_wt_actv_13_13_valid(wt13_actv_pvld[13]),
.io_wt_actv_13_13_bits_nz(wt13_actv_nz[13]),
.io_wt_actv_13_13_bits_data(wt13_actv_data[111:104]),

.io_wt_actv_13_14_valid(wt13_actv_pvld[14]),
.io_wt_actv_13_14_bits_nz(wt13_actv_nz[14]),
.io_wt_actv_13_14_bits_data(wt13_actv_data[119:112]),

.io_wt_actv_13_15_valid(wt13_actv_pvld[15]),
.io_wt_actv_13_15_bits_nz(wt13_actv_nz[15]),
.io_wt_actv_13_15_bits_data(wt13_actv_data[127:120]),

.io_wt_actv_13_16_valid(wt13_actv_pvld[16]),
.io_wt_actv_13_16_bits_nz(wt13_actv_nz[16]),
.io_wt_actv_13_16_bits_data(wt13_actv_data[135:128]),

.io_wt_actv_13_17_valid(wt13_actv_pvld[17]),
.io_wt_actv_13_17_bits_nz(wt13_actv_nz[17]),
.io_wt_actv_13_17_bits_data(wt13_actv_data[143:136]),

.io_wt_actv_13_18_valid(wt13_actv_pvld[18]),
.io_wt_actv_13_18_bits_nz(wt13_actv_nz[18]),
.io_wt_actv_13_18_bits_data(wt13_actv_data[151:144]),

.io_wt_actv_13_19_valid(wt13_actv_pvld[19]),
.io_wt_actv_13_19_bits_nz(wt13_actv_nz[19]),
.io_wt_actv_13_19_bits_data(wt13_actv_data[159:152]),

.io_wt_actv_13_20_valid(wt13_actv_pvld[20]),
.io_wt_actv_13_20_bits_nz(wt13_actv_nz[20]),
.io_wt_actv_13_20_bits_data(wt13_actv_data[167:160]),

.io_wt_actv_13_21_valid(wt13_actv_pvld[21]),
.io_wt_actv_13_21_bits_nz(wt13_actv_nz[21]),
.io_wt_actv_13_21_bits_data(wt13_actv_data[175:168]),

.io_wt_actv_13_22_valid(wt13_actv_pvld[22]),
.io_wt_actv_13_22_bits_nz(wt13_actv_nz[22]),
.io_wt_actv_13_22_bits_data(wt13_actv_data[183:176]),

.io_wt_actv_13_23_valid(wt13_actv_pvld[23]),
.io_wt_actv_13_23_bits_nz(wt13_actv_nz[23]),
.io_wt_actv_13_23_bits_data(wt13_actv_data[191:184]),

.io_wt_actv_13_24_valid(wt13_actv_pvld[24]),
.io_wt_actv_13_24_bits_nz(wt13_actv_nz[24]),
.io_wt_actv_13_24_bits_data(wt13_actv_data[199:192]),

.io_wt_actv_13_25_valid(wt13_actv_pvld[25]),
.io_wt_actv_13_25_bits_nz(wt13_actv_nz[25]),
.io_wt_actv_13_25_bits_data(wt13_actv_data[207:200]),

.io_wt_actv_13_26_valid(wt13_actv_pvld[26]),
.io_wt_actv_13_26_bits_nz(wt13_actv_nz[26]),
.io_wt_actv_13_26_bits_data(wt13_actv_data[215:208]),

.io_wt_actv_13_27_valid(wt13_actv_pvld[27]),
.io_wt_actv_13_27_bits_nz(wt13_actv_nz[27]),
.io_wt_actv_13_27_bits_data(wt13_actv_data[223:216]),

.io_wt_actv_13_28_valid(wt13_actv_pvld[28]),
.io_wt_actv_13_28_bits_nz(wt13_actv_nz[28]),
.io_wt_actv_13_28_bits_data(wt13_actv_data[231:224]),

.io_wt_actv_13_29_valid(wt13_actv_pvld[29]),
.io_wt_actv_13_29_bits_nz(wt13_actv_nz[29]),
.io_wt_actv_13_29_bits_data(wt13_actv_data[239:232]),

.io_wt_actv_13_30_valid(wt13_actv_pvld[30]),
.io_wt_actv_13_30_bits_nz(wt13_actv_nz[30]),
.io_wt_actv_13_30_bits_data(wt13_actv_data[247:240]),

.io_wt_actv_13_31_valid(wt13_actv_pvld[31]),
.io_wt_actv_13_31_bits_nz(wt13_actv_nz[31]),
.io_wt_actv_13_31_bits_data(wt13_actv_data[255:248]),

.io_wt_actv_13_32_valid(wt13_actv_pvld[32]),
.io_wt_actv_13_32_bits_nz(wt13_actv_nz[32]),
.io_wt_actv_13_32_bits_data(wt13_actv_data[263:256]),

.io_wt_actv_13_33_valid(wt13_actv_pvld[33]),
.io_wt_actv_13_33_bits_nz(wt13_actv_nz[33]),
.io_wt_actv_13_33_bits_data(wt13_actv_data[271:264]),

.io_wt_actv_13_34_valid(wt13_actv_pvld[34]),
.io_wt_actv_13_34_bits_nz(wt13_actv_nz[34]),
.io_wt_actv_13_34_bits_data(wt13_actv_data[279:272]),

.io_wt_actv_13_35_valid(wt13_actv_pvld[35]),
.io_wt_actv_13_35_bits_nz(wt13_actv_nz[35]),
.io_wt_actv_13_35_bits_data(wt13_actv_data[287:280]),

.io_wt_actv_13_36_valid(wt13_actv_pvld[36]),
.io_wt_actv_13_36_bits_nz(wt13_actv_nz[36]),
.io_wt_actv_13_36_bits_data(wt13_actv_data[295:288]),

.io_wt_actv_13_37_valid(wt13_actv_pvld[37]),
.io_wt_actv_13_37_bits_nz(wt13_actv_nz[37]),
.io_wt_actv_13_37_bits_data(wt13_actv_data[303:296]),

.io_wt_actv_13_38_valid(wt13_actv_pvld[38]),
.io_wt_actv_13_38_bits_nz(wt13_actv_nz[38]),
.io_wt_actv_13_38_bits_data(wt13_actv_data[311:304]),

.io_wt_actv_13_39_valid(wt13_actv_pvld[39]),
.io_wt_actv_13_39_bits_nz(wt13_actv_nz[39]),
.io_wt_actv_13_39_bits_data(wt13_actv_data[319:312]),

.io_wt_actv_13_40_valid(wt13_actv_pvld[40]),
.io_wt_actv_13_40_bits_nz(wt13_actv_nz[40]),
.io_wt_actv_13_40_bits_data(wt13_actv_data[327:320]),

.io_wt_actv_13_41_valid(wt13_actv_pvld[41]),
.io_wt_actv_13_41_bits_nz(wt13_actv_nz[41]),
.io_wt_actv_13_41_bits_data(wt13_actv_data[335:328]),

.io_wt_actv_13_42_valid(wt13_actv_pvld[42]),
.io_wt_actv_13_42_bits_nz(wt13_actv_nz[42]),
.io_wt_actv_13_42_bits_data(wt13_actv_data[343:336]),

.io_wt_actv_13_43_valid(wt13_actv_pvld[43]),
.io_wt_actv_13_43_bits_nz(wt13_actv_nz[43]),
.io_wt_actv_13_43_bits_data(wt13_actv_data[351:344]),

.io_wt_actv_13_44_valid(wt13_actv_pvld[44]),
.io_wt_actv_13_44_bits_nz(wt13_actv_nz[44]),
.io_wt_actv_13_44_bits_data(wt13_actv_data[359:352]),

.io_wt_actv_13_45_valid(wt13_actv_pvld[45]),
.io_wt_actv_13_45_bits_nz(wt13_actv_nz[45]),
.io_wt_actv_13_45_bits_data(wt13_actv_data[367:360]),

.io_wt_actv_13_46_valid(wt13_actv_pvld[46]),
.io_wt_actv_13_46_bits_nz(wt13_actv_nz[46]),
.io_wt_actv_13_46_bits_data(wt13_actv_data[375:368]),

.io_wt_actv_13_47_valid(wt13_actv_pvld[47]),
.io_wt_actv_13_47_bits_nz(wt13_actv_nz[47]),
.io_wt_actv_13_47_bits_data(wt13_actv_data[383:376]),

.io_wt_actv_13_48_valid(wt13_actv_pvld[48]),
.io_wt_actv_13_48_bits_nz(wt13_actv_nz[48]),
.io_wt_actv_13_48_bits_data(wt13_actv_data[391:384]),

.io_wt_actv_13_49_valid(wt13_actv_pvld[49]),
.io_wt_actv_13_49_bits_nz(wt13_actv_nz[49]),
.io_wt_actv_13_49_bits_data(wt13_actv_data[399:392]),

.io_wt_actv_13_50_valid(wt13_actv_pvld[50]),
.io_wt_actv_13_50_bits_nz(wt13_actv_nz[50]),
.io_wt_actv_13_50_bits_data(wt13_actv_data[407:400]),

.io_wt_actv_13_51_valid(wt13_actv_pvld[51]),
.io_wt_actv_13_51_bits_nz(wt13_actv_nz[51]),
.io_wt_actv_13_51_bits_data(wt13_actv_data[415:408]),

.io_wt_actv_13_52_valid(wt13_actv_pvld[52]),
.io_wt_actv_13_52_bits_nz(wt13_actv_nz[52]),
.io_wt_actv_13_52_bits_data(wt13_actv_data[423:416]),

.io_wt_actv_13_53_valid(wt13_actv_pvld[53]),
.io_wt_actv_13_53_bits_nz(wt13_actv_nz[53]),
.io_wt_actv_13_53_bits_data(wt13_actv_data[431:424]),

.io_wt_actv_13_54_valid(wt13_actv_pvld[54]),
.io_wt_actv_13_54_bits_nz(wt13_actv_nz[54]),
.io_wt_actv_13_54_bits_data(wt13_actv_data[439:432]),

.io_wt_actv_13_55_valid(wt13_actv_pvld[55]),
.io_wt_actv_13_55_bits_nz(wt13_actv_nz[55]),
.io_wt_actv_13_55_bits_data(wt13_actv_data[447:440]),

.io_wt_actv_13_56_valid(wt13_actv_pvld[56]),
.io_wt_actv_13_56_bits_nz(wt13_actv_nz[56]),
.io_wt_actv_13_56_bits_data(wt13_actv_data[455:448]),

.io_wt_actv_13_57_valid(wt13_actv_pvld[57]),
.io_wt_actv_13_57_bits_nz(wt13_actv_nz[57]),
.io_wt_actv_13_57_bits_data(wt13_actv_data[463:456]),

.io_wt_actv_13_58_valid(wt13_actv_pvld[58]),
.io_wt_actv_13_58_bits_nz(wt13_actv_nz[58]),
.io_wt_actv_13_58_bits_data(wt13_actv_data[471:464]),

.io_wt_actv_13_59_valid(wt13_actv_pvld[59]),
.io_wt_actv_13_59_bits_nz(wt13_actv_nz[59]),
.io_wt_actv_13_59_bits_data(wt13_actv_data[479:472]),

.io_wt_actv_13_60_valid(wt13_actv_pvld[60]),
.io_wt_actv_13_60_bits_nz(wt13_actv_nz[60]),
.io_wt_actv_13_60_bits_data(wt13_actv_data[487:480]),

.io_wt_actv_13_61_valid(wt13_actv_pvld[61]),
.io_wt_actv_13_61_bits_nz(wt13_actv_nz[61]),
.io_wt_actv_13_61_bits_data(wt13_actv_data[495:488]),

.io_wt_actv_13_62_valid(wt13_actv_pvld[62]),
.io_wt_actv_13_62_bits_nz(wt13_actv_nz[62]),
.io_wt_actv_13_62_bits_data(wt13_actv_data[503:496]),

.io_wt_actv_13_63_valid(wt13_actv_pvld[63]),
.io_wt_actv_13_63_bits_nz(wt13_actv_nz[63]),
.io_wt_actv_13_63_bits_data(wt13_actv_data[511:504]),

.io_wt_actv_14_0_valid(wt14_actv_pvld[0]),
.io_wt_actv_14_0_bits_nz(wt14_actv_nz[0]),
.io_wt_actv_14_0_bits_data(wt14_actv_data[7:0]),

.io_wt_actv_14_1_valid(wt14_actv_pvld[1]),
.io_wt_actv_14_1_bits_nz(wt14_actv_nz[1]),
.io_wt_actv_14_1_bits_data(wt14_actv_data[15:8]),

.io_wt_actv_14_2_valid(wt14_actv_pvld[2]),
.io_wt_actv_14_2_bits_nz(wt14_actv_nz[2]),
.io_wt_actv_14_2_bits_data(wt14_actv_data[23:16]),

.io_wt_actv_14_3_valid(wt14_actv_pvld[3]),
.io_wt_actv_14_3_bits_nz(wt14_actv_nz[3]),
.io_wt_actv_14_3_bits_data(wt14_actv_data[31:24]),

.io_wt_actv_14_4_valid(wt14_actv_pvld[4]),
.io_wt_actv_14_4_bits_nz(wt14_actv_nz[4]),
.io_wt_actv_14_4_bits_data(wt14_actv_data[39:32]),

.io_wt_actv_14_5_valid(wt14_actv_pvld[5]),
.io_wt_actv_14_5_bits_nz(wt14_actv_nz[5]),
.io_wt_actv_14_5_bits_data(wt14_actv_data[47:40]),

.io_wt_actv_14_6_valid(wt14_actv_pvld[6]),
.io_wt_actv_14_6_bits_nz(wt14_actv_nz[6]),
.io_wt_actv_14_6_bits_data(wt14_actv_data[55:48]),

.io_wt_actv_14_7_valid(wt14_actv_pvld[7]),
.io_wt_actv_14_7_bits_nz(wt14_actv_nz[7]),
.io_wt_actv_14_7_bits_data(wt14_actv_data[63:56]),

.io_wt_actv_14_8_valid(wt14_actv_pvld[8]),
.io_wt_actv_14_8_bits_nz(wt14_actv_nz[8]),
.io_wt_actv_14_8_bits_data(wt14_actv_data[71:64]),

.io_wt_actv_14_9_valid(wt14_actv_pvld[9]),
.io_wt_actv_14_9_bits_nz(wt14_actv_nz[9]),
.io_wt_actv_14_9_bits_data(wt14_actv_data[79:72]),

.io_wt_actv_14_10_valid(wt14_actv_pvld[10]),
.io_wt_actv_14_10_bits_nz(wt14_actv_nz[10]),
.io_wt_actv_14_10_bits_data(wt14_actv_data[87:80]),

.io_wt_actv_14_11_valid(wt14_actv_pvld[11]),
.io_wt_actv_14_11_bits_nz(wt14_actv_nz[11]),
.io_wt_actv_14_11_bits_data(wt14_actv_data[95:88]),

.io_wt_actv_14_12_valid(wt14_actv_pvld[12]),
.io_wt_actv_14_12_bits_nz(wt14_actv_nz[12]),
.io_wt_actv_14_12_bits_data(wt14_actv_data[103:96]),

.io_wt_actv_14_13_valid(wt14_actv_pvld[13]),
.io_wt_actv_14_13_bits_nz(wt14_actv_nz[13]),
.io_wt_actv_14_13_bits_data(wt14_actv_data[111:104]),

.io_wt_actv_14_14_valid(wt14_actv_pvld[14]),
.io_wt_actv_14_14_bits_nz(wt14_actv_nz[14]),
.io_wt_actv_14_14_bits_data(wt14_actv_data[119:112]),

.io_wt_actv_14_15_valid(wt14_actv_pvld[15]),
.io_wt_actv_14_15_bits_nz(wt14_actv_nz[15]),
.io_wt_actv_14_15_bits_data(wt14_actv_data[127:120]),

.io_wt_actv_14_16_valid(wt14_actv_pvld[16]),
.io_wt_actv_14_16_bits_nz(wt14_actv_nz[16]),
.io_wt_actv_14_16_bits_data(wt14_actv_data[135:128]),

.io_wt_actv_14_17_valid(wt14_actv_pvld[17]),
.io_wt_actv_14_17_bits_nz(wt14_actv_nz[17]),
.io_wt_actv_14_17_bits_data(wt14_actv_data[143:136]),

.io_wt_actv_14_18_valid(wt14_actv_pvld[18]),
.io_wt_actv_14_18_bits_nz(wt14_actv_nz[18]),
.io_wt_actv_14_18_bits_data(wt14_actv_data[151:144]),

.io_wt_actv_14_19_valid(wt14_actv_pvld[19]),
.io_wt_actv_14_19_bits_nz(wt14_actv_nz[19]),
.io_wt_actv_14_19_bits_data(wt14_actv_data[159:152]),

.io_wt_actv_14_20_valid(wt14_actv_pvld[20]),
.io_wt_actv_14_20_bits_nz(wt14_actv_nz[20]),
.io_wt_actv_14_20_bits_data(wt14_actv_data[167:160]),

.io_wt_actv_14_21_valid(wt14_actv_pvld[21]),
.io_wt_actv_14_21_bits_nz(wt14_actv_nz[21]),
.io_wt_actv_14_21_bits_data(wt14_actv_data[175:168]),

.io_wt_actv_14_22_valid(wt14_actv_pvld[22]),
.io_wt_actv_14_22_bits_nz(wt14_actv_nz[22]),
.io_wt_actv_14_22_bits_data(wt14_actv_data[183:176]),

.io_wt_actv_14_23_valid(wt14_actv_pvld[23]),
.io_wt_actv_14_23_bits_nz(wt14_actv_nz[23]),
.io_wt_actv_14_23_bits_data(wt14_actv_data[191:184]),

.io_wt_actv_14_24_valid(wt14_actv_pvld[24]),
.io_wt_actv_14_24_bits_nz(wt14_actv_nz[24]),
.io_wt_actv_14_24_bits_data(wt14_actv_data[199:192]),

.io_wt_actv_14_25_valid(wt14_actv_pvld[25]),
.io_wt_actv_14_25_bits_nz(wt14_actv_nz[25]),
.io_wt_actv_14_25_bits_data(wt14_actv_data[207:200]),

.io_wt_actv_14_26_valid(wt14_actv_pvld[26]),
.io_wt_actv_14_26_bits_nz(wt14_actv_nz[26]),
.io_wt_actv_14_26_bits_data(wt14_actv_data[215:208]),

.io_wt_actv_14_27_valid(wt14_actv_pvld[27]),
.io_wt_actv_14_27_bits_nz(wt14_actv_nz[27]),
.io_wt_actv_14_27_bits_data(wt14_actv_data[223:216]),

.io_wt_actv_14_28_valid(wt14_actv_pvld[28]),
.io_wt_actv_14_28_bits_nz(wt14_actv_nz[28]),
.io_wt_actv_14_28_bits_data(wt14_actv_data[231:224]),

.io_wt_actv_14_29_valid(wt14_actv_pvld[29]),
.io_wt_actv_14_29_bits_nz(wt14_actv_nz[29]),
.io_wt_actv_14_29_bits_data(wt14_actv_data[239:232]),

.io_wt_actv_14_30_valid(wt14_actv_pvld[30]),
.io_wt_actv_14_30_bits_nz(wt14_actv_nz[30]),
.io_wt_actv_14_30_bits_data(wt14_actv_data[247:240]),

.io_wt_actv_14_31_valid(wt14_actv_pvld[31]),
.io_wt_actv_14_31_bits_nz(wt14_actv_nz[31]),
.io_wt_actv_14_31_bits_data(wt14_actv_data[255:248]),

.io_wt_actv_14_32_valid(wt14_actv_pvld[32]),
.io_wt_actv_14_32_bits_nz(wt14_actv_nz[32]),
.io_wt_actv_14_32_bits_data(wt14_actv_data[263:256]),

.io_wt_actv_14_33_valid(wt14_actv_pvld[33]),
.io_wt_actv_14_33_bits_nz(wt14_actv_nz[33]),
.io_wt_actv_14_33_bits_data(wt14_actv_data[271:264]),

.io_wt_actv_14_34_valid(wt14_actv_pvld[34]),
.io_wt_actv_14_34_bits_nz(wt14_actv_nz[34]),
.io_wt_actv_14_34_bits_data(wt14_actv_data[279:272]),

.io_wt_actv_14_35_valid(wt14_actv_pvld[35]),
.io_wt_actv_14_35_bits_nz(wt14_actv_nz[35]),
.io_wt_actv_14_35_bits_data(wt14_actv_data[287:280]),

.io_wt_actv_14_36_valid(wt14_actv_pvld[36]),
.io_wt_actv_14_36_bits_nz(wt14_actv_nz[36]),
.io_wt_actv_14_36_bits_data(wt14_actv_data[295:288]),

.io_wt_actv_14_37_valid(wt14_actv_pvld[37]),
.io_wt_actv_14_37_bits_nz(wt14_actv_nz[37]),
.io_wt_actv_14_37_bits_data(wt14_actv_data[303:296]),

.io_wt_actv_14_38_valid(wt14_actv_pvld[38]),
.io_wt_actv_14_38_bits_nz(wt14_actv_nz[38]),
.io_wt_actv_14_38_bits_data(wt14_actv_data[311:304]),

.io_wt_actv_14_39_valid(wt14_actv_pvld[39]),
.io_wt_actv_14_39_bits_nz(wt14_actv_nz[39]),
.io_wt_actv_14_39_bits_data(wt14_actv_data[319:312]),

.io_wt_actv_14_40_valid(wt14_actv_pvld[40]),
.io_wt_actv_14_40_bits_nz(wt14_actv_nz[40]),
.io_wt_actv_14_40_bits_data(wt14_actv_data[327:320]),

.io_wt_actv_14_41_valid(wt14_actv_pvld[41]),
.io_wt_actv_14_41_bits_nz(wt14_actv_nz[41]),
.io_wt_actv_14_41_bits_data(wt14_actv_data[335:328]),

.io_wt_actv_14_42_valid(wt14_actv_pvld[42]),
.io_wt_actv_14_42_bits_nz(wt14_actv_nz[42]),
.io_wt_actv_14_42_bits_data(wt14_actv_data[343:336]),

.io_wt_actv_14_43_valid(wt14_actv_pvld[43]),
.io_wt_actv_14_43_bits_nz(wt14_actv_nz[43]),
.io_wt_actv_14_43_bits_data(wt14_actv_data[351:344]),

.io_wt_actv_14_44_valid(wt14_actv_pvld[44]),
.io_wt_actv_14_44_bits_nz(wt14_actv_nz[44]),
.io_wt_actv_14_44_bits_data(wt14_actv_data[359:352]),

.io_wt_actv_14_45_valid(wt14_actv_pvld[45]),
.io_wt_actv_14_45_bits_nz(wt14_actv_nz[45]),
.io_wt_actv_14_45_bits_data(wt14_actv_data[367:360]),

.io_wt_actv_14_46_valid(wt14_actv_pvld[46]),
.io_wt_actv_14_46_bits_nz(wt14_actv_nz[46]),
.io_wt_actv_14_46_bits_data(wt14_actv_data[375:368]),

.io_wt_actv_14_47_valid(wt14_actv_pvld[47]),
.io_wt_actv_14_47_bits_nz(wt14_actv_nz[47]),
.io_wt_actv_14_47_bits_data(wt14_actv_data[383:376]),

.io_wt_actv_14_48_valid(wt14_actv_pvld[48]),
.io_wt_actv_14_48_bits_nz(wt14_actv_nz[48]),
.io_wt_actv_14_48_bits_data(wt14_actv_data[391:384]),

.io_wt_actv_14_49_valid(wt14_actv_pvld[49]),
.io_wt_actv_14_49_bits_nz(wt14_actv_nz[49]),
.io_wt_actv_14_49_bits_data(wt14_actv_data[399:392]),

.io_wt_actv_14_50_valid(wt14_actv_pvld[50]),
.io_wt_actv_14_50_bits_nz(wt14_actv_nz[50]),
.io_wt_actv_14_50_bits_data(wt14_actv_data[407:400]),

.io_wt_actv_14_51_valid(wt14_actv_pvld[51]),
.io_wt_actv_14_51_bits_nz(wt14_actv_nz[51]),
.io_wt_actv_14_51_bits_data(wt14_actv_data[415:408]),

.io_wt_actv_14_52_valid(wt14_actv_pvld[52]),
.io_wt_actv_14_52_bits_nz(wt14_actv_nz[52]),
.io_wt_actv_14_52_bits_data(wt14_actv_data[423:416]),

.io_wt_actv_14_53_valid(wt14_actv_pvld[53]),
.io_wt_actv_14_53_bits_nz(wt14_actv_nz[53]),
.io_wt_actv_14_53_bits_data(wt14_actv_data[431:424]),

.io_wt_actv_14_54_valid(wt14_actv_pvld[54]),
.io_wt_actv_14_54_bits_nz(wt14_actv_nz[54]),
.io_wt_actv_14_54_bits_data(wt14_actv_data[439:432]),

.io_wt_actv_14_55_valid(wt14_actv_pvld[55]),
.io_wt_actv_14_55_bits_nz(wt14_actv_nz[55]),
.io_wt_actv_14_55_bits_data(wt14_actv_data[447:440]),

.io_wt_actv_14_56_valid(wt14_actv_pvld[56]),
.io_wt_actv_14_56_bits_nz(wt14_actv_nz[56]),
.io_wt_actv_14_56_bits_data(wt14_actv_data[455:448]),

.io_wt_actv_14_57_valid(wt14_actv_pvld[57]),
.io_wt_actv_14_57_bits_nz(wt14_actv_nz[57]),
.io_wt_actv_14_57_bits_data(wt14_actv_data[463:456]),

.io_wt_actv_14_58_valid(wt14_actv_pvld[58]),
.io_wt_actv_14_58_bits_nz(wt14_actv_nz[58]),
.io_wt_actv_14_58_bits_data(wt14_actv_data[471:464]),

.io_wt_actv_14_59_valid(wt14_actv_pvld[59]),
.io_wt_actv_14_59_bits_nz(wt14_actv_nz[59]),
.io_wt_actv_14_59_bits_data(wt14_actv_data[479:472]),

.io_wt_actv_14_60_valid(wt14_actv_pvld[60]),
.io_wt_actv_14_60_bits_nz(wt14_actv_nz[60]),
.io_wt_actv_14_60_bits_data(wt14_actv_data[487:480]),

.io_wt_actv_14_61_valid(wt14_actv_pvld[61]),
.io_wt_actv_14_61_bits_nz(wt14_actv_nz[61]),
.io_wt_actv_14_61_bits_data(wt14_actv_data[495:488]),

.io_wt_actv_14_62_valid(wt14_actv_pvld[62]),
.io_wt_actv_14_62_bits_nz(wt14_actv_nz[62]),
.io_wt_actv_14_62_bits_data(wt14_actv_data[503:496]),

.io_wt_actv_14_63_valid(wt14_actv_pvld[63]),
.io_wt_actv_14_63_bits_nz(wt14_actv_nz[63]),
.io_wt_actv_14_63_bits_data(wt14_actv_data[511:504]),

.io_wt_actv_15_0_valid(wt15_actv_pvld[0]),
.io_wt_actv_15_0_bits_nz(wt15_actv_nz[0]),
.io_wt_actv_15_0_bits_data(wt15_actv_data[7:0]),

.io_wt_actv_15_1_valid(wt15_actv_pvld[1]),
.io_wt_actv_15_1_bits_nz(wt15_actv_nz[1]),
.io_wt_actv_15_1_bits_data(wt15_actv_data[15:8]),

.io_wt_actv_15_2_valid(wt15_actv_pvld[2]),
.io_wt_actv_15_2_bits_nz(wt15_actv_nz[2]),
.io_wt_actv_15_2_bits_data(wt15_actv_data[23:16]),

.io_wt_actv_15_3_valid(wt15_actv_pvld[3]),
.io_wt_actv_15_3_bits_nz(wt15_actv_nz[3]),
.io_wt_actv_15_3_bits_data(wt15_actv_data[31:24]),

.io_wt_actv_15_4_valid(wt15_actv_pvld[4]),
.io_wt_actv_15_4_bits_nz(wt15_actv_nz[4]),
.io_wt_actv_15_4_bits_data(wt15_actv_data[39:32]),

.io_wt_actv_15_5_valid(wt15_actv_pvld[5]),
.io_wt_actv_15_5_bits_nz(wt15_actv_nz[5]),
.io_wt_actv_15_5_bits_data(wt15_actv_data[47:40]),

.io_wt_actv_15_6_valid(wt15_actv_pvld[6]),
.io_wt_actv_15_6_bits_nz(wt15_actv_nz[6]),
.io_wt_actv_15_6_bits_data(wt15_actv_data[55:48]),

.io_wt_actv_15_7_valid(wt15_actv_pvld[7]),
.io_wt_actv_15_7_bits_nz(wt15_actv_nz[7]),
.io_wt_actv_15_7_bits_data(wt15_actv_data[63:56]),

.io_wt_actv_15_8_valid(wt15_actv_pvld[8]),
.io_wt_actv_15_8_bits_nz(wt15_actv_nz[8]),
.io_wt_actv_15_8_bits_data(wt15_actv_data[71:64]),

.io_wt_actv_15_9_valid(wt15_actv_pvld[9]),
.io_wt_actv_15_9_bits_nz(wt15_actv_nz[9]),
.io_wt_actv_15_9_bits_data(wt15_actv_data[79:72]),

.io_wt_actv_15_10_valid(wt15_actv_pvld[10]),
.io_wt_actv_15_10_bits_nz(wt15_actv_nz[10]),
.io_wt_actv_15_10_bits_data(wt15_actv_data[87:80]),

.io_wt_actv_15_11_valid(wt15_actv_pvld[11]),
.io_wt_actv_15_11_bits_nz(wt15_actv_nz[11]),
.io_wt_actv_15_11_bits_data(wt15_actv_data[95:88]),

.io_wt_actv_15_12_valid(wt15_actv_pvld[12]),
.io_wt_actv_15_12_bits_nz(wt15_actv_nz[12]),
.io_wt_actv_15_12_bits_data(wt15_actv_data[103:96]),

.io_wt_actv_15_13_valid(wt15_actv_pvld[13]),
.io_wt_actv_15_13_bits_nz(wt15_actv_nz[13]),
.io_wt_actv_15_13_bits_data(wt15_actv_data[111:104]),

.io_wt_actv_15_14_valid(wt15_actv_pvld[14]),
.io_wt_actv_15_14_bits_nz(wt15_actv_nz[14]),
.io_wt_actv_15_14_bits_data(wt15_actv_data[119:112]),

.io_wt_actv_15_15_valid(wt15_actv_pvld[15]),
.io_wt_actv_15_15_bits_nz(wt15_actv_nz[15]),
.io_wt_actv_15_15_bits_data(wt15_actv_data[127:120]),

.io_wt_actv_15_16_valid(wt15_actv_pvld[16]),
.io_wt_actv_15_16_bits_nz(wt15_actv_nz[16]),
.io_wt_actv_15_16_bits_data(wt15_actv_data[135:128]),

.io_wt_actv_15_17_valid(wt15_actv_pvld[17]),
.io_wt_actv_15_17_bits_nz(wt15_actv_nz[17]),
.io_wt_actv_15_17_bits_data(wt15_actv_data[143:136]),

.io_wt_actv_15_18_valid(wt15_actv_pvld[18]),
.io_wt_actv_15_18_bits_nz(wt15_actv_nz[18]),
.io_wt_actv_15_18_bits_data(wt15_actv_data[151:144]),

.io_wt_actv_15_19_valid(wt15_actv_pvld[19]),
.io_wt_actv_15_19_bits_nz(wt15_actv_nz[19]),
.io_wt_actv_15_19_bits_data(wt15_actv_data[159:152]),

.io_wt_actv_15_20_valid(wt15_actv_pvld[20]),
.io_wt_actv_15_20_bits_nz(wt15_actv_nz[20]),
.io_wt_actv_15_20_bits_data(wt15_actv_data[167:160]),

.io_wt_actv_15_21_valid(wt15_actv_pvld[21]),
.io_wt_actv_15_21_bits_nz(wt15_actv_nz[21]),
.io_wt_actv_15_21_bits_data(wt15_actv_data[175:168]),

.io_wt_actv_15_22_valid(wt15_actv_pvld[22]),
.io_wt_actv_15_22_bits_nz(wt15_actv_nz[22]),
.io_wt_actv_15_22_bits_data(wt15_actv_data[183:176]),

.io_wt_actv_15_23_valid(wt15_actv_pvld[23]),
.io_wt_actv_15_23_bits_nz(wt15_actv_nz[23]),
.io_wt_actv_15_23_bits_data(wt15_actv_data[191:184]),

.io_wt_actv_15_24_valid(wt15_actv_pvld[24]),
.io_wt_actv_15_24_bits_nz(wt15_actv_nz[24]),
.io_wt_actv_15_24_bits_data(wt15_actv_data[199:192]),

.io_wt_actv_15_25_valid(wt15_actv_pvld[25]),
.io_wt_actv_15_25_bits_nz(wt15_actv_nz[25]),
.io_wt_actv_15_25_bits_data(wt15_actv_data[207:200]),

.io_wt_actv_15_26_valid(wt15_actv_pvld[26]),
.io_wt_actv_15_26_bits_nz(wt15_actv_nz[26]),
.io_wt_actv_15_26_bits_data(wt15_actv_data[215:208]),

.io_wt_actv_15_27_valid(wt15_actv_pvld[27]),
.io_wt_actv_15_27_bits_nz(wt15_actv_nz[27]),
.io_wt_actv_15_27_bits_data(wt15_actv_data[223:216]),

.io_wt_actv_15_28_valid(wt15_actv_pvld[28]),
.io_wt_actv_15_28_bits_nz(wt15_actv_nz[28]),
.io_wt_actv_15_28_bits_data(wt15_actv_data[231:224]),

.io_wt_actv_15_29_valid(wt15_actv_pvld[29]),
.io_wt_actv_15_29_bits_nz(wt15_actv_nz[29]),
.io_wt_actv_15_29_bits_data(wt15_actv_data[239:232]),

.io_wt_actv_15_30_valid(wt15_actv_pvld[30]),
.io_wt_actv_15_30_bits_nz(wt15_actv_nz[30]),
.io_wt_actv_15_30_bits_data(wt15_actv_data[247:240]),

.io_wt_actv_15_31_valid(wt15_actv_pvld[31]),
.io_wt_actv_15_31_bits_nz(wt15_actv_nz[31]),
.io_wt_actv_15_31_bits_data(wt15_actv_data[255:248]),

.io_wt_actv_15_32_valid(wt15_actv_pvld[32]),
.io_wt_actv_15_32_bits_nz(wt15_actv_nz[32]),
.io_wt_actv_15_32_bits_data(wt15_actv_data[263:256]),

.io_wt_actv_15_33_valid(wt15_actv_pvld[33]),
.io_wt_actv_15_33_bits_nz(wt15_actv_nz[33]),
.io_wt_actv_15_33_bits_data(wt15_actv_data[271:264]),

.io_wt_actv_15_34_valid(wt15_actv_pvld[34]),
.io_wt_actv_15_34_bits_nz(wt15_actv_nz[34]),
.io_wt_actv_15_34_bits_data(wt15_actv_data[279:272]),

.io_wt_actv_15_35_valid(wt15_actv_pvld[35]),
.io_wt_actv_15_35_bits_nz(wt15_actv_nz[35]),
.io_wt_actv_15_35_bits_data(wt15_actv_data[287:280]),

.io_wt_actv_15_36_valid(wt15_actv_pvld[36]),
.io_wt_actv_15_36_bits_nz(wt15_actv_nz[36]),
.io_wt_actv_15_36_bits_data(wt15_actv_data[295:288]),

.io_wt_actv_15_37_valid(wt15_actv_pvld[37]),
.io_wt_actv_15_37_bits_nz(wt15_actv_nz[37]),
.io_wt_actv_15_37_bits_data(wt15_actv_data[303:296]),

.io_wt_actv_15_38_valid(wt15_actv_pvld[38]),
.io_wt_actv_15_38_bits_nz(wt15_actv_nz[38]),
.io_wt_actv_15_38_bits_data(wt15_actv_data[311:304]),

.io_wt_actv_15_39_valid(wt15_actv_pvld[39]),
.io_wt_actv_15_39_bits_nz(wt15_actv_nz[39]),
.io_wt_actv_15_39_bits_data(wt15_actv_data[319:312]),

.io_wt_actv_15_40_valid(wt15_actv_pvld[40]),
.io_wt_actv_15_40_bits_nz(wt15_actv_nz[40]),
.io_wt_actv_15_40_bits_data(wt15_actv_data[327:320]),

.io_wt_actv_15_41_valid(wt15_actv_pvld[41]),
.io_wt_actv_15_41_bits_nz(wt15_actv_nz[41]),
.io_wt_actv_15_41_bits_data(wt15_actv_data[335:328]),

.io_wt_actv_15_42_valid(wt15_actv_pvld[42]),
.io_wt_actv_15_42_bits_nz(wt15_actv_nz[42]),
.io_wt_actv_15_42_bits_data(wt15_actv_data[343:336]),

.io_wt_actv_15_43_valid(wt15_actv_pvld[43]),
.io_wt_actv_15_43_bits_nz(wt15_actv_nz[43]),
.io_wt_actv_15_43_bits_data(wt15_actv_data[351:344]),

.io_wt_actv_15_44_valid(wt15_actv_pvld[44]),
.io_wt_actv_15_44_bits_nz(wt15_actv_nz[44]),
.io_wt_actv_15_44_bits_data(wt15_actv_data[359:352]),

.io_wt_actv_15_45_valid(wt15_actv_pvld[45]),
.io_wt_actv_15_45_bits_nz(wt15_actv_nz[45]),
.io_wt_actv_15_45_bits_data(wt15_actv_data[367:360]),

.io_wt_actv_15_46_valid(wt15_actv_pvld[46]),
.io_wt_actv_15_46_bits_nz(wt15_actv_nz[46]),
.io_wt_actv_15_46_bits_data(wt15_actv_data[375:368]),

.io_wt_actv_15_47_valid(wt15_actv_pvld[47]),
.io_wt_actv_15_47_bits_nz(wt15_actv_nz[47]),
.io_wt_actv_15_47_bits_data(wt15_actv_data[383:376]),

.io_wt_actv_15_48_valid(wt15_actv_pvld[48]),
.io_wt_actv_15_48_bits_nz(wt15_actv_nz[48]),
.io_wt_actv_15_48_bits_data(wt15_actv_data[391:384]),

.io_wt_actv_15_49_valid(wt15_actv_pvld[49]),
.io_wt_actv_15_49_bits_nz(wt15_actv_nz[49]),
.io_wt_actv_15_49_bits_data(wt15_actv_data[399:392]),

.io_wt_actv_15_50_valid(wt15_actv_pvld[50]),
.io_wt_actv_15_50_bits_nz(wt15_actv_nz[50]),
.io_wt_actv_15_50_bits_data(wt15_actv_data[407:400]),

.io_wt_actv_15_51_valid(wt15_actv_pvld[51]),
.io_wt_actv_15_51_bits_nz(wt15_actv_nz[51]),
.io_wt_actv_15_51_bits_data(wt15_actv_data[415:408]),

.io_wt_actv_15_52_valid(wt15_actv_pvld[52]),
.io_wt_actv_15_52_bits_nz(wt15_actv_nz[52]),
.io_wt_actv_15_52_bits_data(wt15_actv_data[423:416]),

.io_wt_actv_15_53_valid(wt15_actv_pvld[53]),
.io_wt_actv_15_53_bits_nz(wt15_actv_nz[53]),
.io_wt_actv_15_53_bits_data(wt15_actv_data[431:424]),

.io_wt_actv_15_54_valid(wt15_actv_pvld[54]),
.io_wt_actv_15_54_bits_nz(wt15_actv_nz[54]),
.io_wt_actv_15_54_bits_data(wt15_actv_data[439:432]),

.io_wt_actv_15_55_valid(wt15_actv_pvld[55]),
.io_wt_actv_15_55_bits_nz(wt15_actv_nz[55]),
.io_wt_actv_15_55_bits_data(wt15_actv_data[447:440]),

.io_wt_actv_15_56_valid(wt15_actv_pvld[56]),
.io_wt_actv_15_56_bits_nz(wt15_actv_nz[56]),
.io_wt_actv_15_56_bits_data(wt15_actv_data[455:448]),

.io_wt_actv_15_57_valid(wt15_actv_pvld[57]),
.io_wt_actv_15_57_bits_nz(wt15_actv_nz[57]),
.io_wt_actv_15_57_bits_data(wt15_actv_data[463:456]),

.io_wt_actv_15_58_valid(wt15_actv_pvld[58]),
.io_wt_actv_15_58_bits_nz(wt15_actv_nz[58]),
.io_wt_actv_15_58_bits_data(wt15_actv_data[471:464]),

.io_wt_actv_15_59_valid(wt15_actv_pvld[59]),
.io_wt_actv_15_59_bits_nz(wt15_actv_nz[59]),
.io_wt_actv_15_59_bits_data(wt15_actv_data[479:472]),

.io_wt_actv_15_60_valid(wt15_actv_pvld[60]),
.io_wt_actv_15_60_bits_nz(wt15_actv_nz[60]),
.io_wt_actv_15_60_bits_data(wt15_actv_data[487:480]),

.io_wt_actv_15_61_valid(wt15_actv_pvld[61]),
.io_wt_actv_15_61_bits_nz(wt15_actv_nz[61]),
.io_wt_actv_15_61_bits_data(wt15_actv_data[495:488]),

.io_wt_actv_15_62_valid(wt15_actv_pvld[62]),
.io_wt_actv_15_62_bits_nz(wt15_actv_nz[62]),
.io_wt_actv_15_62_bits_data(wt15_actv_data[503:496]),

.io_wt_actv_15_63_valid(wt15_actv_pvld[63]),
.io_wt_actv_15_63_bits_nz(wt15_actv_nz[63]),
.io_wt_actv_15_63_bits_data(wt15_actv_data[511:504])

);
endmodule
