module NV_soDLA_CSC_dl( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input          io_nvdla_core_clk, // @[:@6.4]
  input          io_nvdla_core_ng_clk, // @[:@6.4]
  input  [1:0]   io_sc_state, // @[:@6.4]
  input          io_sg2dl_pd_valid, // @[:@6.4]
  input  [30:0]  io_sg2dl_pd_bits, // @[:@6.4]
  input          io_sg2dl_reuse_rls, // @[:@6.4]
  input          io_cdma2sc_dat_updt_valid, // @[:@6.4]
  input  [14:0]  io_cdma2sc_dat_updt_bits_entries, // @[:@6.4]
  input  [13:0]  io_cdma2sc_dat_updt_bits_slices, // @[:@6.4]
  input          io_sc2cdma_dat_pending_req, // @[:@6.4]
  output         io_sc2cdma_dat_updt_valid, // @[:@6.4]
  output [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@6.4]
  output [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@6.4]
  output         io_sc2buf_dat_rd_addr_valid, // @[:@6.4]
  output [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@6.4]
  input          io_sc2buf_dat_rd_data_valid, // @[:@6.4]
  input  [511:0] io_sc2buf_dat_rd_data_bits, // @[:@6.4]
  output         io_sc2mac_dat_a_valid, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_0, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_1, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_2, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_3, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_4, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_5, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_6, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_7, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_8, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_9, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_10, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_11, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_12, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_13, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_14, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_15, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_16, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_17, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_18, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_19, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_20, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_21, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_22, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_23, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_24, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_25, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_26, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_27, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_28, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_29, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_30, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_31, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_32, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_33, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_34, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_35, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_36, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_37, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_38, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_39, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_40, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_41, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_42, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_43, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_44, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_45, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_46, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_47, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_48, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_49, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_50, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_51, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_52, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_53, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_54, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_55, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_56, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_57, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_58, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_59, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_60, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_61, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_62, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_63, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_a_bits_pd, // @[:@6.4]
  output         io_sc2mac_dat_b_valid, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_0, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_1, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_2, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_3, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_4, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_5, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_6, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_7, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_8, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_9, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_10, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_11, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_12, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_13, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_14, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_15, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_16, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_17, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_18, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_19, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_20, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_21, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_22, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_23, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_24, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_25, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_26, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_27, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_28, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_29, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_30, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_31, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_32, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_33, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_34, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_35, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_36, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_37, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_38, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_39, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_40, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_41, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_42, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_43, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_44, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_45, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_46, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_47, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_48, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_49, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_50, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_51, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_52, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_53, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_54, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_55, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_56, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_57, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_58, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_59, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_60, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_61, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_62, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_63, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_b_bits_pd, // @[:@6.4]
  input          io_reg2dp_op_en, // @[:@6.4]
  input          io_reg2dp_conv_mode, // @[:@6.4]
  input  [4:0]   io_reg2dp_batches, // @[:@6.4]
  input  [1:0]   io_reg2dp_proc_precision, // @[:@6.4]
  input          io_reg2dp_datain_format, // @[:@6.4]
  input          io_reg2dp_skip_data_rls, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_channel_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_height_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_width_ext, // @[:@6.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@6.4]
  input  [12:0]  io_reg2dp_weight_channel_ext, // @[:@6.4]
  input  [13:0]  io_reg2dp_entries, // @[:@6.4]
  input  [12:0]  io_reg2dp_dataout_width, // @[:@6.4]
  input  [11:0]  io_reg2dp_rls_slices, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_x_stride_ext, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_y_stride_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_x_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_y_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_top, // @[:@6.4]
  input  [15:0]  io_reg2dp_pad_value, // @[:@6.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@6.4]
  input  [1:0]   io_reg2dp_pra_truncate, // @[:@6.4]
  output         io_slcg_wg_en // @[:@6.4]
);
  wire  _T_622; // @[NV_NVDLA_CSC_dl.scala 75:31:@8.4]
  wire  _T_626; // @[NV_NVDLA_CSC_dl.scala 77:31:@10.4]
  wire  _T_630; // @[NV_NVDLA_CSC_dl.scala 84:32:@13.4]
  wire  _T_634; // @[NV_NVDLA_CSC_dl.scala 86:35:@15.4]
  wire  _T_635; // @[NV_NVDLA_CSC_dl.scala 87:22:@16.4]
  wire [6:0] _T_640; // @[NV_NVDLA_CSC_dl.scala 94:53:@17.4]
  wire [6:0] _T_642; // @[NV_NVDLA_CSC_dl.scala 94:24:@18.4]
  wire [2:0] _T_643; // @[NV_NVDLA_CSC_dl.scala 94:100:@19.4]
  wire [2:0] _T_645; // @[NV_NVDLA_CSC_dl.scala 95:22:@20.4]
  wire [3:0] _T_647; // @[NV_NVDLA_CSC_dl.scala 96:34:@21.4]
  wire [3:0] _T_648; // @[NV_NVDLA_CSC_dl.scala 96:34:@22.4]
  wire [3:0] _T_650; // @[NV_NVDLA_CSC_dl.scala 97:51:@23.4]
  wire [1:0] _T_651; // @[NV_NVDLA_CSC_dl.scala 98:62:@24.4]
  wire [5:0] _T_654; // @[Cat.scala 30:58:@25.4]
  wire [4:0] _T_657; // @[Cat.scala 30:58:@26.4]
  wire [4:0] _GEN_671; // @[NV_NVDLA_CSC_dl.scala 100:74:@27.4]
  wire [5:0] _T_658; // @[NV_NVDLA_CSC_dl.scala 100:74:@27.4]
  wire  _T_659; // @[Mux.scala 46:19:@28.4]
  wire [5:0] _T_660; // @[Mux.scala 46:16:@29.4]
  wire  _T_661; // @[Mux.scala 46:19:@30.4]
  wire [5:0] _T_662; // @[Mux.scala 46:16:@31.4]
  wire  _T_664; // @[NV_NVDLA_CSC_dl.scala 102:88:@32.4]
  wire [5:0] _T_670; // @[NV_NVDLA_CSC_dl.scala 102:172:@34.4]
  wire [5:0] _T_671; // @[NV_NVDLA_CSC_dl.scala 102:58:@35.4]
  wire [6:0] _T_674; // @[Cat.scala 30:58:@36.4]
  wire [6:0] _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@37.4]
  wire [7:0] _T_675; // @[NV_NVDLA_CSC_dl.scala 103:81:@37.4]
  wire [6:0] _T_676; // @[NV_NVDLA_CSC_dl.scala 103:81:@38.4]
  wire [6:0] _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@40.4]
  wire [7:0] _T_678; // @[NV_NVDLA_CSC_dl.scala 103:100:@40.4]
  wire [6:0] _T_679; // @[NV_NVDLA_CSC_dl.scala 103:100:@41.4]
  wire [6:0] _T_682; // @[NV_NVDLA_CSC_dl.scala 104:58:@43.4]
  wire [5:0] _T_683; // @[NV_NVDLA_CSC_dl.scala 104:58:@44.4]
  wire  _T_684; // @[Mux.scala 46:19:@45.4]
  wire [5:0] _T_685; // @[Mux.scala 46:16:@46.4]
  wire  _T_686; // @[Mux.scala 46:19:@47.4]
  wire [6:0] _T_687; // @[Mux.scala 46:16:@48.4]
  wire [6:0] _T_690; // @[NV_NVDLA_CSC_dl.scala 105:80:@50.4]
  wire [7:0] _T_693; // @[Cat.scala 30:58:@51.4]
  wire [6:0] _T_698; // @[Mux.scala 46:16:@54.4]
  wire [7:0] _T_700; // @[Mux.scala 46:16:@56.4]
  wire [11:0] _T_702; // @[Cat.scala 30:58:@57.4]
  wire [3:0] _T_704; // @[NV_NVDLA_CSC_dl.scala 115:52:@58.4]
  wire [5:0] _T_707; // @[NV_NVDLA_CSC_dl.scala 116:60:@59.4]
  wire [5:0] _T_708; // @[NV_NVDLA_CSC_dl.scala 116:21:@60.4]
  wire [5:0] _T_711; // @[NV_NVDLA_CSC_dl.scala 117:60:@61.4]
  wire [5:0] _T_712; // @[NV_NVDLA_CSC_dl.scala 117:21:@62.4]
  reg  _T_715; // @[NV_NVDLA_CSC_dl.scala 119:26:@63.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_722; // @[NV_NVDLA_CSC_dl.scala 120:25:@65.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_729; // @[NV_NVDLA_CSC_dl.scala 121:25:@67.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_736; // @[NV_NVDLA_CSC_dl.scala 122:29:@69.4]
  reg [31:0] _RAND_3;
  reg [14:0] _T_743; // @[NV_NVDLA_CSC_dl.scala 123:22:@71.4]
  reg [31:0] _RAND_4;
  reg [14:0] _T_750; // @[NV_NVDLA_CSC_dl.scala 124:28:@73.4]
  reg [31:0] _RAND_5;
  reg [12:0] _T_757; // @[NV_NVDLA_CSC_dl.scala 125:32:@75.4]
  reg [31:0] _RAND_6;
  reg [14:0] _T_771; // @[NV_NVDLA_CSC_dl.scala 127:26:@79.4]
  reg [31:0] _RAND_7;
  reg [11:0] _T_778; // @[NV_NVDLA_CSC_dl.scala 128:30:@81.4]
  reg [31:0] _RAND_8;
  reg [11:0] _T_785; // @[NV_NVDLA_CSC_dl.scala 129:30:@83.4]
  reg [31:0] _RAND_9;
  reg [13:0] _T_792; // @[NV_NVDLA_CSC_dl.scala 130:25:@85.4]
  reg [31:0] _RAND_10;
  wire [14:0] _T_794; // @[NV_NVDLA_CSC_dl.scala 133:43:@86.4]
  wire [20:0] _T_796; // @[NV_NVDLA_CSC_dl.scala 134:41:@88.4]
  wire [14:0] _T_797; // @[NV_NVDLA_CSC_dl.scala 134:56:@89.4]
  wire [11:0] _T_798; // @[NV_NVDLA_CSC_dl.scala 136:37:@90.4]
  wire [14:0] _GEN_674; // @[NV_NVDLA_CSC_dl.scala 137:34:@91.4]
  wire [20:0] _T_799; // @[NV_NVDLA_CSC_dl.scala 137:34:@91.4]
  wire [11:0] _T_800; // @[NV_NVDLA_CSC_dl.scala 137:47:@92.4]
  wire [14:0] _GEN_675; // @[NV_NVDLA_CSC_dl.scala 138:34:@93.4]
  wire [28:0] _T_801; // @[NV_NVDLA_CSC_dl.scala 138:34:@93.4]
  wire [11:0] _T_802; // @[NV_NVDLA_CSC_dl.scala 138:51:@94.4]
  wire [12:0] _T_804; // @[NV_NVDLA_CSC_dl.scala 139:41:@95.4]
  wire [11:0] _T_805; // @[NV_NVDLA_CSC_dl.scala 139:41:@96.4]
  wire [13:0] _T_807; // @[NV_NVDLA_CSC_dl.scala 140:77:@97.4]
  wire [12:0] _GEN_676; // @[NV_NVDLA_CSC_dl.scala 140:113:@98.4]
  wire [13:0] _T_808; // @[NV_NVDLA_CSC_dl.scala 140:113:@98.4]
  wire [13:0] _T_809; // @[NV_NVDLA_CSC_dl.scala 140:113:@99.4]
  wire [13:0] _T_810; // @[NV_NVDLA_CSC_dl.scala 140:23:@100.4]
  wire [13:0] _T_811; // @[NV_NVDLA_CSC_dl.scala 141:24:@101.4]
  wire [14:0] _GEN_677; // @[NV_NVDLA_CSC_dl.scala 142:38:@102.4]
  wire [28:0] _T_812; // @[NV_NVDLA_CSC_dl.scala 142:38:@102.4]
  wire [14:0] _T_813; // @[NV_NVDLA_CSC_dl.scala 142:54:@103.4]
  reg [33:0] _T_831; // @[NV_NVDLA_CSC_dl.scala 147:24:@109.4]
  reg [63:0] _RAND_11;
  reg [4:0] _T_838; // @[NV_NVDLA_CSC_dl.scala 148:24:@111.4]
  reg [31:0] _RAND_12;
  reg [13:0] _T_845; // @[NV_NVDLA_CSC_dl.scala 149:27:@113.4]
  reg [31:0] _RAND_13;
  reg [12:0] _T_852; // @[NV_NVDLA_CSC_dl.scala 150:31:@115.4]
  reg [31:0] _RAND_14;
  reg [12:0] _T_859; // @[NV_NVDLA_CSC_dl.scala 151:32:@117.4]
  reg [31:0] _RAND_15;
  reg [10:0] _T_866; // @[NV_NVDLA_CSC_dl.scala 152:33:@119.4]
  reg [31:0] _RAND_16;
  reg [2:0] _T_869; // @[NV_NVDLA_CSC_dl.scala 153:29:@120.4]
  reg [31:0] _RAND_17;
  reg [2:0] _T_872; // @[NV_NVDLA_CSC_dl.scala 154:29:@121.4]
  reg [31:0] _RAND_18;
  reg [2:0] _T_878; // @[NV_NVDLA_CSC_dl.scala 156:29:@123.4]
  reg [31:0] _RAND_19;
  reg [2:0] _T_881; // @[NV_NVDLA_CSC_dl.scala 157:29:@124.4]
  reg [31:0] _RAND_20;
  reg [2:0] _T_884; // @[NV_NVDLA_CSC_dl.scala 158:29:@125.4]
  reg [31:0] _RAND_21;
  reg [2:0] _T_887; // @[NV_NVDLA_CSC_dl.scala 159:29:@126.4]
  reg [31:0] _RAND_22;
  reg [2:0] _T_893; // @[NV_NVDLA_CSC_dl.scala 161:29:@128.4]
  reg [31:0] _RAND_23;
  reg [2:0] _T_896; // @[NV_NVDLA_CSC_dl.scala 162:29:@129.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_902; // @[NV_NVDLA_CSC_dl.scala 164:30:@131.4]
  reg [31:0] _RAND_25;
  reg [2:0] _T_905; // @[NV_NVDLA_CSC_dl.scala 165:27:@132.4]
  reg [31:0] _RAND_26;
  reg [2:0] _T_908; // @[NV_NVDLA_CSC_dl.scala 166:27:@133.4]
  reg [31:0] _RAND_27;
  reg [3:0] _T_915; // @[NV_NVDLA_CSC_dl.scala 167:28:@135.4]
  reg [31:0] _RAND_28;
  reg [3:0] _T_922; // @[NV_NVDLA_CSC_dl.scala 168:28:@137.4]
  reg [31:0] _RAND_29;
  reg [4:0] _T_932; // @[NV_NVDLA_CSC_dl.scala 170:24:@140.4]
  reg [31:0] _RAND_30;
  reg [6:0] _T_939; // @[NV_NVDLA_CSC_dl.scala 171:27:@142.4]
  reg [31:0] _RAND_31;
  reg [6:0] _T_946; // @[NV_NVDLA_CSC_dl.scala 172:34:@144.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_953; // @[NV_NVDLA_CSC_dl.scala 173:26:@146.4]
  reg [31:0] _RAND_33;
  reg [6:0] _T_960; // @[NV_NVDLA_CSC_dl.scala 174:34:@148.4]
  reg [31:0] _RAND_34;
  reg [11:0] _T_967; // @[NV_NVDLA_CSC_dl.scala 175:30:@150.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_974; // @[NV_NVDLA_CSC_dl.scala 176:23:@152.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_981; // @[NV_NVDLA_CSC_dl.scala 177:23:@154.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_988; // @[NV_NVDLA_CSC_dl.scala 178:24:@156.4]
  reg [31:0] _RAND_38;
  reg [14:0] _T_995; // @[NV_NVDLA_CSC_dl.scala 179:26:@158.4]
  reg [31:0] _RAND_39;
  reg [14:0] _T_1002; // @[NV_NVDLA_CSC_dl.scala 180:30:@160.4]
  reg [31:0] _RAND_40;
  reg [14:0] _T_1009; // @[NV_NVDLA_CSC_dl.scala 181:30:@162.4]
  reg [31:0] _RAND_41;
  reg [13:0] _T_1016; // @[NV_NVDLA_CSC_dl.scala 183:26:@164.4]
  reg [31:0] _RAND_42;
  reg [14:0] _T_1023; // @[NV_NVDLA_CSC_dl.scala 184:27:@166.4]
  reg [31:0] _RAND_43;
  wire [33:0] _T_1038; // @[Bitwise.scala 72:12:@174.6]
  wire [5:0] _T_1040; // @[NV_NVDLA_CSC_dl.scala 191:38:@176.6]
  wire [4:0] _T_1041; // @[NV_NVDLA_CSC_dl.scala 191:38:@177.6]
  wire [13:0] _T_1043; // @[NV_NVDLA_CSC_dl.scala 192:48:@179.6]
  wire [6:0] _T_1049; // @[NV_NVDLA_CSC_dl.scala 195:93:@184.6]
  wire [10:0] _T_1050; // @[Cat.scala 30:58:@185.6]
  wire [14:0] _T_1054; // @[Cat.scala 30:58:@218.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [4:0] _GEN_2; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  wire [11:0] _GEN_43; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  wire [11:0] _GEN_44; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  wire [14:0] _GEN_46; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  wire [14:0] _GEN_47; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl.scala 240:17:@238.4]
  wire [14:0] _GEN_49; // @[NV_NVDLA_CSC_dl.scala 240:17:@238.4]
  reg [14:0] _T_1076; // @[NV_NVDLA_CSC_dl.scala 263:59:@250.4]
  reg [31:0] _RAND_44;
  wire  _T_1156; // @[NV_NVDLA_CSC_dl.scala 304:37:@313.4]
  wire  _T_1157; // @[NV_NVDLA_CSC_dl.scala 304:23:@314.4]
  wire  _T_2241; // @[NV_NVDLA_CSC_dl.scala 894:32:@1228.4]
  reg  _T_2217; // @[NV_NVDLA_CSC_dl.scala 879:41:@1196.4]
  reg [31:0] _RAND_45;
  wire  _T_2242; // @[NV_NVDLA_CSC_dl.scala 894:36:@1229.4]
  wire  _T_2243; // @[NV_NVDLA_CSC_dl.scala 895:35:@1230.4]
  reg  _T_2211; // @[NV_NVDLA_CSC_dl.scala 879:41:@1194.4]
  reg [31:0] _RAND_46;
  wire  _T_2244; // @[NV_NVDLA_CSC_dl.scala 895:39:@1231.4]
  wire  _T_2245; // @[NV_NVDLA_CSC_dl.scala 894:57:@1232.4]
  wire  _T_2246; // @[NV_NVDLA_CSC_dl.scala 896:35:@1233.4]
  reg  _T_2208; // @[NV_NVDLA_CSC_dl.scala 879:41:@1193.4]
  reg [31:0] _RAND_47;
  wire  _T_2247; // @[NV_NVDLA_CSC_dl.scala 896:39:@1234.4]
  wire  _T_2248; // @[NV_NVDLA_CSC_dl.scala 895:60:@1235.4]
  wire  _T_2249; // @[NV_NVDLA_CSC_dl.scala 903:42:@1237.4]
  wire [26:0] _T_2253; // @[Bitwise.scala 72:12:@1239.4]
  reg [26:0] _T_2231; // @[NV_NVDLA_CSC_dl.scala 881:41:@1201.4]
  reg [31:0] _RAND_48;
  wire [26:0] _T_2254; // @[NV_NVDLA_CSC_dl.scala 903:47:@1240.4]
  wire  _T_2255; // @[NV_NVDLA_CSC_dl.scala 904:42:@1241.4]
  wire [26:0] _T_2259; // @[Bitwise.scala 72:12:@1243.4]
  reg [26:0] _T_2225; // @[NV_NVDLA_CSC_dl.scala 881:41:@1199.4]
  reg [31:0] _RAND_49;
  wire [26:0] _T_2260; // @[NV_NVDLA_CSC_dl.scala 904:47:@1244.4]
  wire [26:0] _T_2261; // @[NV_NVDLA_CSC_dl.scala 903:66:@1245.4]
  wire  _T_2262; // @[NV_NVDLA_CSC_dl.scala 905:42:@1246.4]
  wire [26:0] _T_2266; // @[Bitwise.scala 72:12:@1248.4]
  reg [26:0] _T_2222; // @[NV_NVDLA_CSC_dl.scala 881:41:@1198.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_2267; // @[NV_NVDLA_CSC_dl.scala 905:47:@1249.4]
  wire [26:0] _T_2268; // @[NV_NVDLA_CSC_dl.scala 904:66:@1250.4]
  wire  _T_2287; // @[NV_NVDLA_CSC_dl.scala 929:26:@1269.4]
  wire  _T_1154; // @[NV_NVDLA_CSC_dl.scala 301:29:@312.4]
  wire  _T_1159; // @[NV_NVDLA_CSC_dl.scala 304:66:@315.4]
  wire  _T_1160; // @[NV_NVDLA_CSC_dl.scala 304:53:@316.4]
  wire  _T_1161; // @[NV_NVDLA_CSC_dl.scala 304:42:@317.4]
  wire [13:0] _T_1162; // @[NV_NVDLA_CSC_dl.scala 305:28:@319.4]
  wire [14:0] _T_1163; // @[NV_NVDLA_CSC_dl.scala 306:29:@321.4]
  wire [14:0] _T_1094; // @[NV_NVDLA_CSC_dl.scala 273:28:@261.4]
  wire [15:0] _T_1102; // @[NV_NVDLA_CSC_dl.scala 278:37:@268.4]
  wire [14:0] _T_1103; // @[NV_NVDLA_CSC_dl.scala 278:37:@269.4]
  wire [13:0] _T_1109; // @[Cat.scala 30:58:@271.4]
  wire [14:0] _GEN_678; // @[NV_NVDLA_CSC_dl.scala 279:46:@272.4]
  wire [15:0] _T_1110; // @[NV_NVDLA_CSC_dl.scala 279:46:@272.4]
  wire [15:0] _T_1111; // @[NV_NVDLA_CSC_dl.scala 279:46:@273.4]
  wire [14:0] _T_1112; // @[NV_NVDLA_CSC_dl.scala 279:46:@274.4]
  wire  _T_1119; // @[NV_NVDLA_CSC_dl.scala 280:45:@277.4]
  wire [14:0] _T_1121; // @[NV_NVDLA_CSC_dl.scala 281:83:@278.4]
  wire [14:0] _T_1122; // @[NV_NVDLA_CSC_dl.scala 281:25:@279.4]
  wire  _T_1148; // @[NV_NVDLA_CSC_dl.scala 292:13:@302.4]
  wire [14:0] _GEN_52; // @[NV_NVDLA_CSC_dl.scala 292:25:@303.4]
  reg  _T_1166; // @[NV_NVDLA_CSC_dl.scala 308:37:@323.4]
  reg [31:0] _RAND_51;
  reg [13:0] _T_1169; // @[Reg.scala 19:20:@326.4]
  reg [31:0] _RAND_52;
  wire [13:0] _GEN_54; // @[Reg.scala 20:19:@327.4]
  reg [14:0] _T_1172; // @[Reg.scala 19:20:@331.4]
  reg [31:0] _RAND_53;
  wire [14:0] _GEN_55; // @[Reg.scala 20:19:@332.4]
  reg  _T_1177; // @[NV_NVDLA_CSC_dl.scala 321:50:@337.4]
  reg [31:0] _RAND_54;
  reg  _T_1180; // @[NV_NVDLA_CSC_dl.scala 321:50:@338.4]
  reg [31:0] _RAND_55;
  reg  _T_1183; // @[NV_NVDLA_CSC_dl.scala 321:50:@339.4]
  reg [31:0] _RAND_56;
  reg  _T_1186; // @[NV_NVDLA_CSC_dl.scala 321:50:@340.4]
  reg [31:0] _RAND_57;
  reg  _T_1189; // @[NV_NVDLA_CSC_dl.scala 321:50:@341.4]
  reg [31:0] _RAND_58;
  reg  _T_1211; // @[NV_NVDLA_CSC_dl.scala 340:36:@371.4]
  reg [31:0] _RAND_59;
  reg  _T_1214; // @[NV_NVDLA_CSC_dl.scala 340:36:@372.4]
  reg [31:0] _RAND_60;
  reg  _T_1217; // @[NV_NVDLA_CSC_dl.scala 340:36:@373.4]
  reg [31:0] _RAND_61;
  reg  _T_1220; // @[NV_NVDLA_CSC_dl.scala 340:36:@374.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_1225; // @[NV_NVDLA_CSC_dl.scala 342:34:@376.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_1228; // @[NV_NVDLA_CSC_dl.scala 342:34:@377.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_1231; // @[NV_NVDLA_CSC_dl.scala 342:34:@378.4]
  reg [31:0] _RAND_65;
  reg [30:0] _T_1234; // @[NV_NVDLA_CSC_dl.scala 342:34:@379.4]
  reg [31:0] _RAND_66;
  wire [30:0] _T_1222; // @[NV_NVDLA_CSC_dl.scala 341:19:@375.4 NV_NVDLA_CSC_dl.scala 345:12:@381.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl.scala 349:23:@383.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl.scala 349:23:@387.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl.scala 349:23:@391.4]
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl.scala 349:23:@395.4]
  wire  _T_1235; // @[NV_NVDLA_CSC_dl.scala 354:30:@398.4]
  wire  _T_1236; // @[NV_NVDLA_CSC_dl.scala 354:34:@399.4]
  wire  _T_1237; // @[NV_NVDLA_CSC_dl.scala 355:30:@400.4]
  wire  _T_1238; // @[NV_NVDLA_CSC_dl.scala 355:34:@401.4]
  wire  _T_1239; // @[NV_NVDLA_CSC_dl.scala 354:50:@402.4]
  wire  _T_1240; // @[NV_NVDLA_CSC_dl.scala 356:30:@403.4]
  wire  _T_1241; // @[NV_NVDLA_CSC_dl.scala 356:34:@404.4]
  wire  _T_1242; // @[NV_NVDLA_CSC_dl.scala 355:50:@405.4]
  wire  _T_1243; // @[NV_NVDLA_CSC_dl.scala 358:37:@406.4]
  wire [30:0] _T_1247; // @[Bitwise.scala 72:12:@408.4]
  wire [30:0] _T_1248; // @[NV_NVDLA_CSC_dl.scala 358:42:@409.4]
  wire  _T_1249; // @[NV_NVDLA_CSC_dl.scala 359:37:@410.4]
  wire [30:0] _T_1253; // @[Bitwise.scala 72:12:@412.4]
  wire [30:0] _T_1254; // @[NV_NVDLA_CSC_dl.scala 359:42:@413.4]
  wire [30:0] _T_1255; // @[NV_NVDLA_CSC_dl.scala 358:56:@414.4]
  wire  _T_1256; // @[NV_NVDLA_CSC_dl.scala 360:37:@415.4]
  wire [30:0] _T_1260; // @[Bitwise.scala 72:12:@417.4]
  wire [30:0] _T_1261; // @[NV_NVDLA_CSC_dl.scala 360:42:@418.4]
  wire [30:0] _T_1262; // @[NV_NVDLA_CSC_dl.scala 359:56:@419.4]
  wire [4:0] _T_1263; // @[NV_NVDLA_CSC_dl.scala 363:24:@420.4]
  wire [4:0] _T_1264; // @[NV_NVDLA_CSC_dl.scala 364:24:@421.4]
  wire [6:0] _T_1265; // @[NV_NVDLA_CSC_dl.scala 365:28:@422.4]
  wire [6:0] _T_1266; // @[NV_NVDLA_CSC_dl.scala 366:29:@423.4]
  wire [1:0] _T_1267; // @[NV_NVDLA_CSC_dl.scala 367:25:@424.4]
  wire  _T_1268; // @[NV_NVDLA_CSC_dl.scala 368:25:@425.4]
  wire  _T_1269; // @[NV_NVDLA_CSC_dl.scala 369:27:@426.4]
  wire  _T_1270; // @[NV_NVDLA_CSC_dl.scala 370:25:@427.4]
  wire  _T_1271; // @[NV_NVDLA_CSC_dl.scala 371:25:@428.4]
  wire  _T_1272; // @[NV_NVDLA_CSC_dl.scala 372:27:@429.4]
  reg [4:0] _T_1279; // @[NV_NVDLA_CSC_dl.scala 377:24:@432.4]
  reg [31:0] _RAND_67;
  wire [5:0] _T_1283; // @[NV_NVDLA_CSC_dl.scala 381:24:@433.4]
  wire [4:0] _T_1284; // @[NV_NVDLA_CSC_dl.scala 381:24:@434.4]
  wire  _T_1287; // @[NV_NVDLA_CSC_dl.scala 383:27:@438.4]
  wire [4:0] _T_1285; // @[NV_NVDLA_CSC_dl.scala 380:17:@435.4]
  wire [4:0] _T_1286; // @[NV_NVDLA_CSC_dl.scala 379:17:@436.4]
  reg [1:0] _T_1290; // @[NV_NVDLA_CSC_dl.scala 386:24:@440.4]
  reg [31:0] _RAND_68;
  wire [2:0] _T_1294; // @[NV_NVDLA_CSC_dl.scala 389:31:@442.4]
  wire [1:0] _T_1295; // @[NV_NVDLA_CSC_dl.scala 389:31:@443.4]
  wire [2:0] _GEN_682; // @[NV_NVDLA_CSC_dl.scala 390:32:@444.4]
  wire  _T_1296; // @[NV_NVDLA_CSC_dl.scala 390:32:@444.4]
  wire  _T_1298; // @[NV_NVDLA_CSC_dl.scala 391:61:@446.4]
  reg [6:0] _T_1306; // @[NV_NVDLA_CSC_dl.scala 397:25:@454.4]
  reg [31:0] _RAND_69;
  wire  _T_1346; // @[NV_NVDLA_CSC_dl.scala 424:37:@483.4]
  wire  _T_1347; // @[NV_NVDLA_CSC_dl.scala 424:24:@484.4]
  wire  _T_1349; // @[NV_NVDLA_CSC_dl.scala 424:56:@485.4]
  wire  _T_1350; // @[NV_NVDLA_CSC_dl.scala 424:44:@486.4]
  wire  _T_1351; // @[NV_NVDLA_CSC_dl.scala 424:42:@487.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_dl.scala 424:75:@488.4]
  wire  _T_1354; // @[NV_NVDLA_CSC_dl.scala 424:63:@489.4]
  wire  _T_1355; // @[NV_NVDLA_CSC_dl.scala 424:61:@490.4]
  reg  _T_1335; // @[NV_NVDLA_CSC_dl.scala 416:32:@476.4]
  reg [31:0] _RAND_70;
  wire  _T_1357; // @[NV_NVDLA_CSC_dl.scala 424:22:@491.4]
  wire  _T_1358; // @[NV_NVDLA_CSC_dl.scala 423:22:@492.4]
  wire  _T_1299; // @[NV_NVDLA_CSC_dl.scala 391:66:@447.4]
  wire  _T_1300; // @[NV_NVDLA_CSC_dl.scala 391:33:@448.4]
  wire  _T_1301; // @[NV_NVDLA_CSC_dl.scala 393:31:@450.6]
  wire [1:0] _T_1303; // @[NV_NVDLA_CSC_dl.scala 393:21:@451.6]
  wire [1:0] _GEN_65; // @[NV_NVDLA_CSC_dl.scala 392:23:@449.4]
  wire [7:0] _T_1312; // @[NV_NVDLA_CSC_dl.scala 401:33:@457.4]
  wire [6:0] _T_1313; // @[NV_NVDLA_CSC_dl.scala 401:33:@458.4]
  wire  _T_1314; // @[NV_NVDLA_CSC_dl.scala 402:51:@459.4]
  wire  _T_1315; // @[NV_NVDLA_CSC_dl.scala 402:33:@460.4]
  wire  _T_1316; // @[NV_NVDLA_CSC_dl.scala 403:34:@462.4]
  wire  _T_1317; // @[NV_NVDLA_CSC_dl.scala 404:52:@464.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_dl.scala 404:34:@465.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_dl.scala 408:41:@467.6]
  wire  _T_1321; // @[NV_NVDLA_CSC_dl.scala 408:39:@468.6]
  wire [6:0] _T_1324; // @[NV_NVDLA_CSC_dl.scala 409:22:@469.6]
  wire [6:0] _T_1325; // @[NV_NVDLA_CSC_dl.scala 408:22:@470.6]
  wire [6:0] _T_1326; // @[NV_NVDLA_CSC_dl.scala 407:22:@471.6]
  wire [6:0] _GEN_66; // @[NV_NVDLA_CSC_dl.scala 406:24:@466.4]
  reg  _T_1329; // @[NV_NVDLA_CSC_dl.scala 414:35:@474.4]
  reg [31:0] _RAND_71;
  reg  _T_1332; // @[NV_NVDLA_CSC_dl.scala 415:32:@475.4]
  reg [31:0] _RAND_72;
  wire  _T_1343; // @[NV_NVDLA_CSC_dl.scala 422:27:@481.4]
  wire  _T_1338; // @[NV_NVDLA_CSC_dl.scala 419:49:@478.4]
  wire  _T_1341; // @[NV_NVDLA_CSC_dl.scala 420:32:@479.4]
  wire  _T_1342; // @[NV_NVDLA_CSC_dl.scala 419:33:@480.4]
  reg [7:0] _T_1361; // @[NV_NVDLA_CSC_dl.scala 432:31:@497.4]
  reg [31:0] _RAND_73;
  wire [7:0] _T_1363; // @[Cat.scala 30:58:@498.4]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CSC_dl.scala 434:21:@499.4]
  reg [12:0] _T_1366; // @[NV_NVDLA_CSC_dl.scala 440:28:@502.4]
  reg [31:0] _RAND_74;
  reg [12:0] _T_1369; // @[NV_NVDLA_CSC_dl.scala 441:28:@503.4]
  reg [31:0] _RAND_75;
  wire [12:0] _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@504.4]
  wire [13:0] _T_1370; // @[NV_NVDLA_CSC_dl.scala 444:39:@504.4]
  wire [12:0] _T_1371; // @[NV_NVDLA_CSC_dl.scala 444:39:@505.4]
  wire  _T_1372; // @[NV_NVDLA_CSC_dl.scala 445:29:@506.4]
  wire  _T_1373; // @[NV_NVDLA_CSC_dl.scala 445:61:@507.4]
  wire  _T_1374; // @[NV_NVDLA_CSC_dl.scala 445:44:@508.4]
  wire  _T_1377; // @[NV_NVDLA_CSC_dl.scala 448:43:@511.4]
  wire  _T_1378; // @[NV_NVDLA_CSC_dl.scala 448:41:@512.4]
  wire [12:0] _T_1379; // @[NV_NVDLA_CSC_dl.scala 449:26:@513.4]
  wire [12:0] _T_1380; // @[NV_NVDLA_CSC_dl.scala 448:26:@514.4]
  wire [12:0] _T_1381; // @[NV_NVDLA_CSC_dl.scala 447:26:@515.4]
  wire  _T_1383; // @[NV_NVDLA_CSC_dl.scala 450:70:@517.4]
  wire  _T_1384; // @[NV_NVDLA_CSC_dl.scala 450:37:@518.4]
  wire  _T_1385; // @[NV_NVDLA_CSC_dl.scala 451:55:@519.4]
  wire  _T_1386; // @[NV_NVDLA_CSC_dl.scala 451:71:@520.4]
  wire  _T_1387; // @[NV_NVDLA_CSC_dl.scala 451:37:@521.4]
  wire [12:0] _GEN_68; // @[NV_NVDLA_CSC_dl.scala 453:27:@522.4]
  wire [12:0] _GEN_69; // @[NV_NVDLA_CSC_dl.scala 456:27:@525.4]
  reg [10:0] _T_1390; // @[NV_NVDLA_CSC_dl.scala 461:27:@528.4]
  reg [31:0] _RAND_76;
  wire  _T_1391; // @[NV_NVDLA_CSC_dl.scala 463:37:@529.4]
  wire  _T_1393; // @[NV_NVDLA_CSC_dl.scala 464:70:@531.4]
  wire  _T_1394; // @[NV_NVDLA_CSC_dl.scala 464:36:@532.4]
  wire [11:0] _T_1398; // @[NV_NVDLA_CSC_dl.scala 469:34:@534.6]
  wire [10:0] _T_1399; // @[NV_NVDLA_CSC_dl.scala 469:34:@535.6]
  wire [10:0] _T_1400; // @[NV_NVDLA_CSC_dl.scala 468:24:@536.6]
  wire [10:0] _T_1401; // @[NV_NVDLA_CSC_dl.scala 467:24:@537.6]
  wire [10:0] _GEN_70; // @[NV_NVDLA_CSC_dl.scala 466:26:@533.4]
  reg [13:0] _T_1404; // @[NV_NVDLA_CSC_dl.scala 473:27:@540.4]
  reg [31:0] _RAND_77;
  reg [13:0] _T_1407; // @[NV_NVDLA_CSC_dl.scala 474:27:@541.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_1410; // @[NV_NVDLA_CSC_dl.scala 475:26:@542.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_1413; // @[NV_NVDLA_CSC_dl.scala 476:26:@543.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_1416; // @[NV_NVDLA_CSC_dl.scala 477:29:@544.4]
  reg [31:0] _RAND_81;
  reg [12:0] _T_1419; // @[NV_NVDLA_CSC_dl.scala 478:29:@545.4]
  reg [31:0] _RAND_82;
  reg  _T_1424; // @[NV_NVDLA_CSC_dl.scala 480:33:@547.4]
  reg [31:0] _RAND_83;
  reg  _T_1427; // @[NV_NVDLA_CSC_dl.scala 481:35:@548.4]
  reg [31:0] _RAND_84;
  wire [12:0] _GEN_684; // @[NV_NVDLA_CSC_dl.scala 484:41:@549.4]
  wire [13:0] _T_1430; // @[NV_NVDLA_CSC_dl.scala 484:41:@549.4]
  wire [13:0] _T_1431; // @[NV_NVDLA_CSC_dl.scala 484:41:@550.4]
  wire [13:0] _T_1432; // @[NV_NVDLA_CSC_dl.scala 483:26:@551.4]
  wire [13:0] _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@552.4]
  wire [14:0] _T_1433; // @[NV_NVDLA_CSC_dl.scala 485:37:@552.4]
  wire [13:0] _T_1434; // @[NV_NVDLA_CSC_dl.scala 485:37:@553.4]
  wire [13:0] _T_1437; // @[NV_NVDLA_CSC_dl.scala 490:25:@556.4]
  wire [13:0] _T_1438; // @[NV_NVDLA_CSC_dl.scala 489:25:@557.4]
  wire [13:0] _T_1439; // @[NV_NVDLA_CSC_dl.scala 488:25:@558.4]
  wire [5:0] _GEN_686; // @[NV_NVDLA_CSC_dl.scala 492:35:@559.4]
  wire [10:0] _T_1440; // @[NV_NVDLA_CSC_dl.scala 492:35:@559.4]
  wire [13:0] _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@560.4]
  wire [14:0] _T_1441; // @[NV_NVDLA_CSC_dl.scala 493:33:@560.4]
  wire [13:0] _T_1442; // @[NV_NVDLA_CSC_dl.scala 493:33:@561.4]
  wire  _T_1445; // @[NV_NVDLA_CSC_dl.scala 494:96:@564.4]
  wire  _T_1446; // @[NV_NVDLA_CSC_dl.scala 494:86:@565.4]
  wire  _T_1447; // @[NV_NVDLA_CSC_dl.scala 494:84:@566.4]
  wire  _T_1448; // @[NV_NVDLA_CSC_dl.scala 494:36:@567.4]
  wire  _T_1451; // @[NV_NVDLA_CSC_dl.scala 495:99:@570.4]
  wire  _T_1452; // @[NV_NVDLA_CSC_dl.scala 495:89:@571.4]
  wire  _T_1453; // @[NV_NVDLA_CSC_dl.scala 495:87:@572.4]
  wire  _T_1454; // @[NV_NVDLA_CSC_dl.scala 495:36:@573.4]
  wire [7:0] _T_1456; // @[NV_NVDLA_CSC_dl.scala 498:26:@574.4]
  wire  _T_1459; // @[NV_NVDLA_CSC_dl.scala 500:79:@576.4]
  wire [7:0] _T_1463; // @[NV_NVDLA_CSC_dl.scala 501:74:@579.4]
  wire [6:0] _T_1464; // @[NV_NVDLA_CSC_dl.scala 501:74:@580.4]
  wire [6:0] _T_1465; // @[NV_NVDLA_CSC_dl.scala 500:27:@581.4]
  wire  _T_1466; // @[NV_NVDLA_CSC_dl.scala 502:37:@582.4]
  wire  _T_1468; // @[NV_NVDLA_CSC_dl.scala 503:35:@583.4]
  wire [13:0] _T_1470; // @[NV_NVDLA_CSC_dl.scala 503:66:@584.4]
  wire [12:0] _T_1471; // @[NV_NVDLA_CSC_dl.scala 503:66:@585.4]
  wire [12:0] _T_1472; // @[NV_NVDLA_CSC_dl.scala 503:22:@586.4]
  wire [12:0] _T_1473; // @[NV_NVDLA_CSC_dl.scala 502:22:@587.4]
  wire [12:0] _GEN_688; // @[NV_NVDLA_CSC_dl.scala 505:44:@589.4]
  wire  _T_1474; // @[NV_NVDLA_CSC_dl.scala 505:44:@589.4]
  wire  _T_1475; // @[NV_NVDLA_CSC_dl.scala 509:39:@590.4]
  wire  _T_1476; // @[NV_NVDLA_CSC_dl.scala 509:54:@591.4]
  wire  _T_1477; // @[NV_NVDLA_CSC_dl.scala 509:71:@592.4]
  wire  _T_1480; // @[NV_NVDLA_CSC_dl.scala 510:73:@595.4]
  wire  _T_1481; // @[NV_NVDLA_CSC_dl.scala 510:71:@596.4]
  wire [15:0] _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@597.4]
  wire [16:0] _T_1482; // @[NV_NVDLA_CSC_dl.scala 510:99:@597.4]
  wire [15:0] _T_1483; // @[NV_NVDLA_CSC_dl.scala 510:99:@598.4]
  wire  _T_1485; // @[NV_NVDLA_CSC_dl.scala 511:54:@600.4]
  wire [15:0] _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@601.4]
  wire [16:0] _T_1486; // @[NV_NVDLA_CSC_dl.scala 511:90:@601.4]
  wire [15:0] _T_1487; // @[NV_NVDLA_CSC_dl.scala 511:90:@602.4]
  wire  _T_1489; // @[NV_NVDLA_CSC_dl.scala 512:56:@604.4]
  wire  _T_1490; // @[NV_NVDLA_CSC_dl.scala 512:54:@605.4]
  wire [16:0] _T_1492; // @[NV_NVDLA_CSC_dl.scala 512:91:@606.4]
  wire [15:0] _T_1493; // @[NV_NVDLA_CSC_dl.scala 512:91:@607.4]
  wire  _T_1494; // @[NV_NVDLA_CSC_dl.scala 513:41:@608.4]
  wire  _T_1495; // @[NV_NVDLA_CSC_dl.scala 513:39:@609.4]
  wire [15:0] _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@610.4]
  wire [16:0] _T_1496; // @[NV_NVDLA_CSC_dl.scala 513:81:@610.4]
  wire [15:0] _T_1497; // @[NV_NVDLA_CSC_dl.scala 513:81:@611.4]
  wire [15:0] _T_1498; // @[NV_NVDLA_CSC_dl.scala 513:24:@612.4]
  wire [15:0] _T_1499; // @[NV_NVDLA_CSC_dl.scala 512:24:@613.4]
  wire [15:0] _T_1500; // @[NV_NVDLA_CSC_dl.scala 511:24:@614.4]
  wire [15:0] _T_1501; // @[NV_NVDLA_CSC_dl.scala 510:24:@615.4]
  wire [15:0] _T_1502; // @[NV_NVDLA_CSC_dl.scala 509:24:@616.4]
  wire [15:0] _T_1503; // @[NV_NVDLA_CSC_dl.scala 508:24:@617.4]
  wire [9:0] _T_1509; // @[NV_NVDLA_CSC_dl.scala 515:68:@619.4]
  wire [14:0] _T_1510; // @[Cat.scala 30:58:@620.4]
  wire  _T_1521; // @[NV_NVDLA_CSC_dl.scala 518:68:@631.4]
  wire  _T_1522; // @[NV_NVDLA_CSC_dl.scala 518:57:@632.4]
  wire  _T_1523; // @[NV_NVDLA_CSC_dl.scala 518:72:@633.4]
  wire  _T_1524; // @[NV_NVDLA_CSC_dl.scala 518:88:@634.4]
  wire  _T_1525; // @[NV_NVDLA_CSC_dl.scala 518:103:@635.4]
  wire  _T_1526; // @[NV_NVDLA_CSC_dl.scala 518:39:@636.4]
  wire  _T_1528; // @[NV_NVDLA_CSC_dl.scala 520:42:@638.4]
  wire  _T_1531; // @[NV_NVDLA_CSC_dl.scala 520:74:@639.4]
  wire  _T_1532; // @[NV_NVDLA_CSC_dl.scala 520:28:@640.4]
  wire  _T_1534; // @[NV_NVDLA_CSC_dl.scala 521:36:@642.4]
  wire  _T_1535; // @[NV_NVDLA_CSC_dl.scala 521:72:@643.4]
  wire  _T_1536; // @[NV_NVDLA_CSC_dl.scala 521:51:@644.4]
  wire [13:0] _GEN_71; // @[NV_NVDLA_CSC_dl.scala 523:26:@645.4]
  wire [15:0] _GEN_72; // @[NV_NVDLA_CSC_dl.scala 523:26:@645.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CSC_dl.scala 527:26:@649.4]
  wire [15:0] _GEN_74; // @[NV_NVDLA_CSC_dl.scala 527:26:@649.4]
  wire [15:0] _GEN_75; // @[NV_NVDLA_CSC_dl.scala 531:26:@653.4]
  reg [13:0] _T_1539; // @[NV_NVDLA_CSC_dl.scala 537:27:@656.4]
  reg [31:0] _RAND_85;
  reg [13:0] _T_1542; // @[NV_NVDLA_CSC_dl.scala 538:27:@657.4]
  reg [31:0] _RAND_86;
  wire [13:0] _GEN_692; // @[NV_NVDLA_CSC_dl.scala 540:41:@658.4]
  wire [14:0] _T_1544; // @[NV_NVDLA_CSC_dl.scala 540:41:@658.4]
  wire [14:0] _T_1545; // @[NV_NVDLA_CSC_dl.scala 540:41:@659.4]
  wire [13:0] _T_1546; // @[NV_NVDLA_CSC_dl.scala 540:41:@660.4]
  wire [13:0] _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@661.4]
  wire [14:0] _T_1547; // @[NV_NVDLA_CSC_dl.scala 541:37:@661.4]
  wire [13:0] _T_1548; // @[NV_NVDLA_CSC_dl.scala 541:37:@662.4]
  wire  _T_1549; // @[NV_NVDLA_CSC_dl.scala 542:52:@663.4]
  wire  _T_1550; // @[NV_NVDLA_CSC_dl.scala 542:35:@664.4]
  wire [13:0] _T_1553; // @[NV_NVDLA_CSC_dl.scala 544:25:@667.4]
  wire [13:0] _T_1554; // @[NV_NVDLA_CSC_dl.scala 543:25:@668.4]
  wire [13:0] _T_1555; // @[NV_NVDLA_CSC_dl.scala 542:25:@669.4]
  wire  _T_1558; // @[NV_NVDLA_CSC_dl.scala 545:91:@672.4]
  wire  _T_1559; // @[NV_NVDLA_CSC_dl.scala 545:54:@673.4]
  wire  _T_1560; // @[NV_NVDLA_CSC_dl.scala 545:36:@674.4]
  wire [5:0] _GEN_694; // @[NV_NVDLA_CSC_dl.scala 547:35:@678.4]
  wire [10:0] _T_1564; // @[NV_NVDLA_CSC_dl.scala 547:35:@678.4]
  wire [13:0] _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@679.4]
  wire [14:0] _T_1565; // @[NV_NVDLA_CSC_dl.scala 548:33:@679.4]
  wire [13:0] _T_1566; // @[NV_NVDLA_CSC_dl.scala 548:33:@680.4]
  wire [13:0] _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@681.4]
  wire [14:0] _T_1567; // @[NV_NVDLA_CSC_dl.scala 548:51:@681.4]
  wire [13:0] _T_1568; // @[NV_NVDLA_CSC_dl.scala 548:51:@682.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CSC_dl.scala 550:26:@683.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CSC_dl.scala 551:26:@686.4]
  wire  _T_1569; // @[NV_NVDLA_CSC_dl.scala 554:39:@689.4]
  wire [13:0] _GEN_697; // @[NV_NVDLA_CSC_dl.scala 554:59:@690.4]
  wire  _T_1570; // @[NV_NVDLA_CSC_dl.scala 554:59:@690.4]
  wire  _T_1571; // @[NV_NVDLA_CSC_dl.scala 554:44:@691.4]
  wire  _T_1572; // @[NV_NVDLA_CSC_dl.scala 554:92:@692.4]
  wire  _T_1573; // @[NV_NVDLA_CSC_dl.scala 554:78:@693.4]
  wire [13:0] _GEN_698; // @[NV_NVDLA_CSC_dl.scala 554:112:@694.4]
  wire  _T_1574; // @[NV_NVDLA_CSC_dl.scala 554:112:@694.4]
  wire  _T_1575; // @[NV_NVDLA_CSC_dl.scala 554:97:@695.4]
  wire  _T_1588; // @[NV_NVDLA_CSC_dl.scala 557:42:@705.4]
  wire  _T_1698; // @[NV_NVDLA_CSC_dl.scala 642:33:@791.4]
  wire  _T_1699; // @[NV_NVDLA_CSC_dl.scala 643:24:@792.4]
  wire [12:0] _T_1701; // @[NV_NVDLA_CSC_dl.scala 643:77:@793.4]
  wire [14:0] _T_1702; // @[Cat.scala 30:58:@794.4]
  wire  _T_1704; // @[NV_NVDLA_CSC_dl.scala 644:38:@795.4]
  wire [11:0] _T_1709; // @[NV_NVDLA_CSC_dl.scala 645:54:@798.4]
  wire [14:0] _T_1710; // @[Cat.scala 30:58:@799.4]
  wire [14:0] _T_1711; // @[NV_NVDLA_CSC_dl.scala 644:23:@800.4]
  wire [14:0] _T_1712; // @[NV_NVDLA_CSC_dl.scala 643:23:@801.4]
  wire [14:0] _T_1713; // @[NV_NVDLA_CSC_dl.scala 642:23:@802.4]
  wire [13:0] _T_1714; // @[NV_NVDLA_CSC_dl.scala 654:24:@804.4]
  wire [11:0] _T_1591; // @[NV_NVDLA_CSC_dl.scala 561:32:@707.4]
  wire [14:0] _GEN_700; // @[NV_NVDLA_CSC_dl.scala 561:40:@708.4]
  wire  _T_1592; // @[NV_NVDLA_CSC_dl.scala 561:40:@708.4]
  wire  _T_1593; // @[NV_NVDLA_CSC_dl.scala 562:34:@709.4]
  wire  _T_1594; // @[NV_NVDLA_CSC_dl.scala 562:24:@710.4]
  wire  _T_1595; // @[NV_NVDLA_CSC_dl.scala 563:29:@711.4]
  wire  _T_1596; // @[NV_NVDLA_CSC_dl.scala 563:33:@712.4]
  wire  _T_1597; // @[NV_NVDLA_CSC_dl.scala 564:39:@713.4]
  wire  _T_1598; // @[NV_NVDLA_CSC_dl.scala 564:37:@714.4]
  wire  _T_1599; // @[NV_NVDLA_CSC_dl.scala 564:56:@715.4]
  wire  _T_1600; // @[NV_NVDLA_CSC_dl.scala 564:54:@716.4]
  wire  _T_1601; // @[NV_NVDLA_CSC_dl.scala 567:37:@717.4]
  wire  _T_1602; // @[NV_NVDLA_CSC_dl.scala 567:27:@718.4]
  wire  _T_1603; // @[NV_NVDLA_CSC_dl.scala 567:54:@719.4]
  wire  _T_1604; // @[NV_NVDLA_CSC_dl.scala 567:26:@720.4]
  wire [1:0] _T_1605; // @[NV_NVDLA_CSC_dl.scala 568:35:@721.4]
  wire  _T_1607; // @[NV_NVDLA_CSC_dl.scala 569:55:@722.4]
  wire  _T_1608; // @[NV_NVDLA_CSC_dl.scala 569:42:@723.4]
  wire  _T_1609; // @[NV_NVDLA_CSC_dl.scala 572:42:@725.4]
  wire [8:0] _T_1613; // @[Cat.scala 30:58:@729.4]
  reg  _T_1616; // @[NV_NVDLA_CSC_dl.scala 579:31:@730.4]
  reg [31:0] _RAND_87;
  reg [1:0] _T_1619; // @[NV_NVDLA_CSC_dl.scala 580:31:@731.4]
  reg [31:0] _RAND_88;
  reg [1:0] _T_1622; // @[NV_NVDLA_CSC_dl.scala 581:31:@732.4]
  reg [31:0] _RAND_89;
  reg  _T_1625; // @[NV_NVDLA_CSC_dl.scala 582:31:@733.4]
  reg [31:0] _RAND_90;
  reg  _T_1628; // @[NV_NVDLA_CSC_dl.scala 583:32:@734.4]
  reg [31:0] _RAND_91;
  reg  _T_1631; // @[NV_NVDLA_CSC_dl.scala 584:31:@735.4]
  reg [31:0] _RAND_92;
  reg [1:0] _T_1634; // @[NV_NVDLA_CSC_dl.scala 585:35:@736.4]
  reg [31:0] _RAND_93;
  reg  _T_1637; // @[NV_NVDLA_CSC_dl.scala 586:34:@737.4]
  reg [31:0] _RAND_94;
  reg [8:0] _T_1640; // @[NV_NVDLA_CSC_dl.scala 587:30:@738.4]
  reg [31:0] _RAND_95;
  reg  _T_1643; // @[NV_NVDLA_CSC_dl.scala 588:29:@739.4]
  reg [31:0] _RAND_96;
  wire  _T_1644; // @[NV_NVDLA_CSC_dl.scala 599:38:@749.6]
  wire  _T_1645; // @[NV_NVDLA_CSC_dl.scala 599:56:@750.6]
  wire [1:0] _GEN_78; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire [1:0] _GEN_79; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_80; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_81; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_82; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire [8:0] _GEN_84; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_87; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  wire  _GEN_88; // @[NV_NVDLA_CSC_dl.scala 603:26:@755.4]
  reg [12:0] _T_1648; // @[NV_NVDLA_CSC_dl.scala 611:21:@758.4]
  reg [31:0] _RAND_97;
  reg [12:0] _T_1651; // @[NV_NVDLA_CSC_dl.scala 612:24:@759.4]
  reg [31:0] _RAND_98;
  reg [12:0] _T_1654; // @[NV_NVDLA_CSC_dl.scala 613:26:@760.4]
  reg [31:0] _RAND_99;
  reg [12:0] _T_1657; // @[NV_NVDLA_CSC_dl.scala 614:26:@761.4]
  reg [31:0] _RAND_100;
  reg [12:0] _T_1660; // @[NV_NVDLA_CSC_dl.scala 615:26:@762.4]
  reg [31:0] _RAND_101;
  reg [12:0] _T_1663; // @[NV_NVDLA_CSC_dl.scala 616:26:@763.4]
  reg [31:0] _RAND_102;
  reg [12:0] _T_1666; // @[NV_NVDLA_CSC_dl.scala 617:24:@764.4]
  reg [31:0] _RAND_103;
  wire  _T_1667; // @[NV_NVDLA_CSC_dl.scala 620:32:@765.4]
  wire  _T_1668; // @[NV_NVDLA_CSC_dl.scala 620:22:@766.4]
  wire [11:0] _T_1669; // @[NV_NVDLA_CSC_dl.scala 620:49:@767.4]
  wire [11:0] _T_1671; // @[NV_NVDLA_CSC_dl.scala 620:21:@768.4]
  wire  _T_1673; // @[NV_NVDLA_CSC_dl.scala 622:34:@769.4]
  wire [12:0] _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@770.4]
  wire [13:0] _T_1675; // @[NV_NVDLA_CSC_dl.scala 622:64:@770.4]
  wire [12:0] _T_1676; // @[NV_NVDLA_CSC_dl.scala 622:64:@771.4]
  wire [12:0] _T_1677; // @[NV_NVDLA_CSC_dl.scala 622:19:@772.4]
  wire [12:0] _T_1678; // @[NV_NVDLA_CSC_dl.scala 621:19:@773.4]
  wire  _T_1682; // @[NV_NVDLA_CSC_dl.scala 624:31:@777.4]
  wire [13:0] _GEN_702; // @[NV_NVDLA_CSC_dl.scala 627:32:@778.4]
  wire [25:0] _T_1683; // @[NV_NVDLA_CSC_dl.scala 627:32:@778.4]
  wire [12:0] _T_1684; // @[NV_NVDLA_CSC_dl.scala 627:50:@779.4]
  wire [11:0] _GEN_703; // @[NV_NVDLA_CSC_dl.scala 628:31:@780.4]
  wire [16:0] _T_1685; // @[NV_NVDLA_CSC_dl.scala 628:31:@780.4]
  wire [12:0] _T_1686; // @[NV_NVDLA_CSC_dl.scala 628:49:@781.4]
  wire [14:0] _GEN_704; // @[NV_NVDLA_CSC_dl.scala 629:29:@782.4]
  wire [19:0] _T_1687; // @[NV_NVDLA_CSC_dl.scala 629:29:@782.4]
  wire [12:0] _T_1688; // @[NV_NVDLA_CSC_dl.scala 629:47:@783.4]
  wire [14:0] _GEN_705; // @[NV_NVDLA_CSC_dl.scala 630:47:@784.4]
  wire [16:0] _T_1690; // @[NV_NVDLA_CSC_dl.scala 630:47:@784.4]
  wire [16:0] _T_1691; // @[NV_NVDLA_CSC_dl.scala 630:21:@785.4]
  wire [12:0] _T_1692; // @[NV_NVDLA_CSC_dl.scala 630:65:@786.4]
  wire  _T_1693; // @[NV_NVDLA_CSC_dl.scala 631:45:@787.4]
  wire  _T_1694; // @[NV_NVDLA_CSC_dl.scala 631:34:@788.4]
  wire [1:0] _T_1695; // @[Cat.scala 30:58:@789.4]
  wire [12:0] _GEN_89; // @[NV_NVDLA_CSC_dl.scala 658:20:@806.4]
  wire [12:0] _GEN_90; // @[NV_NVDLA_CSC_dl.scala 661:23:@809.4]
  wire  _T_1715; // @[NV_NVDLA_CSC_dl.scala 664:19:@812.4]
  wire [12:0] _GEN_91; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  wire [12:0] _GEN_92; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  wire  _T_1716; // @[NV_NVDLA_CSC_dl.scala 669:19:@818.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl.scala 669:23:@819.4]
  wire [13:0] _GEN_95; // @[NV_NVDLA_CSC_dl.scala 672:20:@822.4]
  reg [12:0] _T_1759_0; // @[NV_NVDLA_CSC_dl.scala 680:33:@834.4]
  reg [31:0] _RAND_104;
  reg [12:0] _T_1759_1; // @[NV_NVDLA_CSC_dl.scala 680:33:@834.4]
  reg [31:0] _RAND_105;
  reg [12:0] _T_1759_2; // @[NV_NVDLA_CSC_dl.scala 680:33:@834.4]
  reg [31:0] _RAND_106;
  reg [12:0] _T_1759_3; // @[NV_NVDLA_CSC_dl.scala 680:33:@834.4]
  reg [31:0] _RAND_107;
  reg  _T_1778; // @[NV_NVDLA_CSC_dl.scala 681:35:@835.4]
  reg [31:0] _RAND_108;
  reg [14:0] _T_1785; // @[NV_NVDLA_CSC_dl.scala 682:37:@837.4]
  reg [31:0] _RAND_109;
  reg  _T_1788; // @[NV_NVDLA_CSC_dl.scala 683:32:@838.4]
  reg [31:0] _RAND_110;
  reg [1:0] _T_1794; // @[NV_NVDLA_CSC_dl.scala 685:33:@840.4]
  reg [31:0] _RAND_111;
  reg [1:0] _T_1797; // @[NV_NVDLA_CSC_dl.scala 686:33:@841.4]
  reg [31:0] _RAND_112;
  reg  _T_1800; // @[NV_NVDLA_CSC_dl.scala 687:33:@842.4]
  reg [31:0] _RAND_113;
  reg  _T_1803; // @[NV_NVDLA_CSC_dl.scala 688:34:@843.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_1806; // @[NV_NVDLA_CSC_dl.scala 689:33:@844.4]
  reg [31:0] _RAND_115;
  reg  _T_1809; // @[NV_NVDLA_CSC_dl.scala 690:33:@845.4]
  reg [31:0] _RAND_116;
  reg [1:0] _T_1812; // @[NV_NVDLA_CSC_dl.scala 691:37:@846.4]
  reg [31:0] _RAND_117;
  reg  _T_1815; // @[NV_NVDLA_CSC_dl.scala 692:36:@847.4]
  reg [31:0] _RAND_118;
  reg  _T_1818; // @[NV_NVDLA_CSC_dl.scala 693:31:@848.4]
  reg [31:0] _RAND_119;
  reg [8:0] _T_1821; // @[NV_NVDLA_CSC_dl.scala 694:32:@849.4]
  reg [31:0] _RAND_120;
  wire [13:0] _T_1822; // @[NV_NVDLA_CSC_dl.scala 696:29:@850.4]
  wire [12:0] _T_1823; // @[NV_NVDLA_CSC_dl.scala 696:29:@851.4]
  wire [13:0] _T_1824; // @[NV_NVDLA_CSC_dl.scala 696:43:@852.4]
  wire [12:0] _T_1825; // @[NV_NVDLA_CSC_dl.scala 696:43:@853.4]
  wire [13:0] _T_1826; // @[NV_NVDLA_CSC_dl.scala 696:57:@854.4]
  wire [12:0] _T_1827; // @[NV_NVDLA_CSC_dl.scala 696:57:@855.4]
  wire [14:0] _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@856.4]
  wire [15:0] _T_1828; // @[NV_NVDLA_CSC_dl.scala 697:40:@856.4]
  wire [14:0] _T_1829; // @[NV_NVDLA_CSC_dl.scala 697:40:@857.4]
  wire [14:0] _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@858.4]
  wire [15:0] _T_1830; // @[NV_NVDLA_CSC_dl.scala 697:52:@858.4]
  wire [14:0] _T_1831; // @[NV_NVDLA_CSC_dl.scala 697:52:@859.4]
  wire [14:0] _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@860.4]
  wire [15:0] _T_1832; // @[NV_NVDLA_CSC_dl.scala 697:64:@860.4]
  wire [14:0] _T_1833; // @[NV_NVDLA_CSC_dl.scala 697:64:@861.4]
  wire  _T_1840; // @[NV_NVDLA_CSC_dl.scala 698:45:@864.4]
  wire [15:0] _T_1847; // @[NV_NVDLA_CSC_dl.scala 699:42:@867.4]
  wire [15:0] _T_1848; // @[NV_NVDLA_CSC_dl.scala 699:42:@868.4]
  wire [14:0] _T_1849; // @[NV_NVDLA_CSC_dl.scala 699:42:@869.4]
  wire  _T_1850; // @[NV_NVDLA_CSC_dl.scala 700:35:@870.4]
  wire [14:0] _T_1856; // @[NV_NVDLA_CSC_dl.scala 701:25:@872.4]
  wire [14:0] _T_1857; // @[NV_NVDLA_CSC_dl.scala 700:25:@873.4]
  wire  _T_1881; // @[Mux.scala 46:19:@883.4]
  wire [12:0] _T_1882; // @[Mux.scala 46:16:@884.4]
  wire  _T_1883; // @[Mux.scala 46:19:@885.4]
  wire [12:0] _T_1884; // @[Mux.scala 46:16:@886.4]
  wire  _T_1885; // @[Mux.scala 46:19:@887.4]
  wire [12:0] _T_1886; // @[Mux.scala 46:16:@888.4]
  wire  _T_1887; // @[Mux.scala 46:19:@889.4]
  wire [12:0] _T_1888; // @[Mux.scala 46:16:@890.4]
  wire [14:0] _GEN_712; // @[NV_NVDLA_CSC_dl.scala 708:65:@891.4]
  wire  _T_1889; // @[NV_NVDLA_CSC_dl.scala 708:65:@891.4]
  wire  _T_1890; // @[NV_NVDLA_CSC_dl.scala 708:85:@892.4]
  wire  _T_1891; // @[NV_NVDLA_CSC_dl.scala 708:43:@893.4]
  wire  _T_1892; // @[NV_NVDLA_CSC_dl.scala 710:38:@894.4]
  wire  _T_1894; // @[NV_NVDLA_CSC_dl.scala 710:78:@895.4]
  wire  _T_1895; // @[NV_NVDLA_CSC_dl.scala 710:58:@896.4]
  wire  _T_1896; // @[NV_NVDLA_CSC_dl.scala 710:17:@897.4]
  wire  _T_1899; // @[NV_NVDLA_CSC_dl.scala 710:78:@899.4]
  wire  _T_1900; // @[NV_NVDLA_CSC_dl.scala 710:58:@900.4]
  wire  _T_1901; // @[NV_NVDLA_CSC_dl.scala 710:17:@901.4]
  wire  _T_1904; // @[NV_NVDLA_CSC_dl.scala 710:78:@903.4]
  wire  _T_1905; // @[NV_NVDLA_CSC_dl.scala 710:58:@904.4]
  wire  _T_1906; // @[NV_NVDLA_CSC_dl.scala 710:17:@905.4]
  wire  _T_1909; // @[NV_NVDLA_CSC_dl.scala 710:78:@907.4]
  wire  _T_1910; // @[NV_NVDLA_CSC_dl.scala 710:58:@908.4]
  wire  _T_1911; // @[NV_NVDLA_CSC_dl.scala 710:17:@909.4]
  wire [14:0] _GEN_96; // @[NV_NVDLA_CSC_dl.scala 717:35:@915.4]
  wire [14:0] _GEN_97; // @[NV_NVDLA_CSC_dl.scala 717:35:@918.4]
  wire [14:0] _GEN_98; // @[NV_NVDLA_CSC_dl.scala 717:35:@921.4]
  wire [14:0] _GEN_99; // @[NV_NVDLA_CSC_dl.scala 717:35:@924.4]
  wire  _T_1922; // @[NV_NVDLA_CSC_dl.scala 723:14:@928.4]
  wire [14:0] _GEN_100; // @[NV_NVDLA_CSC_dl.scala 723:34:@929.4]
  wire [1:0] _GEN_101; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire [1:0] _GEN_102; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire  _GEN_103; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire  _GEN_104; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire  _GEN_106; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire [1:0] _GEN_107; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire  _GEN_109; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire [8:0] _GEN_110; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  wire [6:0] _T_1932; // @[Cat.scala 30:58:@956.4]
  wire [28:0] _T_1938; // @[Cat.scala 30:58:@962.4]
  reg  _T_1943; // @[NV_NVDLA_CSC_dl.scala 757:73:@964.4]
  reg [31:0] _RAND_121;
  reg  _T_1946; // @[NV_NVDLA_CSC_dl.scala 757:73:@965.4]
  reg [31:0] _RAND_122;
  reg  _T_1949; // @[NV_NVDLA_CSC_dl.scala 757:73:@966.4]
  reg [31:0] _RAND_123;
  reg  _T_1952; // @[NV_NVDLA_CSC_dl.scala 757:73:@967.4]
  reg [31:0] _RAND_124;
  reg  _T_1955; // @[NV_NVDLA_CSC_dl.scala 757:73:@968.4]
  reg [31:0] _RAND_125;
  reg  _T_1958; // @[NV_NVDLA_CSC_dl.scala 757:73:@969.4]
  reg [31:0] _RAND_126;
  reg [28:0] _T_1963; // @[NV_NVDLA_CSC_dl.scala 759:71:@971.4]
  reg [31:0] _RAND_127;
  reg [28:0] _T_1966; // @[NV_NVDLA_CSC_dl.scala 759:71:@972.4]
  reg [31:0] _RAND_128;
  reg [28:0] _T_1969; // @[NV_NVDLA_CSC_dl.scala 759:71:@973.4]
  reg [31:0] _RAND_129;
  reg [28:0] _T_1972; // @[NV_NVDLA_CSC_dl.scala 759:71:@974.4]
  reg [31:0] _RAND_130;
  reg [28:0] _T_1975; // @[NV_NVDLA_CSC_dl.scala 759:71:@975.4]
  reg [31:0] _RAND_131;
  reg [28:0] _T_1978; // @[NV_NVDLA_CSC_dl.scala 759:71:@976.4]
  reg [31:0] _RAND_132;
  wire [28:0] _GEN_111; // @[NV_NVDLA_CSC_dl.scala 775:33:@1004.4]
  wire [28:0] _GEN_114; // @[NV_NVDLA_CSC_dl.scala 775:33:@1013.4]
  wire [28:0] _GEN_117; // @[NV_NVDLA_CSC_dl.scala 775:33:@1022.4]
  wire [28:0] _GEN_120; // @[NV_NVDLA_CSC_dl.scala 775:33:@1031.4]
  wire [28:0] _GEN_123; // @[NV_NVDLA_CSC_dl.scala 775:33:@1040.4]
  wire [28:0] _GEN_126; // @[NV_NVDLA_CSC_dl.scala 775:33:@1049.4]
  wire [1:0] _T_2039; // @[NV_NVDLA_CSC_dl.scala 792:41:@1057.4]
  wire [1:0] _T_2040; // @[NV_NVDLA_CSC_dl.scala 793:41:@1058.4]
  wire  _T_2041; // @[NV_NVDLA_CSC_dl.scala 794:41:@1059.4]
  wire  _T_2042; // @[NV_NVDLA_CSC_dl.scala 795:42:@1060.4]
  wire [7:0] _T_2043; // @[NV_NVDLA_CSC_dl.scala 796:41:@1061.4]
  wire [1:0] _T_2044; // @[NV_NVDLA_CSC_dl.scala 797:45:@1062.4]
  wire  _T_2047; // @[NV_NVDLA_CSC_dl.scala 800:39:@1065.4]
  wire [8:0] _T_2048; // @[NV_NVDLA_CSC_dl.scala 801:40:@1066.4]
  reg  _T_2051; // @[NV_NVDLA_CSC_dl.scala 806:29:@1067.4]
  reg [31:0] _RAND_133;
  reg  _T_2063; // @[NV_NVDLA_CSC_dl.scala 810:29:@1071.4]
  reg [31:0] _RAND_134;
  reg [511:0] _T_2074; // @[NV_NVDLA_CSC_dl.scala 815:19:@1075.4]
  reg [511:0] _RAND_135;
  reg [511:0] _T_2082; // @[NV_NVDLA_CSC_dl.scala 819:19:@1079.4]
  reg [511:0] _RAND_136;
  wire  _T_2105; // @[NV_NVDLA_CSC_dl.scala 831:69:@1094.4]
  wire  _T_2106; // @[NV_NVDLA_CSC_dl.scala 831:74:@1095.4]
  wire  _T_2107; // @[NV_NVDLA_CSC_dl.scala 831:90:@1096.4]
  wire  _T_2108; // @[NV_NVDLA_CSC_dl.scala 831:88:@1097.4]
  wire  _T_2148; // @[NV_NVDLA_CSC_dl.scala 846:22:@1131.4]
  wire  _T_2162; // @[NV_NVDLA_CSC_dl.scala 850:48:@1142.4]
  wire  _T_2163; // @[NV_NVDLA_CSC_dl.scala 850:22:@1143.4]
  reg [7:0] _T_2182; // @[NV_NVDLA_CSC_dl.scala 867:29:@1184.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_2185; // @[NV_NVDLA_CSC_dl.scala 868:29:@1185.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_2188; // @[NV_NVDLA_CSC_dl.scala 869:29:@1186.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_2191; // @[NV_NVDLA_CSC_dl.scala 870:29:@1187.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_2194; // @[NV_NVDLA_CSC_dl.scala 871:33:@1188.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_2197; // @[NV_NVDLA_CSC_dl.scala 872:33:@1189.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_2200; // @[NV_NVDLA_CSC_dl.scala 873:33:@1190.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_2203; // @[NV_NVDLA_CSC_dl.scala 874:33:@1191.4]
  reg [31:0] _RAND_144;
  reg  _T_2214; // @[NV_NVDLA_CSC_dl.scala 879:41:@1195.4]
  reg [31:0] _RAND_145;
  reg [26:0] _T_2228; // @[NV_NVDLA_CSC_dl.scala 881:41:@1200.4]
  reg [31:0] _RAND_146;
  wire [26:0] _T_2240; // @[Cat.scala 30:58:@1210.4]
  wire [26:0] _GEN_137; // @[NV_NVDLA_CSC_dl.scala 889:28:@1213.4]
  wire [26:0] _GEN_138; // @[NV_NVDLA_CSC_dl.scala 889:28:@1217.4]
  wire [26:0] _GEN_139; // @[NV_NVDLA_CSC_dl.scala 889:28:@1221.4]
  wire [26:0] _GEN_140; // @[NV_NVDLA_CSC_dl.scala 889:28:@1225.4]
  wire  _T_2269; // @[NV_NVDLA_CSC_dl.scala 907:39:@1251.4]
  wire  _T_2270; // @[NV_NVDLA_CSC_dl.scala 908:39:@1252.4]
  wire  _T_2271; // @[NV_NVDLA_CSC_dl.scala 909:39:@1253.4]
  wire  _T_2272; // @[NV_NVDLA_CSC_dl.scala 910:39:@1254.4]
  wire [8:0] _T_2273; // @[NV_NVDLA_CSC_dl.scala 912:38:@1255.4]
  wire [8:0] _T_2274; // @[NV_NVDLA_CSC_dl.scala 913:38:@1256.4]
  wire [8:0] _T_2275; // @[NV_NVDLA_CSC_dl.scala 914:38:@1257.4]
  wire [8:0] _T_2276; // @[NV_NVDLA_CSC_dl.scala 915:38:@1258.4]
  wire  _T_2277; // @[NV_NVDLA_CSC_dl.scala 917:44:@1259.4]
  wire  _T_2278; // @[NV_NVDLA_CSC_dl.scala 918:44:@1260.4]
  wire  _T_2279; // @[NV_NVDLA_CSC_dl.scala 919:44:@1261.4]
  wire  _T_2280; // @[NV_NVDLA_CSC_dl.scala 920:44:@1262.4]
  wire [1:0] _T_2281; // @[NV_NVDLA_CSC_dl.scala 923:31:@1263.4]
  wire [7:0] _T_2285; // @[NV_NVDLA_CSC_dl.scala 927:31:@1267.4]
  wire [1:0] _T_2286; // @[NV_NVDLA_CSC_dl.scala 928:35:@1268.4]
  wire [7:0] _T_2296; // @[NV_NVDLA_CSC_dl.scala 939:29:@1277.4]
  wire  _T_2307; // @[NV_NVDLA_CSC_dl.scala 944:50:@1281.4]
  wire [7:0] _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@1282.4]
  wire [8:0] _T_2309; // @[NV_NVDLA_CSC_dl.scala 944:111:@1282.4]
  wire [7:0] _T_2310; // @[NV_NVDLA_CSC_dl.scala 944:111:@1283.4]
  wire [8:0] _T_2311; // @[NV_NVDLA_CSC_dl.scala 944:133:@1284.4]
  wire [8:0] _T_2312; // @[NV_NVDLA_CSC_dl.scala 944:133:@1285.4]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_dl.scala 944:133:@1286.4]
  wire [7:0] _T_2314; // @[NV_NVDLA_CSC_dl.scala 944:29:@1287.4]
  wire [8:0] _T_2318; // @[NV_NVDLA_CSC_dl.scala 945:111:@1289.4]
  wire [7:0] _T_2319; // @[NV_NVDLA_CSC_dl.scala 945:111:@1290.4]
  wire [8:0] _T_2320; // @[NV_NVDLA_CSC_dl.scala 945:133:@1291.4]
  wire [8:0] _T_2321; // @[NV_NVDLA_CSC_dl.scala 945:133:@1292.4]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_dl.scala 945:133:@1293.4]
  wire [7:0] _T_2323; // @[NV_NVDLA_CSC_dl.scala 945:29:@1294.4]
  wire [8:0] _T_2327; // @[NV_NVDLA_CSC_dl.scala 946:111:@1296.4]
  wire [7:0] _T_2328; // @[NV_NVDLA_CSC_dl.scala 946:111:@1297.4]
  wire [8:0] _T_2329; // @[NV_NVDLA_CSC_dl.scala 946:133:@1298.4]
  wire [8:0] _T_2330; // @[NV_NVDLA_CSC_dl.scala 946:133:@1299.4]
  wire [7:0] _T_2331; // @[NV_NVDLA_CSC_dl.scala 946:133:@1300.4]
  wire [7:0] _T_2332; // @[NV_NVDLA_CSC_dl.scala 946:29:@1301.4]
  wire [8:0] _T_2336; // @[NV_NVDLA_CSC_dl.scala 947:111:@1303.4]
  wire [7:0] _T_2337; // @[NV_NVDLA_CSC_dl.scala 947:111:@1304.4]
  wire [8:0] _T_2338; // @[NV_NVDLA_CSC_dl.scala 947:133:@1305.4]
  wire [8:0] _T_2339; // @[NV_NVDLA_CSC_dl.scala 947:133:@1306.4]
  wire [7:0] _T_2340; // @[NV_NVDLA_CSC_dl.scala 947:133:@1307.4]
  wire [7:0] _T_2341; // @[NV_NVDLA_CSC_dl.scala 947:29:@1308.4]
  wire  _T_2343; // @[NV_NVDLA_CSC_dl.scala 956:52:@1309.4]
  wire  _T_2344; // @[NV_NVDLA_CSC_dl.scala 956:50:@1310.4]
  wire  _T_2345; // @[NV_NVDLA_CSC_dl.scala 957:50:@1311.4]
  wire [7:0] _T_2350; // @[NV_NVDLA_CSC_dl.scala 957:27:@1314.4]
  wire [7:0] _T_2351; // @[NV_NVDLA_CSC_dl.scala 956:27:@1315.4]
  wire [7:0] _T_2352; // @[NV_NVDLA_CSC_dl.scala 955:27:@1316.4]
  wire  _T_2354; // @[NV_NVDLA_CSC_dl.scala 961:52:@1317.4]
  wire  _T_2355; // @[NV_NVDLA_CSC_dl.scala 961:50:@1318.4]
  wire  _T_2356; // @[NV_NVDLA_CSC_dl.scala 962:50:@1319.4]
  wire [7:0] _T_2361; // @[NV_NVDLA_CSC_dl.scala 962:27:@1322.4]
  wire [7:0] _T_2362; // @[NV_NVDLA_CSC_dl.scala 961:27:@1323.4]
  wire [7:0] _T_2363; // @[NV_NVDLA_CSC_dl.scala 960:27:@1324.4]
  wire  _T_2365; // @[NV_NVDLA_CSC_dl.scala 966:52:@1325.4]
  wire  _T_2366; // @[NV_NVDLA_CSC_dl.scala 966:50:@1326.4]
  wire  _T_2367; // @[NV_NVDLA_CSC_dl.scala 967:50:@1327.4]
  wire [7:0] _T_2372; // @[NV_NVDLA_CSC_dl.scala 967:27:@1330.4]
  wire [7:0] _T_2373; // @[NV_NVDLA_CSC_dl.scala 966:27:@1331.4]
  wire [7:0] _T_2374; // @[NV_NVDLA_CSC_dl.scala 965:27:@1332.4]
  wire  _T_2376; // @[NV_NVDLA_CSC_dl.scala 971:52:@1333.4]
  wire  _T_2377; // @[NV_NVDLA_CSC_dl.scala 971:50:@1334.4]
  wire  _T_2378; // @[NV_NVDLA_CSC_dl.scala 972:50:@1335.4]
  wire [7:0] _T_2383; // @[NV_NVDLA_CSC_dl.scala 972:27:@1338.4]
  wire [7:0] _T_2384; // @[NV_NVDLA_CSC_dl.scala 971:27:@1339.4]
  wire [7:0] _T_2385; // @[NV_NVDLA_CSC_dl.scala 970:27:@1340.4]
  wire  _T_2386; // @[NV_NVDLA_CSC_dl.scala 976:46:@1341.4]
  wire  _T_2387; // @[NV_NVDLA_CSC_dl.scala 976:51:@1342.4]
  wire  _T_2388; // @[NV_NVDLA_CSC_dl.scala 976:34:@1343.4]
  wire  _T_2389; // @[NV_NVDLA_CSC_dl.scala 977:46:@1344.4]
  wire  _T_2390; // @[NV_NVDLA_CSC_dl.scala 977:51:@1345.4]
  wire  _T_2392; // @[NV_NVDLA_CSC_dl.scala 977:87:@1346.4]
  wire  _T_2393; // @[NV_NVDLA_CSC_dl.scala 977:69:@1347.4]
  wire  _T_2394; // @[NV_NVDLA_CSC_dl.scala 977:34:@1348.4]
  wire  _T_2395; // @[NV_NVDLA_CSC_dl.scala 978:46:@1349.4]
  wire  _T_2396; // @[NV_NVDLA_CSC_dl.scala 978:51:@1350.4]
  wire  _T_2398; // @[NV_NVDLA_CSC_dl.scala 978:87:@1351.4]
  wire  _T_2399; // @[NV_NVDLA_CSC_dl.scala 978:69:@1352.4]
  wire  _T_2400; // @[NV_NVDLA_CSC_dl.scala 978:34:@1353.4]
  wire  _T_2401; // @[NV_NVDLA_CSC_dl.scala 979:46:@1354.4]
  wire  _T_2402; // @[NV_NVDLA_CSC_dl.scala 979:51:@1355.4]
  wire  _T_2405; // @[NV_NVDLA_CSC_dl.scala 979:69:@1357.4]
  wire  _T_2406; // @[NV_NVDLA_CSC_dl.scala 979:34:@1358.4]
  wire  _T_2407; // @[NV_NVDLA_CSC_dl.scala 981:50:@1359.4]
  wire  _T_2408; // @[NV_NVDLA_CSC_dl.scala 981:55:@1360.4]
  wire  _T_2409; // @[NV_NVDLA_CSC_dl.scala 981:73:@1361.4]
  wire  _T_2410; // @[NV_NVDLA_CSC_dl.scala 981:97:@1362.4]
  wire  _T_2411; // @[NV_NVDLA_CSC_dl.scala 981:38:@1363.4]
  wire  _T_2412; // @[NV_NVDLA_CSC_dl.scala 982:50:@1364.4]
  wire  _T_2413; // @[NV_NVDLA_CSC_dl.scala 982:55:@1365.4]
  wire  _T_2414; // @[NV_NVDLA_CSC_dl.scala 982:73:@1366.4]
  wire  _T_2415; // @[NV_NVDLA_CSC_dl.scala 982:97:@1367.4]
  wire  _T_2417; // @[NV_NVDLA_CSC_dl.scala 982:138:@1368.4]
  wire  _T_2418; // @[NV_NVDLA_CSC_dl.scala 982:120:@1369.4]
  wire  _T_2419; // @[NV_NVDLA_CSC_dl.scala 982:38:@1370.4]
  wire  _T_2420; // @[NV_NVDLA_CSC_dl.scala 983:50:@1371.4]
  wire  _T_2421; // @[NV_NVDLA_CSC_dl.scala 983:55:@1372.4]
  wire  _T_2422; // @[NV_NVDLA_CSC_dl.scala 983:73:@1373.4]
  wire  _T_2423; // @[NV_NVDLA_CSC_dl.scala 983:97:@1374.4]
  wire  _T_2425; // @[NV_NVDLA_CSC_dl.scala 983:138:@1375.4]
  wire  _T_2426; // @[NV_NVDLA_CSC_dl.scala 983:120:@1376.4]
  wire  _T_2427; // @[NV_NVDLA_CSC_dl.scala 983:38:@1377.4]
  wire  _T_2428; // @[NV_NVDLA_CSC_dl.scala 984:50:@1378.4]
  wire  _T_2429; // @[NV_NVDLA_CSC_dl.scala 984:55:@1379.4]
  wire  _T_2430; // @[NV_NVDLA_CSC_dl.scala 984:73:@1380.4]
  wire  _T_2431; // @[NV_NVDLA_CSC_dl.scala 984:97:@1381.4]
  wire  _T_2434; // @[NV_NVDLA_CSC_dl.scala 984:120:@1383.4]
  wire  _T_2435; // @[NV_NVDLA_CSC_dl.scala 984:38:@1384.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_dl.scala 986:24:@1385.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_dl.scala 987:24:@1388.4]
  wire [7:0] _GEN_143; // @[NV_NVDLA_CSC_dl.scala 988:24:@1391.4]
  wire [7:0] _GEN_144; // @[NV_NVDLA_CSC_dl.scala 989:24:@1394.4]
  wire [7:0] _GEN_145; // @[NV_NVDLA_CSC_dl.scala 990:28:@1397.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl.scala 991:28:@1400.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl.scala 992:28:@1403.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl.scala 993:28:@1406.4]
  wire [7:0] _T_2436; // @[NV_NVDLA_CSC_dl.scala 1002:55:@1409.4]
  wire [63:0] _T_2439; // @[Cat.scala 30:58:@1412.4]
  wire [127:0] _T_2440; // @[Cat.scala 30:58:@1413.4]
  wire [255:0] _T_2441; // @[Cat.scala 30:58:@1414.4]
  wire [511:0] _T_2442; // @[Cat.scala 30:58:@1415.4]
  wire [511:0] _T_2443; // @[NV_NVDLA_CSC_dl.scala 1004:23:@1416.4]
  wire [511:0] _T_2447; // @[NV_NVDLA_CSC_dl.scala 1009:23:@1420.4]
  wire  _T_2453; // @[NV_NVDLA_CSC_dl.scala 1022:37:@1425.4]
  wire  _T_2456; // @[NV_NVDLA_CSC_dl.scala 1023:43:@1426.4]
  wire  _T_2457; // @[NV_NVDLA_CSC_dl.scala 1023:87:@1427.4]
  wire  _T_2459; // @[NV_NVDLA_CSC_dl.scala 1023:91:@1428.4]
  wire  _T_2460; // @[NV_NVDLA_CSC_dl.scala 1023:72:@1429.4]
  wire [255:0] _T_2462; // @[NV_NVDLA_CSC_dl.scala 1023:171:@1430.4]
  wire [511:0] _T_2463; // @[Cat.scala 30:58:@1431.4]
  wire  _T_2469; // @[NV_NVDLA_CSC_dl.scala 1024:72:@1435.4]
  wire [255:0] _T_2471; // @[NV_NVDLA_CSC_dl.scala 1024:171:@1436.4]
  wire [511:0] _T_2472; // @[Cat.scala 30:58:@1437.4]
  wire [511:0] _T_2473; // @[NV_NVDLA_CSC_dl.scala 1024:27:@1438.4]
  wire [511:0] _T_2474; // @[NV_NVDLA_CSC_dl.scala 1023:27:@1439.4]
  wire [511:0] _T_2475; // @[NV_NVDLA_CSC_dl.scala 1022:27:@1440.4]
  wire [7:0] _T_2546; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1443.4]
  wire [7:0] _T_2547; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1445.4]
  wire [7:0] _T_2548; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1447.4]
  wire [7:0] _T_2549; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1449.4]
  wire [7:0] _T_2550; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1451.4]
  wire [7:0] _T_2551; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1453.4]
  wire [7:0] _T_2552; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1455.4]
  wire [7:0] _T_2553; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1457.4]
  wire [7:0] _T_2554; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1459.4]
  wire [7:0] _T_2555; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1461.4]
  wire [7:0] _T_2556; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1463.4]
  wire [7:0] _T_2557; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1465.4]
  wire [7:0] _T_2558; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1467.4]
  wire [7:0] _T_2559; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1469.4]
  wire [7:0] _T_2560; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1471.4]
  wire [7:0] _T_2561; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1473.4]
  wire [7:0] _T_2562; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1475.4]
  wire [7:0] _T_2563; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1477.4]
  wire [7:0] _T_2564; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1479.4]
  wire [7:0] _T_2565; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1481.4]
  wire [7:0] _T_2566; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1483.4]
  wire [7:0] _T_2567; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1485.4]
  wire [7:0] _T_2568; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1487.4]
  wire [7:0] _T_2569; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1489.4]
  wire [7:0] _T_2570; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1491.4]
  wire [7:0] _T_2571; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1493.4]
  wire [7:0] _T_2572; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1495.4]
  wire [7:0] _T_2573; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1497.4]
  wire [7:0] _T_2574; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1499.4]
  wire [7:0] _T_2575; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1501.4]
  wire [7:0] _T_2576; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1503.4]
  wire [7:0] _T_2577; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1505.4]
  wire [7:0] _T_2578; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1507.4]
  wire [7:0] _T_2579; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1509.4]
  wire [7:0] _T_2580; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1511.4]
  wire [7:0] _T_2581; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1513.4]
  wire [7:0] _T_2582; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1515.4]
  wire [7:0] _T_2583; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1517.4]
  wire [7:0] _T_2584; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1519.4]
  wire [7:0] _T_2585; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1521.4]
  wire [7:0] _T_2586; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1523.4]
  wire [7:0] _T_2587; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1525.4]
  wire [7:0] _T_2588; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1527.4]
  wire [7:0] _T_2589; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1529.4]
  wire [7:0] _T_2590; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1531.4]
  wire [7:0] _T_2591; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1533.4]
  wire [7:0] _T_2592; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1535.4]
  wire [7:0] _T_2593; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1537.4]
  wire [7:0] _T_2594; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1539.4]
  wire [7:0] _T_2595; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1541.4]
  wire [7:0] _T_2596; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1543.4]
  wire [7:0] _T_2597; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1545.4]
  wire [7:0] _T_2598; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1547.4]
  wire [7:0] _T_2599; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1549.4]
  wire [7:0] _T_2600; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1551.4]
  wire [7:0] _T_2601; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1553.4]
  wire [7:0] _T_2602; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1555.4]
  wire [7:0] _T_2603; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1557.4]
  wire [7:0] _T_2604; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1559.4]
  wire [7:0] _T_2605; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1561.4]
  wire [7:0] _T_2606; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1563.4]
  wire [7:0] _T_2607; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1565.4]
  wire [7:0] _T_2608; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1567.4]
  wire [7:0] _T_2609; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1569.4]
  reg [255:0] _T_2611; // @[NV_NVDLA_CSC_dl.scala 1044:28:@1571.4]
  reg [255:0] _RAND_147;
  reg [127:0] _T_2613; // @[NV_NVDLA_CSC_dl.scala 1045:28:@1572.4]
  reg [127:0] _RAND_148;
  reg [127:0] _T_2615; // @[NV_NVDLA_CSC_dl.scala 1046:28:@1573.4]
  reg [127:0] _RAND_149;
  reg [127:0] _T_2617; // @[NV_NVDLA_CSC_dl.scala 1048:28:@1574.4]
  reg [127:0] _RAND_150;
  reg [127:0] _T_2619; // @[NV_NVDLA_CSC_dl.scala 1049:28:@1575.4]
  reg [127:0] _RAND_151;
  reg [127:0] _T_2621; // @[NV_NVDLA_CSC_dl.scala 1051:28:@1576.4]
  reg [127:0] _RAND_152;
  wire  _T_2622; // @[NV_NVDLA_CSC_dl.scala 1053:39:@1577.4]
  wire  _T_2623; // @[NV_NVDLA_CSC_dl.scala 1053:29:@1578.4]
  wire [1023:0] _T_2625; // @[Cat.scala 30:58:@1579.4]
  wire [1023:0] _T_2626; // @[NV_NVDLA_CSC_dl.scala 1053:28:@1580.4]
  wire  _T_2627; // @[NV_NVDLA_CSC_dl.scala 1054:39:@1581.4]
  wire  _T_2628; // @[NV_NVDLA_CSC_dl.scala 1054:29:@1582.4]
  wire [1023:0] _T_2630; // @[Cat.scala 30:58:@1583.4]
  wire [1023:0] _T_2631; // @[NV_NVDLA_CSC_dl.scala 1054:28:@1584.4]
  wire  _T_2632; // @[NV_NVDLA_CSC_dl.scala 1055:39:@1585.4]
  wire  _T_2633; // @[NV_NVDLA_CSC_dl.scala 1055:29:@1586.4]
  wire [1023:0] _T_2636; // @[NV_NVDLA_CSC_dl.scala 1055:28:@1588.4]
  wire  _T_2637; // @[NV_NVDLA_CSC_dl.scala 1056:39:@1589.4]
  wire  _T_2638; // @[NV_NVDLA_CSC_dl.scala 1056:29:@1590.4]
  wire [1023:0] _T_2641; // @[NV_NVDLA_CSC_dl.scala 1056:28:@1592.4]
  wire [10:0] _T_2643; // @[Cat.scala 30:58:@1593.4]
  wire [1023:0] _T_2644; // @[NV_NVDLA_CSC_dl.scala 1058:41:@1594.4]
  wire [511:0] _T_2645; // @[NV_NVDLA_CSC_dl.scala 1058:82:@1595.4]
  wire [10:0] _T_2647; // @[Cat.scala 30:58:@1596.4]
  wire [1023:0] _T_2648; // @[NV_NVDLA_CSC_dl.scala 1059:41:@1597.4]
  wire [511:0] _T_2649; // @[NV_NVDLA_CSC_dl.scala 1059:82:@1598.4]
  wire [10:0] _T_2651; // @[Cat.scala 30:58:@1599.4]
  wire [1023:0] _T_2652; // @[NV_NVDLA_CSC_dl.scala 1060:41:@1600.4]
  wire [511:0] _T_2653; // @[NV_NVDLA_CSC_dl.scala 1060:82:@1601.4]
  wire [10:0] _T_2655; // @[Cat.scala 30:58:@1602.4]
  wire [1023:0] _T_2656; // @[NV_NVDLA_CSC_dl.scala 1061:41:@1603.4]
  wire [511:0] _T_2657; // @[NV_NVDLA_CSC_dl.scala 1061:82:@1604.4]
  wire  _T_2658; // @[NV_NVDLA_CSC_dl.scala 1063:36:@1605.4]
  wire  _T_2659; // @[NV_NVDLA_CSC_dl.scala 1063:26:@1606.4]
  wire  _T_2662; // @[NV_NVDLA_CSC_dl.scala 1064:41:@1607.4]
  wire [127:0] _T_2663; // @[NV_NVDLA_CSC_dl.scala 1064:81:@1608.4]
  wire [511:0] _T_2669; // @[Cat.scala 30:58:@1614.4]
  wire  _T_2671; // @[NV_NVDLA_CSC_dl.scala 1065:41:@1615.4]
  wire [255:0] _T_2672; // @[NV_NVDLA_CSC_dl.scala 1065:81:@1616.4]
  wire [511:0] _T_2674; // @[Cat.scala 30:58:@1618.4]
  wire [511:0] _T_2676; // @[NV_NVDLA_CSC_dl.scala 1065:25:@1620.4]
  wire [511:0] _T_2677; // @[NV_NVDLA_CSC_dl.scala 1064:25:@1621.4]
  wire [511:0] _T_2678; // @[NV_NVDLA_CSC_dl.scala 1063:25:@1622.4]
  wire [7:0] _T_2749; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1624.4]
  wire [7:0] _T_2750; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1626.4]
  wire [7:0] _T_2751; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1628.4]
  wire [7:0] _T_2752; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1630.4]
  wire [7:0] _T_2753; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1632.4]
  wire [7:0] _T_2754; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1634.4]
  wire [7:0] _T_2755; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1636.4]
  wire [7:0] _T_2756; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1638.4]
  wire [7:0] _T_2757; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1640.4]
  wire [7:0] _T_2758; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1642.4]
  wire [7:0] _T_2759; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1644.4]
  wire [7:0] _T_2760; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1646.4]
  wire [7:0] _T_2761; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1648.4]
  wire [7:0] _T_2762; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1650.4]
  wire [7:0] _T_2763; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1652.4]
  wire [7:0] _T_2764; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1654.4]
  wire [7:0] _T_2765; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1656.4]
  wire [7:0] _T_2766; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1658.4]
  wire [7:0] _T_2767; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1660.4]
  wire [7:0] _T_2768; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1662.4]
  wire [7:0] _T_2769; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1664.4]
  wire [7:0] _T_2770; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1666.4]
  wire [7:0] _T_2771; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1668.4]
  wire [7:0] _T_2772; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1670.4]
  wire [7:0] _T_2773; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1672.4]
  wire [7:0] _T_2774; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1674.4]
  wire [7:0] _T_2775; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1676.4]
  wire [7:0] _T_2776; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1678.4]
  wire [7:0] _T_2777; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1680.4]
  wire [7:0] _T_2778; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1682.4]
  wire [7:0] _T_2779; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1684.4]
  wire [7:0] _T_2780; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1686.4]
  wire [7:0] _T_2781; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1688.4]
  wire [7:0] _T_2782; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1690.4]
  wire [7:0] _T_2783; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1692.4]
  wire [7:0] _T_2784; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1694.4]
  wire [7:0] _T_2785; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1696.4]
  wire [7:0] _T_2786; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1698.4]
  wire [7:0] _T_2787; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1700.4]
  wire [7:0] _T_2788; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1702.4]
  wire [7:0] _T_2789; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1704.4]
  wire [7:0] _T_2790; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1706.4]
  wire [7:0] _T_2791; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1708.4]
  wire [7:0] _T_2792; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1710.4]
  wire [7:0] _T_2793; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1712.4]
  wire [7:0] _T_2794; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1714.4]
  wire [7:0] _T_2795; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1716.4]
  wire [7:0] _T_2796; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1718.4]
  wire [7:0] _T_2797; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1720.4]
  wire [7:0] _T_2798; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1722.4]
  wire [7:0] _T_2799; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1724.4]
  wire [7:0] _T_2800; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1726.4]
  wire [7:0] _T_2801; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1728.4]
  wire [7:0] _T_2802; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1730.4]
  wire [7:0] _T_2803; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1732.4]
  wire [7:0] _T_2804; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1734.4]
  wire [7:0] _T_2805; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1736.4]
  wire [7:0] _T_2806; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1738.4]
  wire [7:0] _T_2807; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1740.4]
  wire [7:0] _T_2808; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1742.4]
  wire [7:0] _T_2809; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1744.4]
  wire [7:0] _T_2810; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1746.4]
  wire [7:0] _T_2811; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1748.4]
  wire [7:0] _T_2812; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1750.4]
  wire  _T_2814; // @[NV_NVDLA_CSC_dl.scala 1074:59:@1752.4]
  wire  _T_2815; // @[NV_NVDLA_CSC_dl.scala 1074:41:@1753.4]
  wire  _T_2817; // @[NV_NVDLA_CSC_dl.scala 1075:59:@1754.4]
  wire  _T_2818; // @[NV_NVDLA_CSC_dl.scala 1075:41:@1755.4]
  wire  _T_2821; // @[NV_NVDLA_CSC_dl.scala 1076:41:@1757.4]
  wire [511:0] _GEN_149; // @[NV_NVDLA_CSC_dl.scala 1078:24:@1758.4]
  wire [255:0] _GEN_150; // @[NV_NVDLA_CSC_dl.scala 1081:24:@1761.4]
  wire [511:0] _GEN_151; // @[NV_NVDLA_CSC_dl.scala 1081:24:@1761.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl.scala 1085:24:@1765.4]
  wire [318:0] _T_2827; // @[NV_NVDLA_CSC_dl.scala 1094:56:@1771.4]
  wire [63:0] _T_2828; // @[NV_NVDLA_CSC_dl.scala 1094:73:@1772.4]
  wire [63:0] _T_2829; // @[NV_NVDLA_CSC_dl.scala 1094:24:@1773.4]
  wire  _T_2831; // @[NV_NVDLA_CSC_dl.scala 1096:51:@1774.4]
  wire [63:0] _T_2838; // @[NV_NVDLA_CSC_dl.scala 1096:32:@1776.4]
  wire  _T_2840; // @[NV_NVDLA_CSC_dl.scala 1097:51:@1777.4]
  wire [31:0] _T_2847; // @[NV_NVDLA_CSC_dl.scala 1097:32:@1779.4]
  wire  _T_2849; // @[NV_NVDLA_CSC_dl.scala 1098:51:@1780.4]
  wire [31:0] _T_2856; // @[NV_NVDLA_CSC_dl.scala 1098:32:@1782.4]
  wire [31:0] _T_2857; // @[NV_NVDLA_CSC_dl.scala 1100:57:@1783.4]
  wire [63:0] _T_2863; // @[Cat.scala 30:58:@1785.4]
  wire [15:0] _T_2864; // @[NV_NVDLA_CSC_dl.scala 1101:57:@1786.4]
  wire [15:0] _T_2865; // @[NV_NVDLA_CSC_dl.scala 1101:106:@1787.4]
  wire [15:0] _T_2866; // @[NV_NVDLA_CSC_dl.scala 1101:155:@1788.4]
  wire [63:0] _T_2874; // @[Cat.scala 30:58:@1792.4]
  wire  _T_2876; // @[NV_NVDLA_CSC_dl.scala 1103:43:@1793.4]
  wire [15:0] _T_2877; // @[NV_NVDLA_CSC_dl.scala 1103:89:@1794.4]
  wire [63:0] _T_2879; // @[Cat.scala 30:58:@1796.4]
  wire [63:0] _T_2880; // @[NV_NVDLA_CSC_dl.scala 1103:116:@1797.4]
  wire  _T_2882; // @[NV_NVDLA_CSC_dl.scala 1104:43:@1798.4]
  wire [31:0] _T_2883; // @[NV_NVDLA_CSC_dl.scala 1104:89:@1799.4]
  wire [63:0] _T_2884; // @[Cat.scala 30:58:@1800.4]
  wire [63:0] _T_2885; // @[NV_NVDLA_CSC_dl.scala 1104:116:@1801.4]
  wire [63:0] _T_2886; // @[NV_NVDLA_CSC_dl.scala 1104:26:@1802.4]
  wire [63:0] _T_2887; // @[NV_NVDLA_CSC_dl.scala 1103:26:@1803.4]
  wire  _T_2888; // @[NV_NVDLA_CSC_dl.scala 1108:35:@1804.4]
  wire [7:0] _T_2889_0; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_1; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_2; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_3; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_4; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_5; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_6; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_7; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_8; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_9; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_10; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_11; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_12; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_13; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_14; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_15; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_16; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_17; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_18; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_19; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_20; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_21; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_22; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_23; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_24; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_25; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_26; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_27; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_28; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_29; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_30; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_31; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_32; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_33; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_34; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_35; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_36; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_37; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_38; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_39; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_40; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_41; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_42; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_43; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_44; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_45; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_46; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_47; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_48; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_49; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_50; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_51; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_52; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_53; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_54; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_55; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_56; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_57; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_58; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_59; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_60; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_61; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_62; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire [7:0] _T_2889_63; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  wire  _T_3022; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1806.4]
  wire  _T_3024; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1807.4]
  wire  _T_3026; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1808.4]
  wire  _T_3028; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1809.4]
  wire  _T_3030; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1810.4]
  wire  _T_3032; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1811.4]
  wire  _T_3034; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1812.4]
  wire  _T_3036; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1813.4]
  wire  _T_3038; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1814.4]
  wire  _T_3040; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1815.4]
  wire  _T_3042; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1816.4]
  wire  _T_3044; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1817.4]
  wire  _T_3046; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1818.4]
  wire  _T_3048; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1819.4]
  wire  _T_3050; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1820.4]
  wire  _T_3052; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1821.4]
  wire  _T_3054; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1822.4]
  wire  _T_3056; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1823.4]
  wire  _T_3058; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1824.4]
  wire  _T_3060; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1825.4]
  wire  _T_3062; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1826.4]
  wire  _T_3064; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1827.4]
  wire  _T_3066; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1828.4]
  wire  _T_3068; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1829.4]
  wire  _T_3070; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1830.4]
  wire  _T_3072; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1831.4]
  wire  _T_3074; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1832.4]
  wire  _T_3076; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1833.4]
  wire  _T_3078; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1834.4]
  wire  _T_3080; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1835.4]
  wire  _T_3082; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1836.4]
  wire  _T_3084; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1837.4]
  wire  _T_3086; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1838.4]
  wire  _T_3088; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1839.4]
  wire  _T_3090; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1840.4]
  wire  _T_3092; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1841.4]
  wire  _T_3094; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1842.4]
  wire  _T_3096; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1843.4]
  wire  _T_3098; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1844.4]
  wire  _T_3100; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1845.4]
  wire  _T_3102; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1846.4]
  wire  _T_3104; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1847.4]
  wire  _T_3106; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1848.4]
  wire  _T_3108; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1849.4]
  wire  _T_3110; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1850.4]
  wire  _T_3112; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1851.4]
  wire  _T_3114; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1852.4]
  wire  _T_3116; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1853.4]
  wire  _T_3118; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1854.4]
  wire  _T_3120; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1855.4]
  wire  _T_3122; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1856.4]
  wire  _T_3124; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1857.4]
  wire  _T_3126; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1858.4]
  wire  _T_3128; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1859.4]
  wire  _T_3130; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1860.4]
  wire  _T_3132; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1861.4]
  wire  _T_3134; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1862.4]
  wire  _T_3136; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1863.4]
  wire  _T_3138; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1864.4]
  wire  _T_3140; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1865.4]
  wire  _T_3142; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1866.4]
  wire  _T_3144; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1867.4]
  wire  _T_3146; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1868.4]
  wire  _T_3148; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1869.4]
  wire  _T_3219; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1935.4]
  wire  _T_3220; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1936.4]
  wire  _T_3221; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1937.4]
  wire  _T_3222; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1938.4]
  wire  _T_3223; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1939.4]
  wire  _T_3224; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1940.4]
  wire  _T_3225; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1941.4]
  wire  _T_3226; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1942.4]
  wire  _T_3227; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1943.4]
  wire  _T_3228; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1944.4]
  wire  _T_3229; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1945.4]
  wire  _T_3230; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1946.4]
  wire  _T_3231; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1947.4]
  wire  _T_3232; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1948.4]
  wire  _T_3233; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1949.4]
  wire  _T_3234; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1950.4]
  wire  _T_3235; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1951.4]
  wire  _T_3236; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1952.4]
  wire  _T_3237; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1953.4]
  wire  _T_3238; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1954.4]
  wire  _T_3239; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1955.4]
  wire  _T_3240; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1956.4]
  wire  _T_3241; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1957.4]
  wire  _T_3242; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1958.4]
  wire  _T_3243; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1959.4]
  wire  _T_3244; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1960.4]
  wire  _T_3245; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1961.4]
  wire  _T_3246; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1962.4]
  wire  _T_3247; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1963.4]
  wire  _T_3248; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1964.4]
  wire  _T_3249; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1965.4]
  wire  _T_3250; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1966.4]
  wire  _T_3251; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1967.4]
  wire  _T_3252; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1968.4]
  wire  _T_3253; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1969.4]
  wire  _T_3254; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1970.4]
  wire  _T_3255; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1971.4]
  wire  _T_3256; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1972.4]
  wire  _T_3257; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1973.4]
  wire  _T_3258; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1974.4]
  wire  _T_3259; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1975.4]
  wire  _T_3260; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1976.4]
  wire  _T_3261; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1977.4]
  wire  _T_3262; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1978.4]
  wire  _T_3263; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1979.4]
  wire  _T_3264; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1980.4]
  wire  _T_3265; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1981.4]
  wire  _T_3266; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1982.4]
  wire  _T_3267; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1983.4]
  wire  _T_3268; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1984.4]
  wire  _T_3269; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1985.4]
  wire  _T_3270; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1986.4]
  wire  _T_3271; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1987.4]
  wire  _T_3272; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1988.4]
  wire  _T_3273; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1989.4]
  wire  _T_3274; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1990.4]
  wire  _T_3275; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1991.4]
  wire  _T_3276; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1992.4]
  wire  _T_3277; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1993.4]
  wire  _T_3278; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1994.4]
  wire  _T_3279; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1995.4]
  wire  _T_3280; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1996.4]
  wire  _T_3281; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1997.4]
  wire  _T_3282; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1998.4]
  wire  _T_3283; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1999.4]
  wire  _T_3284; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2000.4]
  wire  _T_3285; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2001.4]
  wire  _T_3286; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2002.4]
  wire  _T_3287; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2003.4]
  wire  _T_3288; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2004.4]
  wire  _T_3289; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2005.4]
  wire  _T_3290; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2006.4]
  wire  _T_3291; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2007.4]
  wire  _T_3292; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2008.4]
  wire  _T_3293; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2009.4]
  wire  _T_3294; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2010.4]
  wire  _T_3295; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2011.4]
  wire  _T_3296; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2012.4]
  wire  _T_3297; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2013.4]
  wire  _T_3298; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2014.4]
  wire  _T_3299; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2015.4]
  wire  _T_3300; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2016.4]
  wire  _T_3301; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2017.4]
  wire  _T_3302; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2018.4]
  wire  _T_3303; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2019.4]
  wire  _T_3304; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2020.4]
  wire  _T_3305; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2021.4]
  wire  _T_3306; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2022.4]
  wire  _T_3307; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2023.4]
  wire  _T_3308; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2024.4]
  wire  _T_3309; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2025.4]
  wire  _T_3310; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2026.4]
  wire  _T_3311; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2027.4]
  wire  _T_3312; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2028.4]
  wire  _T_3313; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2029.4]
  wire  _T_3314; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2030.4]
  wire  _T_3315; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2031.4]
  wire  _T_3316; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2032.4]
  wire  _T_3317; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2033.4]
  wire  _T_3318; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2034.4]
  wire  _T_3319; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2035.4]
  wire  _T_3320; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2036.4]
  wire  _T_3321; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2037.4]
  wire  _T_3322; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2038.4]
  wire  _T_3323; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2039.4]
  wire  _T_3324; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2040.4]
  wire  _T_3325; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2041.4]
  wire  _T_3326; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2042.4]
  wire  _T_3327; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2043.4]
  wire  _T_3328; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2044.4]
  wire  _T_3329; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2045.4]
  wire  _T_3330; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2046.4]
  wire  _T_3331; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2047.4]
  wire  _T_3332; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2048.4]
  wire  _T_3333; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2049.4]
  wire  _T_3334; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2050.4]
  wire  _T_3335; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2051.4]
  wire  _T_3336; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2052.4]
  wire  _T_3337; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2053.4]
  wire  _T_3338; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2054.4]
  wire  _T_3339; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2055.4]
  wire  _T_3340; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2056.4]
  wire  _T_3341; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2057.4]
  wire  _T_3342; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2058.4]
  wire  _T_3343; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2059.4]
  wire  _T_3344; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2060.4]
  wire  _T_3345; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2061.4]
  wire  _T_3346; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2062.4]
  reg  _T_3419; // @[NV_NVDLA_CSC_dl.scala 1117:27:@2128.4]
  reg [31:0] _RAND_153;
  reg  _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_154;
  reg  _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_155;
  reg  _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_156;
  reg  _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_157;
  reg  _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_158;
  reg  _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_159;
  reg  _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_160;
  reg  _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_161;
  reg  _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_162;
  reg  _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_163;
  reg  _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_164;
  reg  _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_165;
  reg  _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_166;
  reg  _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_167;
  reg  _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_168;
  reg  _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_169;
  reg  _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_170;
  reg  _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_171;
  reg  _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_172;
  reg  _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_173;
  reg  _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_174;
  reg  _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_175;
  reg  _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_176;
  reg  _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_177;
  reg  _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_178;
  reg  _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_179;
  reg  _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_180;
  reg  _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_181;
  reg  _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_182;
  reg  _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_183;
  reg  _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_184;
  reg  _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_185;
  reg  _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_186;
  reg  _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_187;
  reg  _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_188;
  reg  _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_189;
  reg  _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_190;
  reg  _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_191;
  reg  _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_192;
  reg  _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_193;
  reg  _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_194;
  reg  _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_195;
  reg  _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_196;
  reg  _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_197;
  reg  _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_198;
  reg  _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_199;
  reg  _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_200;
  reg  _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_201;
  reg  _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_202;
  reg  _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_203;
  reg  _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_204;
  reg  _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_205;
  reg  _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_206;
  reg  _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_207;
  reg  _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_208;
  reg  _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_209;
  reg  _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_210;
  reg  _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_211;
  reg  _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_212;
  reg  _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_213;
  reg  _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_214;
  reg  _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_215;
  reg  _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_216;
  reg  _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1119:34:@2195.4]
  reg [31:0] _RAND_217;
  reg [7:0] _T_3889_0; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_218;
  reg [7:0] _T_3889_1; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_219;
  reg [7:0] _T_3889_2; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_220;
  reg [7:0] _T_3889_3; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_221;
  reg [7:0] _T_3889_4; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_222;
  reg [7:0] _T_3889_5; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_3889_6; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_224;
  reg [7:0] _T_3889_7; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_225;
  reg [7:0] _T_3889_8; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_226;
  reg [7:0] _T_3889_9; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_227;
  reg [7:0] _T_3889_10; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_228;
  reg [7:0] _T_3889_11; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_229;
  reg [7:0] _T_3889_12; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_230;
  reg [7:0] _T_3889_13; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_231;
  reg [7:0] _T_3889_14; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_232;
  reg [7:0] _T_3889_15; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_233;
  reg [7:0] _T_3889_16; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_234;
  reg [7:0] _T_3889_17; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_235;
  reg [7:0] _T_3889_18; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_236;
  reg [7:0] _T_3889_19; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_237;
  reg [7:0] _T_3889_20; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_238;
  reg [7:0] _T_3889_21; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_239;
  reg [7:0] _T_3889_22; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_240;
  reg [7:0] _T_3889_23; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_241;
  reg [7:0] _T_3889_24; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_242;
  reg [7:0] _T_3889_25; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_243;
  reg [7:0] _T_3889_26; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_244;
  reg [7:0] _T_3889_27; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_245;
  reg [7:0] _T_3889_28; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_246;
  reg [7:0] _T_3889_29; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_247;
  reg [7:0] _T_3889_30; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_248;
  reg [7:0] _T_3889_31; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_249;
  reg [7:0] _T_3889_32; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_250;
  reg [7:0] _T_3889_33; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_251;
  reg [7:0] _T_3889_34; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_252;
  reg [7:0] _T_3889_35; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_253;
  reg [7:0] _T_3889_36; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_254;
  reg [7:0] _T_3889_37; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_255;
  reg [7:0] _T_3889_38; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_256;
  reg [7:0] _T_3889_39; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_3889_40; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_3889_41; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_3889_42; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_3889_43; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_3889_44; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_3889_45; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_3889_46; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_3889_47; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_3889_48; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_3889_49; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_3889_50; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_3889_51; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_3889_52; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_3889_53; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_3889_54; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_3889_55; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_3889_56; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_3889_57; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_3889_58; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_3889_59; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_3889_60; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_3889_61; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_3889_62; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_3889_63; // @[NV_NVDLA_CSC_dl.scala 1120:30:@2196.4]
  reg [31:0] _RAND_281;
  wire  _GEN_156; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  wire  _T_3956; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2267.4]
  wire  _T_3957; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2271.4]
  wire  _T_3958; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2275.4]
  wire  _T_3959; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2279.4]
  wire  _T_3960; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2283.4]
  wire  _T_3961; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2287.4]
  wire  _T_3962; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2291.4]
  wire  _T_3963; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2295.4]
  wire  _T_3964; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2299.4]
  wire  _T_3965; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2303.4]
  wire  _T_3966; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2307.4]
  wire  _T_3967; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2311.4]
  wire  _T_3968; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2315.4]
  wire  _T_3969; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2319.4]
  wire  _T_3970; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2323.4]
  wire  _T_3971; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2327.4]
  wire  _T_3972; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2331.4]
  wire  _T_3973; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2335.4]
  wire  _T_3974; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2339.4]
  wire  _T_3975; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2343.4]
  wire  _T_3976; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2347.4]
  wire  _T_3977; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2351.4]
  wire  _T_3978; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2355.4]
  wire  _T_3979; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2359.4]
  wire  _T_3980; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2363.4]
  wire  _T_3981; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2367.4]
  wire  _T_3982; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2371.4]
  wire  _T_3983; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2375.4]
  wire  _T_3984; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2379.4]
  wire  _T_3985; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2383.4]
  wire  _T_3986; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2387.4]
  wire  _T_3987; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2391.4]
  wire  _T_3988; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2395.4]
  wire  _T_3989; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2399.4]
  wire  _T_3990; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2403.4]
  wire  _T_3991; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2407.4]
  wire  _T_3992; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2411.4]
  wire  _T_3993; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2415.4]
  wire  _T_3994; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2419.4]
  wire  _T_3995; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2423.4]
  wire  _T_3996; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2427.4]
  wire  _T_3997; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2431.4]
  wire  _T_3998; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2435.4]
  wire  _T_3999; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2439.4]
  wire  _T_4000; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2443.4]
  wire  _T_4001; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2447.4]
  wire  _T_4002; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2451.4]
  wire  _T_4003; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2455.4]
  wire  _T_4004; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2459.4]
  wire  _T_4005; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2463.4]
  wire  _T_4006; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2467.4]
  wire  _T_4007; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2471.4]
  wire  _T_4008; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2475.4]
  wire  _T_4009; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2479.4]
  wire  _T_4010; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2483.4]
  wire  _T_4011; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2487.4]
  wire  _T_4012; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2491.4]
  wire  _T_4013; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2495.4]
  wire  _T_4014; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2499.4]
  wire  _T_4015; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2503.4]
  wire  _T_4016; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2507.4]
  wire  _T_4017; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2511.4]
  wire  _T_4018; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2515.4]
  wire  _T_4019; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2519.4]
  reg  _T_4022; // @[NV_NVDLA_CSC_dl.scala 1145:26:@2523.4]
  reg [31:0] _RAND_282;
  reg  _T_4289_0; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_283;
  reg  _T_4289_1; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_284;
  reg  _T_4289_2; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_285;
  reg  _T_4289_3; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_286;
  reg  _T_4289_4; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_287;
  reg  _T_4289_5; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_288;
  reg  _T_4289_6; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_289;
  reg  _T_4289_7; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_290;
  reg  _T_4289_8; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_291;
  reg  _T_4289_9; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_292;
  reg  _T_4289_10; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_293;
  reg  _T_4289_11; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_294;
  reg  _T_4289_12; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_295;
  reg  _T_4289_13; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_296;
  reg  _T_4289_14; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_297;
  reg  _T_4289_15; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_298;
  reg  _T_4289_16; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_299;
  reg  _T_4289_17; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_300;
  reg  _T_4289_18; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_301;
  reg  _T_4289_19; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_302;
  reg  _T_4289_20; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_303;
  reg  _T_4289_21; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_304;
  reg  _T_4289_22; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_305;
  reg  _T_4289_23; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_306;
  reg  _T_4289_24; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_307;
  reg  _T_4289_25; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_308;
  reg  _T_4289_26; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_309;
  reg  _T_4289_27; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_310;
  reg  _T_4289_28; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_311;
  reg  _T_4289_29; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_312;
  reg  _T_4289_30; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_313;
  reg  _T_4289_31; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_314;
  reg  _T_4289_32; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_315;
  reg  _T_4289_33; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_316;
  reg  _T_4289_34; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_317;
  reg  _T_4289_35; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_318;
  reg  _T_4289_36; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_319;
  reg  _T_4289_37; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_320;
  reg  _T_4289_38; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_321;
  reg  _T_4289_39; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_322;
  reg  _T_4289_40; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_323;
  reg  _T_4289_41; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_324;
  reg  _T_4289_42; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_325;
  reg  _T_4289_43; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_326;
  reg  _T_4289_44; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_327;
  reg  _T_4289_45; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_328;
  reg  _T_4289_46; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_329;
  reg  _T_4289_47; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_330;
  reg  _T_4289_48; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_331;
  reg  _T_4289_49; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_332;
  reg  _T_4289_50; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_333;
  reg  _T_4289_51; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_334;
  reg  _T_4289_52; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_335;
  reg  _T_4289_53; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_336;
  reg  _T_4289_54; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_337;
  reg  _T_4289_55; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_338;
  reg  _T_4289_56; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_339;
  reg  _T_4289_57; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_340;
  reg  _T_4289_58; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_341;
  reg  _T_4289_59; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_342;
  reg  _T_4289_60; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_343;
  reg  _T_4289_61; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_344;
  reg  _T_4289_62; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_345;
  reg  _T_4289_63; // @[NV_NVDLA_CSC_dl.scala 1146:26:@2589.4]
  reg [31:0] _RAND_346;
  reg [8:0] _T_4488; // @[NV_NVDLA_CSC_dl.scala 1147:26:@2590.4]
  reg [31:0] _RAND_347;
  reg [7:0] _T_4492_0; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_348;
  reg [7:0] _T_4492_1; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_349;
  reg [7:0] _T_4492_2; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_350;
  reg [7:0] _T_4492_3; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_351;
  reg [7:0] _T_4492_4; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_352;
  reg [7:0] _T_4492_5; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_353;
  reg [7:0] _T_4492_6; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_354;
  reg [7:0] _T_4492_7; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_355;
  reg [7:0] _T_4492_8; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_356;
  reg [7:0] _T_4492_9; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_357;
  reg [7:0] _T_4492_10; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_358;
  reg [7:0] _T_4492_11; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_359;
  reg [7:0] _T_4492_12; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_360;
  reg [7:0] _T_4492_13; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_361;
  reg [7:0] _T_4492_14; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_362;
  reg [7:0] _T_4492_15; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_363;
  reg [7:0] _T_4492_16; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_364;
  reg [7:0] _T_4492_17; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_365;
  reg [7:0] _T_4492_18; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_366;
  reg [7:0] _T_4492_19; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_367;
  reg [7:0] _T_4492_20; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_368;
  reg [7:0] _T_4492_21; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_369;
  reg [7:0] _T_4492_22; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_370;
  reg [7:0] _T_4492_23; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_371;
  reg [7:0] _T_4492_24; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_372;
  reg [7:0] _T_4492_25; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_373;
  reg [7:0] _T_4492_26; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_374;
  reg [7:0] _T_4492_27; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_375;
  reg [7:0] _T_4492_28; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_376;
  reg [7:0] _T_4492_29; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_377;
  reg [7:0] _T_4492_30; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_378;
  reg [7:0] _T_4492_31; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_379;
  reg [7:0] _T_4492_32; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_380;
  reg [7:0] _T_4492_33; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_381;
  reg [7:0] _T_4492_34; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_382;
  reg [7:0] _T_4492_35; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_383;
  reg [7:0] _T_4492_36; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_384;
  reg [7:0] _T_4492_37; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_385;
  reg [7:0] _T_4492_38; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_386;
  reg [7:0] _T_4492_39; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_387;
  reg [7:0] _T_4492_40; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_388;
  reg [7:0] _T_4492_41; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_389;
  reg [7:0] _T_4492_42; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4492_43; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4492_44; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4492_45; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4492_46; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4492_47; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4492_48; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4492_49; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4492_50; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4492_51; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4492_52; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4492_53; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4492_54; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4492_55; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4492_56; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4492_57; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4492_58; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4492_59; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4492_60; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4492_61; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4492_62; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4492_63; // @[NV_NVDLA_CSC_dl.scala 1148:22:@2591.4]
  reg [31:0] _RAND_411;
  wire  _T_4559; // @[NV_NVDLA_CSC_dl.scala 1151:24:@2592.4]
  wire  _T_4694_0; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_1; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_2; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_3; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_4; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_5; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_6; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_7; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_8; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_9; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_10; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_11; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_12; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_13; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_14; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_15; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_16; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_17; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_18; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_19; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_20; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_21; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_22; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_23; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_24; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_25; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_26; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_27; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_28; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_29; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_30; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_31; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_32; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_33; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_34; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_35; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_36; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_37; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_38; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_39; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_40; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_41; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_42; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_43; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_44; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_45; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_46; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_47; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_48; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_49; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_50; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_51; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_52; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_53; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_54; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_55; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_56; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_57; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_58; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_59; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_60; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_61; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_62; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4694_63; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  wire  _T_4826; // @[NV_NVDLA_CSC_dl.scala 1155:19:@2660.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_289; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  wire [8:0] _GEN_348; // @[NV_NVDLA_CSC_dl.scala 1158:19:@2727.4]
  reg  _T_4829; // @[NV_NVDLA_CSC_dl.scala 1171:29:@2922.4]
  reg [31:0] _RAND_412;
  wire  _T_4830; // @[NV_NVDLA_CSC_dl.scala 1172:27:@2924.4]
  wire [8:0] _T_4832; // @[NV_NVDLA_CSC_dl.scala 1172:26:@2925.4]
  reg  _T_4835; // @[NV_NVDLA_CSC_dl.scala 1174:33:@2926.4]
  reg [31:0] _RAND_413;
  reg  _T_4838; // @[NV_NVDLA_CSC_dl.scala 1175:33:@2929.4]
  reg [31:0] _RAND_414;
  wire  _T_4840; // @[NV_NVDLA_CSC_dl.scala 1176:85:@2932.4]
  reg [8:0] _T_4842; // @[Reg.scala 19:20:@2933.4]
  reg [31:0] _RAND_415;
  wire [8:0] _GEN_413; // @[Reg.scala 20:19:@2934.4]
  reg [8:0] _T_4846; // @[Reg.scala 19:20:@2939.4]
  reg [31:0] _RAND_416;
  wire [8:0] _GEN_414; // @[Reg.scala 20:19:@2940.4]
  reg  _T_5114_0; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_417;
  reg  _T_5114_1; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_418;
  reg  _T_5114_2; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_419;
  reg  _T_5114_3; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_420;
  reg  _T_5114_4; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_421;
  reg  _T_5114_5; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_422;
  reg  _T_5114_6; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_423;
  reg  _T_5114_7; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_424;
  reg  _T_5114_8; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_425;
  reg  _T_5114_9; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_426;
  reg  _T_5114_10; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_427;
  reg  _T_5114_11; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_428;
  reg  _T_5114_12; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_429;
  reg  _T_5114_13; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_430;
  reg  _T_5114_14; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_431;
  reg  _T_5114_15; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_432;
  reg  _T_5114_16; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_433;
  reg  _T_5114_17; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_434;
  reg  _T_5114_18; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_435;
  reg  _T_5114_19; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_436;
  reg  _T_5114_20; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_437;
  reg  _T_5114_21; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_438;
  reg  _T_5114_22; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_439;
  reg  _T_5114_23; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_440;
  reg  _T_5114_24; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_441;
  reg  _T_5114_25; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_442;
  reg  _T_5114_26; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_443;
  reg  _T_5114_27; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_444;
  reg  _T_5114_28; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_445;
  reg  _T_5114_29; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_446;
  reg  _T_5114_30; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_447;
  reg  _T_5114_31; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_448;
  reg  _T_5114_32; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_449;
  reg  _T_5114_33; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_450;
  reg  _T_5114_34; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_451;
  reg  _T_5114_35; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_452;
  reg  _T_5114_36; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_453;
  reg  _T_5114_37; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_454;
  reg  _T_5114_38; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_455;
  reg  _T_5114_39; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_456;
  reg  _T_5114_40; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_457;
  reg  _T_5114_41; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_458;
  reg  _T_5114_42; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_459;
  reg  _T_5114_43; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_460;
  reg  _T_5114_44; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_461;
  reg  _T_5114_45; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_462;
  reg  _T_5114_46; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_463;
  reg  _T_5114_47; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_464;
  reg  _T_5114_48; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_465;
  reg  _T_5114_49; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_466;
  reg  _T_5114_50; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_467;
  reg  _T_5114_51; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_468;
  reg  _T_5114_52; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_469;
  reg  _T_5114_53; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_470;
  reg  _T_5114_54; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_471;
  reg  _T_5114_55; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_472;
  reg  _T_5114_56; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_473;
  reg  _T_5114_57; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_474;
  reg  _T_5114_58; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_475;
  reg  _T_5114_59; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_476;
  reg  _T_5114_60; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_477;
  reg  _T_5114_61; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_478;
  reg  _T_5114_62; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_479;
  reg  _T_5114_63; // @[Reg.scala 19:20:@3010.4]
  reg [31:0] _RAND_480;
  wire  _GEN_415; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_416; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_417; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_418; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_419; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_420; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_421; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_422; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_423; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_424; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_425; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@3011.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@3011.4]
  reg  _T_5578_0; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_481;
  reg  _T_5578_1; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_482;
  reg  _T_5578_2; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_483;
  reg  _T_5578_3; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_484;
  reg  _T_5578_4; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_485;
  reg  _T_5578_5; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_486;
  reg  _T_5578_6; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_487;
  reg  _T_5578_7; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_488;
  reg  _T_5578_8; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_489;
  reg  _T_5578_9; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_490;
  reg  _T_5578_10; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_491;
  reg  _T_5578_11; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_492;
  reg  _T_5578_12; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_493;
  reg  _T_5578_13; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_494;
  reg  _T_5578_14; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_495;
  reg  _T_5578_15; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_496;
  reg  _T_5578_16; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_497;
  reg  _T_5578_17; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_498;
  reg  _T_5578_18; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_499;
  reg  _T_5578_19; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_500;
  reg  _T_5578_20; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_501;
  reg  _T_5578_21; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_502;
  reg  _T_5578_22; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_503;
  reg  _T_5578_23; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_504;
  reg  _T_5578_24; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_505;
  reg  _T_5578_25; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_506;
  reg  _T_5578_26; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_507;
  reg  _T_5578_27; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_508;
  reg  _T_5578_28; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_509;
  reg  _T_5578_29; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_510;
  reg  _T_5578_30; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_511;
  reg  _T_5578_31; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_512;
  reg  _T_5578_32; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_513;
  reg  _T_5578_33; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_514;
  reg  _T_5578_34; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_515;
  reg  _T_5578_35; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_516;
  reg  _T_5578_36; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_517;
  reg  _T_5578_37; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_518;
  reg  _T_5578_38; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_519;
  reg  _T_5578_39; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_520;
  reg  _T_5578_40; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_521;
  reg  _T_5578_41; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_522;
  reg  _T_5578_42; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_523;
  reg  _T_5578_43; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_524;
  reg  _T_5578_44; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_525;
  reg  _T_5578_45; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_526;
  reg  _T_5578_46; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_527;
  reg  _T_5578_47; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_528;
  reg  _T_5578_48; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_529;
  reg  _T_5578_49; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_530;
  reg  _T_5578_50; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_531;
  reg  _T_5578_51; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_532;
  reg  _T_5578_52; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_533;
  reg  _T_5578_53; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_534;
  reg  _T_5578_54; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_535;
  reg  _T_5578_55; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_536;
  reg  _T_5578_56; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_537;
  reg  _T_5578_57; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_538;
  reg  _T_5578_58; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_539;
  reg  _T_5578_59; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_540;
  reg  _T_5578_60; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_541;
  reg  _T_5578_61; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_542;
  reg  _T_5578_62; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_543;
  reg  _T_5578_63; // @[Reg.scala 19:20:@3207.4]
  reg [31:0] _RAND_544;
  wire  _GEN_479; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_489; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@3208.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@3208.4]
  reg [7:0] _T_5776; // @[Reg.scala 11:16:@3338.4]
  reg [31:0] _RAND_545;
  reg [7:0] _T_5778; // @[Reg.scala 11:16:@3343.4]
  reg [31:0] _RAND_546;
  reg [7:0] _T_5780; // @[Reg.scala 11:16:@3348.4]
  reg [31:0] _RAND_547;
  reg [7:0] _T_5782; // @[Reg.scala 11:16:@3353.4]
  reg [31:0] _RAND_548;
  reg [7:0] _T_5784; // @[Reg.scala 11:16:@3358.4]
  reg [31:0] _RAND_549;
  reg [7:0] _T_5786; // @[Reg.scala 11:16:@3363.4]
  reg [31:0] _RAND_550;
  reg [7:0] _T_5788; // @[Reg.scala 11:16:@3368.4]
  reg [31:0] _RAND_551;
  reg [7:0] _T_5790; // @[Reg.scala 11:16:@3373.4]
  reg [31:0] _RAND_552;
  reg [7:0] _T_5792; // @[Reg.scala 11:16:@3378.4]
  reg [31:0] _RAND_553;
  reg [7:0] _T_5794; // @[Reg.scala 11:16:@3383.4]
  reg [31:0] _RAND_554;
  reg [7:0] _T_5796; // @[Reg.scala 11:16:@3388.4]
  reg [31:0] _RAND_555;
  reg [7:0] _T_5798; // @[Reg.scala 11:16:@3393.4]
  reg [31:0] _RAND_556;
  reg [7:0] _T_5800; // @[Reg.scala 11:16:@3398.4]
  reg [31:0] _RAND_557;
  reg [7:0] _T_5802; // @[Reg.scala 11:16:@3403.4]
  reg [31:0] _RAND_558;
  reg [7:0] _T_5804; // @[Reg.scala 11:16:@3408.4]
  reg [31:0] _RAND_559;
  reg [7:0] _T_5806; // @[Reg.scala 11:16:@3413.4]
  reg [31:0] _RAND_560;
  reg [7:0] _T_5808; // @[Reg.scala 11:16:@3418.4]
  reg [31:0] _RAND_561;
  reg [7:0] _T_5810; // @[Reg.scala 11:16:@3423.4]
  reg [31:0] _RAND_562;
  reg [7:0] _T_5812; // @[Reg.scala 11:16:@3428.4]
  reg [31:0] _RAND_563;
  reg [7:0] _T_5814; // @[Reg.scala 11:16:@3433.4]
  reg [31:0] _RAND_564;
  reg [7:0] _T_5816; // @[Reg.scala 11:16:@3438.4]
  reg [31:0] _RAND_565;
  reg [7:0] _T_5818; // @[Reg.scala 11:16:@3443.4]
  reg [31:0] _RAND_566;
  reg [7:0] _T_5820; // @[Reg.scala 11:16:@3448.4]
  reg [31:0] _RAND_567;
  reg [7:0] _T_5822; // @[Reg.scala 11:16:@3453.4]
  reg [31:0] _RAND_568;
  reg [7:0] _T_5824; // @[Reg.scala 11:16:@3458.4]
  reg [31:0] _RAND_569;
  reg [7:0] _T_5826; // @[Reg.scala 11:16:@3463.4]
  reg [31:0] _RAND_570;
  reg [7:0] _T_5828; // @[Reg.scala 11:16:@3468.4]
  reg [31:0] _RAND_571;
  reg [7:0] _T_5830; // @[Reg.scala 11:16:@3473.4]
  reg [31:0] _RAND_572;
  reg [7:0] _T_5832; // @[Reg.scala 11:16:@3478.4]
  reg [31:0] _RAND_573;
  reg [7:0] _T_5834; // @[Reg.scala 11:16:@3483.4]
  reg [31:0] _RAND_574;
  reg [7:0] _T_5836; // @[Reg.scala 11:16:@3488.4]
  reg [31:0] _RAND_575;
  reg [7:0] _T_5838; // @[Reg.scala 11:16:@3493.4]
  reg [31:0] _RAND_576;
  reg [7:0] _T_5840; // @[Reg.scala 11:16:@3498.4]
  reg [31:0] _RAND_577;
  reg [7:0] _T_5842; // @[Reg.scala 11:16:@3503.4]
  reg [31:0] _RAND_578;
  reg [7:0] _T_5844; // @[Reg.scala 11:16:@3508.4]
  reg [31:0] _RAND_579;
  reg [7:0] _T_5846; // @[Reg.scala 11:16:@3513.4]
  reg [31:0] _RAND_580;
  reg [7:0] _T_5848; // @[Reg.scala 11:16:@3518.4]
  reg [31:0] _RAND_581;
  reg [7:0] _T_5850; // @[Reg.scala 11:16:@3523.4]
  reg [31:0] _RAND_582;
  reg [7:0] _T_5852; // @[Reg.scala 11:16:@3528.4]
  reg [31:0] _RAND_583;
  reg [7:0] _T_5854; // @[Reg.scala 11:16:@3533.4]
  reg [31:0] _RAND_584;
  reg [7:0] _T_5856; // @[Reg.scala 11:16:@3538.4]
  reg [31:0] _RAND_585;
  reg [7:0] _T_5858; // @[Reg.scala 11:16:@3543.4]
  reg [31:0] _RAND_586;
  reg [7:0] _T_5860; // @[Reg.scala 11:16:@3548.4]
  reg [31:0] _RAND_587;
  reg [7:0] _T_5862; // @[Reg.scala 11:16:@3553.4]
  reg [31:0] _RAND_588;
  reg [7:0] _T_5864; // @[Reg.scala 11:16:@3558.4]
  reg [31:0] _RAND_589;
  reg [7:0] _T_5866; // @[Reg.scala 11:16:@3563.4]
  reg [31:0] _RAND_590;
  reg [7:0] _T_5868; // @[Reg.scala 11:16:@3568.4]
  reg [31:0] _RAND_591;
  reg [7:0] _T_5870; // @[Reg.scala 11:16:@3573.4]
  reg [31:0] _RAND_592;
  reg [7:0] _T_5872; // @[Reg.scala 11:16:@3578.4]
  reg [31:0] _RAND_593;
  reg [7:0] _T_5874; // @[Reg.scala 11:16:@3583.4]
  reg [31:0] _RAND_594;
  reg [7:0] _T_5876; // @[Reg.scala 11:16:@3588.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5878; // @[Reg.scala 11:16:@3593.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5880; // @[Reg.scala 11:16:@3598.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5882; // @[Reg.scala 11:16:@3603.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5884; // @[Reg.scala 11:16:@3608.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5886; // @[Reg.scala 11:16:@3613.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5888; // @[Reg.scala 11:16:@3618.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5890; // @[Reg.scala 11:16:@3623.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5892; // @[Reg.scala 11:16:@3628.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5894; // @[Reg.scala 11:16:@3633.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5896; // @[Reg.scala 11:16:@3638.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5898; // @[Reg.scala 11:16:@3643.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5900; // @[Reg.scala 11:16:@3648.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5902; // @[Reg.scala 11:16:@3653.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5904; // @[Reg.scala 11:16:@3658.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5906; // @[Reg.scala 11:16:@3663.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5908; // @[Reg.scala 11:16:@3668.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5910; // @[Reg.scala 11:16:@3673.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5912; // @[Reg.scala 11:16:@3678.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5914; // @[Reg.scala 11:16:@3683.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5916; // @[Reg.scala 11:16:@3688.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5918; // @[Reg.scala 11:16:@3693.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5920; // @[Reg.scala 11:16:@3698.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5922; // @[Reg.scala 11:16:@3703.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5924; // @[Reg.scala 11:16:@3708.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5926; // @[Reg.scala 11:16:@3713.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5928; // @[Reg.scala 11:16:@3718.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5930; // @[Reg.scala 11:16:@3723.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5932; // @[Reg.scala 11:16:@3728.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5934; // @[Reg.scala 11:16:@3733.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5936; // @[Reg.scala 11:16:@3738.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5938; // @[Reg.scala 11:16:@3743.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5940; // @[Reg.scala 11:16:@3748.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5942; // @[Reg.scala 11:16:@3753.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5944; // @[Reg.scala 11:16:@3758.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5946; // @[Reg.scala 11:16:@3763.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5948; // @[Reg.scala 11:16:@3768.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5950; // @[Reg.scala 11:16:@3773.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5952; // @[Reg.scala 11:16:@3778.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5954; // @[Reg.scala 11:16:@3783.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5956; // @[Reg.scala 11:16:@3788.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5958; // @[Reg.scala 11:16:@3793.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5960; // @[Reg.scala 11:16:@3798.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5962; // @[Reg.scala 11:16:@3803.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5964; // @[Reg.scala 11:16:@3808.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5966; // @[Reg.scala 11:16:@3813.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5968; // @[Reg.scala 11:16:@3818.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5970; // @[Reg.scala 11:16:@3823.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5972; // @[Reg.scala 11:16:@3828.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5974; // @[Reg.scala 11:16:@3833.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5976; // @[Reg.scala 11:16:@3838.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5978; // @[Reg.scala 11:16:@3843.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5980; // @[Reg.scala 11:16:@3848.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5982; // @[Reg.scala 11:16:@3853.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5984; // @[Reg.scala 11:16:@3858.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5986; // @[Reg.scala 11:16:@3863.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5988; // @[Reg.scala 11:16:@3868.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5990; // @[Reg.scala 11:16:@3873.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5992; // @[Reg.scala 11:16:@3878.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5994; // @[Reg.scala 11:16:@3883.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5996; // @[Reg.scala 11:16:@3888.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_5998; // @[Reg.scala 11:16:@3893.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_6000; // @[Reg.scala 11:16:@3898.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_6002; // @[Reg.scala 11:16:@3903.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_6004; // @[Reg.scala 11:16:@3908.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_6006; // @[Reg.scala 11:16:@3913.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_6008; // @[Reg.scala 11:16:@3918.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_6010; // @[Reg.scala 11:16:@3923.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_6012; // @[Reg.scala 11:16:@3928.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_6014; // @[Reg.scala 11:16:@3933.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_6016; // @[Reg.scala 11:16:@3938.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_6018; // @[Reg.scala 11:16:@3943.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_6020; // @[Reg.scala 11:16:@3948.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_6022; // @[Reg.scala 11:16:@3953.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_6024; // @[Reg.scala 11:16:@3958.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_6026; // @[Reg.scala 11:16:@3963.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_6028; // @[Reg.scala 11:16:@3968.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_6030; // @[Reg.scala 11:16:@3973.4]
  reg [31:0] _RAND_672;
  assign _T_622 = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_dl.scala 75:31:@8.4]
  assign _T_626 = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_dl.scala 77:31:@10.4]
  assign _T_630 = io_reg2dp_op_en & _T_622; // @[NV_NVDLA_CSC_dl.scala 84:32:@13.4]
  assign _T_634 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl.scala 86:35:@15.4]
  assign _T_635 = _T_634 & io_reg2dp_datain_format; // @[NV_NVDLA_CSC_dl.scala 87:22:@16.4]
  assign _T_640 = 7'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_dl.scala 94:53:@17.4]
  assign _T_642 = _T_635 ? _T_640 : 7'h8; // @[NV_NVDLA_CSC_dl.scala 94:24:@18.4]
  assign _T_643 = _T_642[5:3]; // @[NV_NVDLA_CSC_dl.scala 94:100:@19.4]
  assign _T_645 = _T_635 ? _T_643 : 3'h1; // @[NV_NVDLA_CSC_dl.scala 95:22:@20.4]
  assign _T_647 = _T_645 - 3'h1; // @[NV_NVDLA_CSC_dl.scala 96:34:@21.4]
  assign _T_648 = $unsigned(_T_647); // @[NV_NVDLA_CSC_dl.scala 96:34:@22.4]
  assign _T_650 = io_reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl.scala 97:51:@23.4]
  assign _T_651 = io_reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl.scala 98:62:@24.4]
  assign _T_654 = {_T_650,2'h0}; // @[Cat.scala 30:58:@25.4]
  assign _T_657 = {_T_650,1'h0}; // @[Cat.scala 30:58:@26.4]
  assign _GEN_671 = {{1'd0}, _T_650}; // @[NV_NVDLA_CSC_dl.scala 100:74:@27.4]
  assign _T_658 = _T_657 + _GEN_671; // @[NV_NVDLA_CSC_dl.scala 100:74:@27.4]
  assign _T_659 = 2'h2 == _T_651; // @[Mux.scala 46:19:@28.4]
  assign _T_660 = _T_659 ? _T_658 : {{2'd0}, _T_650}; // @[Mux.scala 46:16:@29.4]
  assign _T_661 = 2'h3 == _T_651; // @[Mux.scala 46:19:@30.4]
  assign _T_662 = _T_661 ? _T_654 : _T_660; // @[Mux.scala 46:16:@31.4]
  assign _T_664 = io_reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl.scala 102:88:@32.4]
  assign _T_670 = io_reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl.scala 102:172:@34.4]
  assign _T_671 = _T_664 ? 6'h3f : _T_670; // @[NV_NVDLA_CSC_dl.scala 102:58:@35.4]
  assign _T_674 = {_T_662,1'h0}; // @[Cat.scala 30:58:@36.4]
  assign _GEN_672 = {{1'd0}, _T_662}; // @[NV_NVDLA_CSC_dl.scala 103:81:@37.4]
  assign _T_675 = _T_674 + _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@37.4]
  assign _T_676 = _T_674 + _GEN_672; // @[NV_NVDLA_CSC_dl.scala 103:81:@38.4]
  assign _GEN_673 = {{1'd0}, _T_670}; // @[NV_NVDLA_CSC_dl.scala 103:100:@40.4]
  assign _T_678 = _T_676 + _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@40.4]
  assign _T_679 = _T_676 + _GEN_673; // @[NV_NVDLA_CSC_dl.scala 103:100:@41.4]
  assign _T_682 = _T_662 + _T_670; // @[NV_NVDLA_CSC_dl.scala 104:58:@43.4]
  assign _T_683 = _T_662 + _T_670; // @[NV_NVDLA_CSC_dl.scala 104:58:@44.4]
  assign _T_684 = 2'h1 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@45.4]
  assign _T_685 = _T_684 ? _T_683 : _T_671; // @[Mux.scala 46:16:@46.4]
  assign _T_686 = 2'h2 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@47.4]
  assign _T_687 = _T_686 ? _T_679 : {{1'd0}, _T_685}; // @[Mux.scala 46:16:@48.4]
  assign _T_690 = _T_670 + 6'h1; // @[NV_NVDLA_CSC_dl.scala 105:80:@50.4]
  assign _T_693 = {_T_662,2'h0}; // @[Cat.scala 30:58:@51.4]
  assign _T_698 = _T_684 ? _T_674 : {{1'd0}, _T_662}; // @[Mux.scala 46:16:@54.4]
  assign _T_700 = _T_686 ? _T_693 : {{1'd0}, _T_698}; // @[Mux.scala 46:16:@56.4]
  assign _T_702 = {_T_662,6'h0}; // @[Cat.scala 30:58:@57.4]
  assign _T_704 = io_reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl.scala 115:52:@58.4]
  assign _T_707 = io_reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl.scala 116:60:@59.4]
  assign _T_708 = _T_635 ? 6'h1 : _T_707; // @[NV_NVDLA_CSC_dl.scala 116:21:@60.4]
  assign _T_711 = io_reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl.scala 117:60:@61.4]
  assign _T_712 = _T_635 ? 6'h1 : _T_711; // @[NV_NVDLA_CSC_dl.scala 117:21:@62.4]
  assign _T_794 = io_reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl.scala 133:43:@86.4]
  assign _T_796 = _T_794 * 15'h1; // @[NV_NVDLA_CSC_dl.scala 134:41:@88.4]
  assign _T_797 = _T_796[14:0]; // @[NV_NVDLA_CSC_dl.scala 134:56:@89.4]
  assign _T_798 = 6'h1 * _T_712; // @[NV_NVDLA_CSC_dl.scala 136:37:@90.4]
  assign _GEN_674 = {{9'd0}, _T_722}; // @[NV_NVDLA_CSC_dl.scala 137:34:@91.4]
  assign _T_799 = _T_743 * _GEN_674; // @[NV_NVDLA_CSC_dl.scala 137:34:@91.4]
  assign _T_800 = _T_799[11:0]; // @[NV_NVDLA_CSC_dl.scala 137:47:@92.4]
  assign _GEN_675 = {{1'd0}, _T_736}; // @[NV_NVDLA_CSC_dl.scala 138:34:@93.4]
  assign _T_801 = _T_743 * _GEN_675; // @[NV_NVDLA_CSC_dl.scala 138:34:@93.4]
  assign _T_802 = _T_801[11:0]; // @[NV_NVDLA_CSC_dl.scala 138:51:@94.4]
  assign _T_804 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl.scala 139:41:@95.4]
  assign _T_805 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl.scala 139:41:@96.4]
  assign _T_807 = io_reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl.scala 140:77:@97.4]
  assign _GEN_676 = {{1'd0}, io_reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl.scala 140:113:@98.4]
  assign _T_808 = io_reg2dp_datain_height_ext - _GEN_676; // @[NV_NVDLA_CSC_dl.scala 140:113:@98.4]
  assign _T_809 = $unsigned(_T_808); // @[NV_NVDLA_CSC_dl.scala 140:113:@99.4]
  assign _T_810 = io_reg2dp_skip_data_rls ? _T_807 : _T_809; // @[NV_NVDLA_CSC_dl.scala 140:23:@100.4]
  assign _T_811 = _T_715 ? _T_729 : _T_792; // @[NV_NVDLA_CSC_dl.scala 141:24:@101.4]
  assign _GEN_677 = {{1'd0}, _T_811}; // @[NV_NVDLA_CSC_dl.scala 142:38:@102.4]
  assign _T_812 = _T_750 * _GEN_677; // @[NV_NVDLA_CSC_dl.scala 142:38:@102.4]
  assign _T_813 = _T_812[14:0]; // @[NV_NVDLA_CSC_dl.scala 142:54:@103.4]
  assign _T_1038 = _T_635 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@174.6]
  assign _T_1040 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl.scala 191:38:@176.6]
  assign _T_1041 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl.scala 191:38:@177.6]
  assign _T_1043 = io_reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl.scala 192:48:@179.6]
  assign _T_1049 = io_reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl.scala 195:93:@184.6]
  assign _T_1050 = {4'h0,_T_1049}; // @[Cat.scala 30:58:@185.6]
  assign _T_1054 = {1'h0,io_reg2dp_entries}; // @[Cat.scala 30:58:@218.6]
  assign _GEN_1 = _T_630 ? _T_1038 : _T_831; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_2 = _T_630 ? _T_1041 : _T_838; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_3 = _T_630 ? _T_1043 : _T_845; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_4 = _T_630 ? io_reg2dp_datain_width_ext : _T_852; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_5 = _T_630 ? io_reg2dp_datain_height_ext : _T_859; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_6 = _T_630 ? _T_1050 : _T_866; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_7 = _T_630 ? _T_643 : _T_869; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_8 = _T_630 ? _T_643 : _T_872; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_10 = _T_630 ? _T_643 : _T_878; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_11 = _T_630 ? _T_643 : _T_881; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_12 = _T_630 ? _T_643 : _T_884; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_13 = _T_630 ? _T_643 : _T_887; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_15 = _T_630 ? _T_643 : _T_893; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_16 = _T_630 ? _T_643 : _T_896; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_18 = _T_630 ? _T_643 : _T_902; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_19 = _T_630 ? _T_645 : _T_905; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_20 = _T_630 ? _T_645 : _T_908; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_21 = _T_630 ? _T_650 : _T_915; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_22 = _T_630 ? _T_704 : _T_922; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_24 = _T_630 ? 6'h1 : _T_722; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_25 = _T_630 ? 5'h0 : _T_932; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_26 = _T_630 ? _T_687 : _T_939; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_27 = _T_630 ? _T_690 : _T_946; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_28 = _T_630 ? _T_700 : _T_953; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_29 = _T_630 ? {{1'd0}, _T_662} : _T_960; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_30 = _T_630 ? _T_702 : _T_967; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_31 = _T_630 ? _T_708 : _T_974; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_32 = _T_630 ? _T_712 : _T_981; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_33 = _T_630 ? io_reg2dp_pad_value : _T_988; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_34 = _T_630 ? _T_794 : _T_743; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_35 = _T_630 ? _T_797 : _T_750; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_36 = _T_630 ? _T_1054 : _T_995; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_37 = _T_630 ? {{2'd0}, _T_798} : _T_736; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_38 = _T_630 ? {{2'd0}, _T_805} : _T_729; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_39 = _T_630 ? _T_810 : _T_792; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_40 = _T_630 ? io_reg2dp_dataout_width : _T_757; // @[NV_NVDLA_CSC_dl.scala 188:15:@170.4]
  assign _GEN_43 = _T_715 ? _T_800 : _T_778; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  assign _GEN_44 = _T_715 ? _T_802 : _T_785; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  assign _GEN_45 = _T_715 ? _T_743 : _T_1002; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  assign _GEN_46 = _T_715 ? _T_743 : _T_1009; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  assign _GEN_47 = _T_715 ? _T_813 : _T_771; // @[NV_NVDLA_CSC_dl.scala 233:18:@231.4]
  assign _GEN_48 = _T_626 ? _T_792 : _T_1016; // @[NV_NVDLA_CSC_dl.scala 240:17:@238.4]
  assign _GEN_49 = _T_626 ? _T_813 : _T_1023; // @[NV_NVDLA_CSC_dl.scala 240:17:@238.4]
  assign _T_1156 = _T_1016 != 14'h0; // @[NV_NVDLA_CSC_dl.scala 304:37:@313.4]
  assign _T_1157 = io_sg2dl_reuse_rls & _T_1156; // @[NV_NVDLA_CSC_dl.scala 304:23:@314.4]
  assign _T_2241 = _T_878[2]; // @[NV_NVDLA_CSC_dl.scala 894:32:@1228.4]
  assign _T_2242 = _T_2241 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 894:36:@1229.4]
  assign _T_2243 = _T_878[1]; // @[NV_NVDLA_CSC_dl.scala 895:35:@1230.4]
  assign _T_2244 = _T_2243 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 895:39:@1231.4]
  assign _T_2245 = _T_2242 | _T_2244; // @[NV_NVDLA_CSC_dl.scala 894:57:@1232.4]
  assign _T_2246 = _T_878[0]; // @[NV_NVDLA_CSC_dl.scala 896:35:@1233.4]
  assign _T_2247 = _T_2246 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 896:39:@1234.4]
  assign _T_2248 = _T_2245 | _T_2247; // @[NV_NVDLA_CSC_dl.scala 895:60:@1235.4]
  assign _T_2249 = _T_881[2]; // @[NV_NVDLA_CSC_dl.scala 903:42:@1237.4]
  assign _T_2253 = _T_2249 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1239.4]
  assign _T_2254 = _T_2253 & _T_2231; // @[NV_NVDLA_CSC_dl.scala 903:47:@1240.4]
  assign _T_2255 = _T_881[1]; // @[NV_NVDLA_CSC_dl.scala 904:42:@1241.4]
  assign _T_2259 = _T_2255 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1243.4]
  assign _T_2260 = _T_2259 & _T_2225; // @[NV_NVDLA_CSC_dl.scala 904:47:@1244.4]
  assign _T_2261 = _T_2254 | _T_2260; // @[NV_NVDLA_CSC_dl.scala 903:66:@1245.4]
  assign _T_2262 = _T_881[0]; // @[NV_NVDLA_CSC_dl.scala 905:42:@1246.4]
  assign _T_2266 = _T_2262 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1248.4]
  assign _T_2267 = _T_2266 & _T_2222; // @[NV_NVDLA_CSC_dl.scala 905:47:@1249.4]
  assign _T_2268 = _T_2261 | _T_2267; // @[NV_NVDLA_CSC_dl.scala 904:66:@1250.4]
  assign _T_2287 = _T_2268[17]; // @[NV_NVDLA_CSC_dl.scala 929:26:@1269.4]
  assign _T_1154 = _T_2248 & _T_2287; // @[NV_NVDLA_CSC_dl.scala 301:29:@312.4]
  assign _T_1159 = _T_729 != 14'h0; // @[NV_NVDLA_CSC_dl.scala 304:66:@315.4]
  assign _T_1160 = _T_1154 & _T_1159; // @[NV_NVDLA_CSC_dl.scala 304:53:@316.4]
  assign _T_1161 = _T_1157 | _T_1160; // @[NV_NVDLA_CSC_dl.scala 304:42:@317.4]
  assign _T_1162 = _T_1154 ? _T_729 : _T_1016; // @[NV_NVDLA_CSC_dl.scala 305:28:@319.4]
  assign _T_1163 = _T_1154 ? _T_771 : _T_1023; // @[NV_NVDLA_CSC_dl.scala 306:29:@321.4]
  assign _T_1094 = _T_1161 ? _T_1163 : 15'h0; // @[NV_NVDLA_CSC_dl.scala 273:28:@261.4]
  assign _T_1102 = _T_1076 + _T_1094; // @[NV_NVDLA_CSC_dl.scala 278:37:@268.4]
  assign _T_1103 = _T_1076 + _T_1094; // @[NV_NVDLA_CSC_dl.scala 278:37:@269.4]
  assign _T_1109 = {_T_838,9'h0}; // @[Cat.scala 30:58:@271.4]
  assign _GEN_678 = {{1'd0}, _T_1109}; // @[NV_NVDLA_CSC_dl.scala 279:46:@272.4]
  assign _T_1110 = _T_1103 - _GEN_678; // @[NV_NVDLA_CSC_dl.scala 279:46:@272.4]
  assign _T_1111 = $unsigned(_T_1110); // @[NV_NVDLA_CSC_dl.scala 279:46:@273.4]
  assign _T_1112 = _T_1111[14:0]; // @[NV_NVDLA_CSC_dl.scala 279:46:@274.4]
  assign _T_1119 = _T_1103 >= _GEN_678; // @[NV_NVDLA_CSC_dl.scala 280:45:@277.4]
  assign _T_1121 = _T_1119 ? _T_1112 : _T_1103; // @[NV_NVDLA_CSC_dl.scala 281:83:@278.4]
  assign _T_1122 = io_sc2cdma_dat_pending_req ? 15'h0 : _T_1121; // @[NV_NVDLA_CSC_dl.scala 281:25:@279.4]
  assign _T_1148 = _T_1161 | io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl.scala 292:13:@302.4]
  assign _GEN_52 = _T_1148 ? _T_1122 : _T_1076; // @[NV_NVDLA_CSC_dl.scala 292:25:@303.4]
  assign _GEN_54 = _T_1161 ? _T_1162 : _T_1169; // @[Reg.scala 20:19:@327.4]
  assign _GEN_55 = _T_1161 ? _T_1163 : _T_1172; // @[Reg.scala 20:19:@332.4]
  assign _T_1222 = {{30'd0}, _T_1189}; // @[NV_NVDLA_CSC_dl.scala 341:19:@375.4 NV_NVDLA_CSC_dl.scala 345:12:@381.4]
  assign _GEN_61 = _T_1189 ? _T_1222 : _T_1225; // @[NV_NVDLA_CSC_dl.scala 349:23:@383.4]
  assign _GEN_62 = _T_1211 ? _T_1225 : _T_1228; // @[NV_NVDLA_CSC_dl.scala 349:23:@387.4]
  assign _GEN_63 = _T_1214 ? _T_1228 : _T_1231; // @[NV_NVDLA_CSC_dl.scala 349:23:@391.4]
  assign _GEN_64 = _T_1217 ? _T_1231 : _T_1234; // @[NV_NVDLA_CSC_dl.scala 349:23:@395.4]
  assign _T_1235 = _T_869[2]; // @[NV_NVDLA_CSC_dl.scala 354:30:@398.4]
  assign _T_1236 = _T_1235 & _T_1211; // @[NV_NVDLA_CSC_dl.scala 354:34:@399.4]
  assign _T_1237 = _T_869[1]; // @[NV_NVDLA_CSC_dl.scala 355:30:@400.4]
  assign _T_1238 = _T_1237 & _T_1217; // @[NV_NVDLA_CSC_dl.scala 355:34:@401.4]
  assign _T_1239 = _T_1236 | _T_1238; // @[NV_NVDLA_CSC_dl.scala 354:50:@402.4]
  assign _T_1240 = _T_869[0]; // @[NV_NVDLA_CSC_dl.scala 356:30:@403.4]
  assign _T_1241 = _T_1240 & _T_1220; // @[NV_NVDLA_CSC_dl.scala 356:34:@404.4]
  assign _T_1242 = _T_1239 | _T_1241; // @[NV_NVDLA_CSC_dl.scala 355:50:@405.4]
  assign _T_1243 = _T_872[2]; // @[NV_NVDLA_CSC_dl.scala 358:37:@406.4]
  assign _T_1247 = _T_1243 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@408.4]
  assign _T_1248 = _T_1247 & _T_1225; // @[NV_NVDLA_CSC_dl.scala 358:42:@409.4]
  assign _T_1249 = _T_872[1]; // @[NV_NVDLA_CSC_dl.scala 359:37:@410.4]
  assign _T_1253 = _T_1249 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@412.4]
  assign _T_1254 = _T_1253 & _T_1231; // @[NV_NVDLA_CSC_dl.scala 359:42:@413.4]
  assign _T_1255 = _T_1248 | _T_1254; // @[NV_NVDLA_CSC_dl.scala 358:56:@414.4]
  assign _T_1256 = _T_872[0]; // @[NV_NVDLA_CSC_dl.scala 360:37:@415.4]
  assign _T_1260 = _T_1256 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@417.4]
  assign _T_1261 = _T_1260 & _T_1234; // @[NV_NVDLA_CSC_dl.scala 360:42:@418.4]
  assign _T_1262 = _T_1255 | _T_1261; // @[NV_NVDLA_CSC_dl.scala 359:56:@419.4]
  assign _T_1263 = _T_1262[4:0]; // @[NV_NVDLA_CSC_dl.scala 363:24:@420.4]
  assign _T_1264 = _T_1262[9:5]; // @[NV_NVDLA_CSC_dl.scala 364:24:@421.4]
  assign _T_1265 = _T_1262[16:10]; // @[NV_NVDLA_CSC_dl.scala 365:28:@422.4]
  assign _T_1266 = _T_1262[23:17]; // @[NV_NVDLA_CSC_dl.scala 366:29:@423.4]
  assign _T_1267 = _T_1262[25:24]; // @[NV_NVDLA_CSC_dl.scala 367:25:@424.4]
  assign _T_1268 = _T_1262[26]; // @[NV_NVDLA_CSC_dl.scala 368:25:@425.4]
  assign _T_1269 = _T_1262[27]; // @[NV_NVDLA_CSC_dl.scala 369:27:@426.4]
  assign _T_1270 = _T_1262[28]; // @[NV_NVDLA_CSC_dl.scala 370:25:@427.4]
  assign _T_1271 = _T_1262[29]; // @[NV_NVDLA_CSC_dl.scala 371:25:@428.4]
  assign _T_1272 = _T_1262[30]; // @[NV_NVDLA_CSC_dl.scala 372:27:@429.4]
  assign _T_1283 = _T_1279 + 5'h1; // @[NV_NVDLA_CSC_dl.scala 381:24:@433.4]
  assign _T_1284 = _T_1279 + 5'h1; // @[NV_NVDLA_CSC_dl.scala 381:24:@434.4]
  assign _T_1287 = _T_1279 == _T_932; // @[NV_NVDLA_CSC_dl.scala 383:27:@438.4]
  assign _T_1285 = _T_1287 ? 5'h0 : _T_1284; // @[NV_NVDLA_CSC_dl.scala 380:17:@435.4]
  assign _T_1286 = _T_630 ? 5'h0 : _T_1285; // @[NV_NVDLA_CSC_dl.scala 379:17:@436.4]
  assign _T_1294 = _T_1290 + 2'h1; // @[NV_NVDLA_CSC_dl.scala 389:31:@442.4]
  assign _T_1295 = _T_1290 + 2'h1; // @[NV_NVDLA_CSC_dl.scala 389:31:@443.4]
  assign _GEN_682 = {{1'd0}, _T_1295}; // @[NV_NVDLA_CSC_dl.scala 390:32:@444.4]
  assign _T_1296 = _GEN_682 == _T_905; // @[NV_NVDLA_CSC_dl.scala 390:32:@444.4]
  assign _T_1298 = io_reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl.scala 391:61:@446.4]
  assign _T_1346 = _T_1306 != 7'h0; // @[NV_NVDLA_CSC_dl.scala 424:37:@483.4]
  assign _T_1347 = ~ _T_1346; // @[NV_NVDLA_CSC_dl.scala 424:24:@484.4]
  assign _T_1349 = _T_1290 != 2'h0; // @[NV_NVDLA_CSC_dl.scala 424:56:@485.4]
  assign _T_1350 = ~ _T_1349; // @[NV_NVDLA_CSC_dl.scala 424:44:@486.4]
  assign _T_1351 = _T_1347 & _T_1350; // @[NV_NVDLA_CSC_dl.scala 424:42:@487.4]
  assign _T_1353 = _T_1279 != 5'h0; // @[NV_NVDLA_CSC_dl.scala 424:75:@488.4]
  assign _T_1354 = ~ _T_1353; // @[NV_NVDLA_CSC_dl.scala 424:63:@489.4]
  assign _T_1355 = _T_1351 & _T_1354; // @[NV_NVDLA_CSC_dl.scala 424:61:@490.4]
  assign _T_1357 = _T_1355 ? 1'h0 : _T_1335; // @[NV_NVDLA_CSC_dl.scala 424:22:@491.4]
  assign _T_1358 = _T_1242 ? 1'h1 : _T_1357; // @[NV_NVDLA_CSC_dl.scala 423:22:@492.4]
  assign _T_1299 = _T_1298 & _T_1358; // @[NV_NVDLA_CSC_dl.scala 391:66:@447.4]
  assign _T_1300 = _T_630 | _T_1299; // @[NV_NVDLA_CSC_dl.scala 391:33:@448.4]
  assign _T_1301 = _T_630 | _T_1296; // @[NV_NVDLA_CSC_dl.scala 393:31:@450.6]
  assign _T_1303 = _T_1301 ? 2'h0 : _T_1295; // @[NV_NVDLA_CSC_dl.scala 393:21:@451.6]
  assign _GEN_65 = _T_1300 ? _T_1303 : _T_1290; // @[NV_NVDLA_CSC_dl.scala 392:23:@449.4]
  assign _T_1312 = _T_1306 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 401:33:@457.4]
  assign _T_1313 = _T_1306 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 401:33:@458.4]
  assign _T_1314 = _T_1313 == _T_1266; // @[NV_NVDLA_CSC_dl.scala 402:51:@459.4]
  assign _T_1315 = _T_1287 & _T_1314; // @[NV_NVDLA_CSC_dl.scala 402:33:@460.4]
  assign _T_1316 = _T_1315 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 403:34:@462.4]
  assign _T_1317 = _T_1358 & _T_1287; // @[NV_NVDLA_CSC_dl.scala 404:52:@464.4]
  assign _T_1318 = _T_630 | _T_1317; // @[NV_NVDLA_CSC_dl.scala 404:34:@465.4]
  assign _T_1320 = ~ _T_1296; // @[NV_NVDLA_CSC_dl.scala 408:41:@467.6]
  assign _T_1321 = _T_1315 & _T_1320; // @[NV_NVDLA_CSC_dl.scala 408:39:@468.6]
  assign _T_1324 = _T_1316 ? 7'h0 : _T_1313; // @[NV_NVDLA_CSC_dl.scala 409:22:@469.6]
  assign _T_1325 = _T_1321 ? 7'h0 : _T_1324; // @[NV_NVDLA_CSC_dl.scala 408:22:@470.6]
  assign _T_1326 = _T_630 ? 7'h0 : _T_1325; // @[NV_NVDLA_CSC_dl.scala 407:22:@471.6]
  assign _GEN_66 = _T_1318 ? _T_1326 : _T_1306; // @[NV_NVDLA_CSC_dl.scala 406:24:@466.4]
  assign _T_1343 = _T_1242 | _T_1329; // @[NV_NVDLA_CSC_dl.scala 422:27:@481.4]
  assign _T_1338 = _T_1343 & _T_1315; // @[NV_NVDLA_CSC_dl.scala 419:49:@478.4]
  assign _T_1341 = _T_1242 ? 1'h1 : _T_1329; // @[NV_NVDLA_CSC_dl.scala 420:32:@479.4]
  assign _T_1342 = _T_1338 ? 1'h0 : _T_1341; // @[NV_NVDLA_CSC_dl.scala 419:33:@480.4]
  assign _T_1363 = {1'h0,_T_1265}; // @[Cat.scala 30:58:@498.4]
  assign _GEN_67 = _T_1358 ? _T_1363 : _T_1361; // @[NV_NVDLA_CSC_dl.scala 434:21:@499.4]
  assign _GEN_683 = {{10'd0}, _T_908}; // @[NV_NVDLA_CSC_dl.scala 444:39:@504.4]
  assign _T_1370 = _T_1366 + _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@504.4]
  assign _T_1371 = _T_1366 + _GEN_683; // @[NV_NVDLA_CSC_dl.scala 444:39:@505.4]
  assign _T_1372 = _T_1287 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 445:29:@506.4]
  assign _T_1373 = _T_1366 >= _T_757; // @[NV_NVDLA_CSC_dl.scala 445:61:@507.4]
  assign _T_1374 = _T_1372 & _T_1373; // @[NV_NVDLA_CSC_dl.scala 445:44:@508.4]
  assign _T_1377 = ~ _T_1269; // @[NV_NVDLA_CSC_dl.scala 448:43:@511.4]
  assign _T_1378 = _T_1316 & _T_1377; // @[NV_NVDLA_CSC_dl.scala 448:41:@512.4]
  assign _T_1379 = _T_1374 ? {{9'd0}, _T_648} : _T_1371; // @[NV_NVDLA_CSC_dl.scala 449:26:@513.4]
  assign _T_1380 = _T_1378 ? _T_1369 : _T_1379; // @[NV_NVDLA_CSC_dl.scala 448:26:@514.4]
  assign _T_1381 = _T_630 ? {{9'd0}, _T_648} : _T_1380; // @[NV_NVDLA_CSC_dl.scala 447:26:@515.4]
  assign _T_1383 = _T_1317 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 450:70:@517.4]
  assign _T_1384 = _T_630 | _T_1383; // @[NV_NVDLA_CSC_dl.scala 450:37:@518.4]
  assign _T_1385 = _T_1358 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 451:55:@519.4]
  assign _T_1386 = _T_1385 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 451:71:@520.4]
  assign _T_1387 = _T_630 | _T_1386; // @[NV_NVDLA_CSC_dl.scala 451:37:@521.4]
  assign _GEN_68 = _T_1384 ? _T_1381 : _T_1366; // @[NV_NVDLA_CSC_dl.scala 453:27:@522.4]
  assign _GEN_69 = _T_1387 ? _T_1381 : _T_1369; // @[NV_NVDLA_CSC_dl.scala 456:27:@525.4]
  assign _T_1391 = _T_1390 == _T_866; // @[NV_NVDLA_CSC_dl.scala 463:37:@529.4]
  assign _T_1393 = _T_1385 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 464:70:@531.4]
  assign _T_1394 = _T_630 | _T_1393; // @[NV_NVDLA_CSC_dl.scala 464:36:@532.4]
  assign _T_1398 = _T_1390 + 11'h1; // @[NV_NVDLA_CSC_dl.scala 469:34:@534.6]
  assign _T_1399 = _T_1390 + 11'h1; // @[NV_NVDLA_CSC_dl.scala 469:34:@535.6]
  assign _T_1400 = _T_1269 ? 11'h0 : _T_1399; // @[NV_NVDLA_CSC_dl.scala 468:24:@536.6]
  assign _T_1401 = _T_630 ? 11'h0 : _T_1400; // @[NV_NVDLA_CSC_dl.scala 467:24:@537.6]
  assign _GEN_70 = _T_1394 ? _T_1401 : _T_1390; // @[NV_NVDLA_CSC_dl.scala 466:26:@533.4]
  assign _GEN_684 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl.scala 484:41:@549.4]
  assign _T_1430 = 13'h0 - _GEN_684; // @[NV_NVDLA_CSC_dl.scala 484:41:@549.4]
  assign _T_1431 = $unsigned(_T_1430); // @[NV_NVDLA_CSC_dl.scala 484:41:@550.4]
  assign _T_1432 = _T_635 ? 14'h0 : _T_1431; // @[NV_NVDLA_CSC_dl.scala 483:26:@551.4]
  assign _GEN_685 = {{10'd0}, _T_915}; // @[NV_NVDLA_CSC_dl.scala 485:37:@552.4]
  assign _T_1433 = _T_1404 + _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@552.4]
  assign _T_1434 = _T_1404 + _GEN_685; // @[NV_NVDLA_CSC_dl.scala 485:37:@553.4]
  assign _T_1437 = _T_1374 ? _T_1432 : _T_1434; // @[NV_NVDLA_CSC_dl.scala 490:25:@556.4]
  assign _T_1438 = _T_1378 ? _T_1407 : _T_1437; // @[NV_NVDLA_CSC_dl.scala 489:25:@557.4]
  assign _T_1439 = _T_630 ? _T_1432 : _T_1438; // @[NV_NVDLA_CSC_dl.scala 488:25:@558.4]
  assign _GEN_686 = {{1'd0}, _T_1263}; // @[NV_NVDLA_CSC_dl.scala 492:35:@559.4]
  assign _T_1440 = _GEN_686 * _T_974; // @[NV_NVDLA_CSC_dl.scala 492:35:@559.4]
  assign _GEN_687 = {{3'd0}, _T_1440}; // @[NV_NVDLA_CSC_dl.scala 493:33:@560.4]
  assign _T_1441 = _T_1404 + _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@560.4]
  assign _T_1442 = _T_1404 + _GEN_687; // @[NV_NVDLA_CSC_dl.scala 493:33:@561.4]
  assign _T_1445 = _T_831[0]; // @[NV_NVDLA_CSC_dl.scala 494:96:@564.4]
  assign _T_1446 = ~ _T_1445; // @[NV_NVDLA_CSC_dl.scala 494:86:@565.4]
  assign _T_1447 = _T_1383 & _T_1446; // @[NV_NVDLA_CSC_dl.scala 494:84:@566.4]
  assign _T_1448 = _T_630 | _T_1447; // @[NV_NVDLA_CSC_dl.scala 494:36:@567.4]
  assign _T_1451 = _T_831[1]; // @[NV_NVDLA_CSC_dl.scala 495:99:@570.4]
  assign _T_1452 = ~ _T_1451; // @[NV_NVDLA_CSC_dl.scala 495:89:@571.4]
  assign _T_1453 = _T_1386 & _T_1452; // @[NV_NVDLA_CSC_dl.scala 495:87:@572.4]
  assign _T_1454 = _T_630 | _T_1453; // @[NV_NVDLA_CSC_dl.scala 495:36:@573.4]
  assign _T_1456 = _T_1296 ? _T_953 : 8'h0; // @[NV_NVDLA_CSC_dl.scala 498:26:@574.4]
  assign _T_1459 = _T_670 == 6'h0; // @[NV_NVDLA_CSC_dl.scala 500:79:@576.4]
  assign _T_1463 = _T_1049 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 501:74:@579.4]
  assign _T_1464 = _T_1049 + 7'h1; // @[NV_NVDLA_CSC_dl.scala 501:74:@580.4]
  assign _T_1465 = _T_1459 ? _T_1049 : _T_1464; // @[NV_NVDLA_CSC_dl.scala 500:27:@581.4]
  assign _T_1466 = _T_1269 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 502:37:@582.4]
  assign _T_1468 = _T_1268 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 503:35:@583.4]
  assign _T_1470 = _T_1419 + 13'h1; // @[NV_NVDLA_CSC_dl.scala 503:66:@584.4]
  assign _T_1471 = _T_1419 + 13'h1; // @[NV_NVDLA_CSC_dl.scala 503:66:@585.4]
  assign _T_1472 = _T_1468 ? _T_1471 : _T_1419; // @[NV_NVDLA_CSC_dl.scala 503:22:@586.4]
  assign _T_1473 = _T_1466 ? 13'h2 : _T_1472; // @[NV_NVDLA_CSC_dl.scala 502:22:@587.4]
  assign _GEN_688 = {{6'd0}, _T_1465}; // @[NV_NVDLA_CSC_dl.scala 505:44:@589.4]
  assign _T_1474 = _T_1419 >= _GEN_688; // @[NV_NVDLA_CSC_dl.scala 505:44:@589.4]
  assign _T_1475 = _T_1316 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 509:39:@590.4]
  assign _T_1476 = _T_1475 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 509:54:@591.4]
  assign _T_1477 = _T_1476 & _T_1374; // @[NV_NVDLA_CSC_dl.scala 509:71:@592.4]
  assign _T_1480 = ~ _T_1374; // @[NV_NVDLA_CSC_dl.scala 510:73:@595.4]
  assign _T_1481 = _T_1476 & _T_1480; // @[NV_NVDLA_CSC_dl.scala 510:71:@596.4]
  assign _GEN_689 = {{4'd0}, _T_967}; // @[NV_NVDLA_CSC_dl.scala 510:99:@597.4]
  assign _T_1482 = _T_1416 + _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@597.4]
  assign _T_1483 = _T_1416 + _GEN_689; // @[NV_NVDLA_CSC_dl.scala 510:99:@598.4]
  assign _T_1485 = _T_1475 & _T_1474; // @[NV_NVDLA_CSC_dl.scala 511:54:@600.4]
  assign _GEN_690 = {{9'd0}, _T_946}; // @[NV_NVDLA_CSC_dl.scala 511:90:@601.4]
  assign _T_1486 = _T_1413 + _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@601.4]
  assign _T_1487 = _T_1413 + _GEN_690; // @[NV_NVDLA_CSC_dl.scala 511:90:@602.4]
  assign _T_1489 = ~ _T_1474; // @[NV_NVDLA_CSC_dl.scala 512:56:@604.4]
  assign _T_1490 = _T_1475 & _T_1489; // @[NV_NVDLA_CSC_dl.scala 512:54:@605.4]
  assign _T_1492 = _T_1413 + 16'h40; // @[NV_NVDLA_CSC_dl.scala 512:91:@606.4]
  assign _T_1493 = _T_1413 + 16'h40; // @[NV_NVDLA_CSC_dl.scala 512:91:@607.4]
  assign _T_1494 = ~ _T_1268; // @[NV_NVDLA_CSC_dl.scala 513:41:@608.4]
  assign _T_1495 = _T_1316 & _T_1494; // @[NV_NVDLA_CSC_dl.scala 513:39:@609.4]
  assign _GEN_691 = {{8'd0}, _T_1456}; // @[NV_NVDLA_CSC_dl.scala 513:81:@610.4]
  assign _T_1496 = _T_1410 + _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@610.4]
  assign _T_1497 = _T_1410 + _GEN_691; // @[NV_NVDLA_CSC_dl.scala 513:81:@611.4]
  assign _T_1498 = _T_1495 ? _T_1413 : _T_1497; // @[NV_NVDLA_CSC_dl.scala 513:24:@612.4]
  assign _T_1499 = _T_1490 ? _T_1493 : _T_1498; // @[NV_NVDLA_CSC_dl.scala 512:24:@613.4]
  assign _T_1500 = _T_1485 ? _T_1487 : _T_1499; // @[NV_NVDLA_CSC_dl.scala 511:24:@614.4]
  assign _T_1501 = _T_1481 ? _T_1483 : _T_1500; // @[NV_NVDLA_CSC_dl.scala 510:24:@615.4]
  assign _T_1502 = _T_1477 ? {{9'd0}, _T_939} : _T_1501; // @[NV_NVDLA_CSC_dl.scala 509:24:@616.4]
  assign _T_1503 = _T_715 ? {{9'd0}, _T_939} : _T_1502; // @[NV_NVDLA_CSC_dl.scala 508:24:@617.4]
  assign _T_1509 = _T_1410[15:6]; // @[NV_NVDLA_CSC_dl.scala 515:68:@619.4]
  assign _T_1510 = {5'h0,_T_1509}; // @[Cat.scala 30:58:@620.4]
  assign _T_1521 = _T_831[4]; // @[NV_NVDLA_CSC_dl.scala 518:68:@631.4]
  assign _T_1522 = _T_1358 & _T_1521; // @[NV_NVDLA_CSC_dl.scala 518:57:@632.4]
  assign _T_1523 = _T_1522 & _T_1316; // @[NV_NVDLA_CSC_dl.scala 518:72:@633.4]
  assign _T_1524 = _T_1523 & _T_1268; // @[NV_NVDLA_CSC_dl.scala 518:88:@634.4]
  assign _T_1525 = _T_1524 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 518:103:@635.4]
  assign _T_1526 = _T_715 | _T_1525; // @[NV_NVDLA_CSC_dl.scala 518:39:@636.4]
  assign _T_1528 = _T_1445 & _T_1242; // @[NV_NVDLA_CSC_dl.scala 520:42:@638.4]
  assign _T_1531 = _T_1424 ? 1'h0 : _T_1427; // @[NV_NVDLA_CSC_dl.scala 520:74:@639.4]
  assign _T_1532 = _T_1528 ? 1'h1 : _T_1531; // @[NV_NVDLA_CSC_dl.scala 520:28:@640.4]
  assign _T_1534 = _T_1445 & _T_1296; // @[NV_NVDLA_CSC_dl.scala 521:36:@642.4]
  assign _T_1535 = _T_1532 | _T_1427; // @[NV_NVDLA_CSC_dl.scala 521:72:@643.4]
  assign _T_1536 = _T_1534 & _T_1535; // @[NV_NVDLA_CSC_dl.scala 521:51:@644.4]
  assign _GEN_71 = _T_1448 ? _T_1439 : _T_1404; // @[NV_NVDLA_CSC_dl.scala 523:26:@645.4]
  assign _GEN_72 = _T_1448 ? _T_1503 : _T_1410; // @[NV_NVDLA_CSC_dl.scala 523:26:@645.4]
  assign _GEN_73 = _T_1454 ? _T_1439 : _T_1407; // @[NV_NVDLA_CSC_dl.scala 527:26:@649.4]
  assign _GEN_74 = _T_1454 ? _T_1503 : _T_1413; // @[NV_NVDLA_CSC_dl.scala 527:26:@649.4]
  assign _GEN_75 = _T_1526 ? _T_1503 : _T_1416; // @[NV_NVDLA_CSC_dl.scala 531:26:@653.4]
  assign _GEN_692 = {{9'd0}, io_reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl.scala 540:41:@658.4]
  assign _T_1544 = 14'h0 - _GEN_692; // @[NV_NVDLA_CSC_dl.scala 540:41:@658.4]
  assign _T_1545 = $unsigned(_T_1544); // @[NV_NVDLA_CSC_dl.scala 540:41:@659.4]
  assign _T_1546 = _T_1545[13:0]; // @[NV_NVDLA_CSC_dl.scala 540:41:@660.4]
  assign _GEN_693 = {{10'd0}, _T_922}; // @[NV_NVDLA_CSC_dl.scala 541:37:@661.4]
  assign _T_1547 = _T_1539 + _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@661.4]
  assign _T_1548 = _T_1539 + _GEN_693; // @[NV_NVDLA_CSC_dl.scala 541:37:@662.4]
  assign _T_1549 = _T_1316 & _T_1270; // @[NV_NVDLA_CSC_dl.scala 542:52:@663.4]
  assign _T_1550 = _T_630 | _T_1549; // @[NV_NVDLA_CSC_dl.scala 542:35:@664.4]
  assign _T_1553 = _T_1374 ? _T_1548 : _T_1539; // @[NV_NVDLA_CSC_dl.scala 544:25:@667.4]
  assign _T_1554 = _T_1378 ? _T_1542 : _T_1553; // @[NV_NVDLA_CSC_dl.scala 543:25:@668.4]
  assign _T_1555 = _T_1550 ? _T_1546 : _T_1554; // @[NV_NVDLA_CSC_dl.scala 542:25:@669.4]
  assign _T_1558 = _T_1378 | _T_1374; // @[NV_NVDLA_CSC_dl.scala 545:91:@672.4]
  assign _T_1559 = _T_1358 & _T_1558; // @[NV_NVDLA_CSC_dl.scala 545:54:@673.4]
  assign _T_1560 = _T_630 | _T_1559; // @[NV_NVDLA_CSC_dl.scala 545:36:@674.4]
  assign _GEN_694 = {{1'd0}, _T_1264}; // @[NV_NVDLA_CSC_dl.scala 547:35:@678.4]
  assign _T_1564 = _GEN_694 * _T_981; // @[NV_NVDLA_CSC_dl.scala 547:35:@678.4]
  assign _GEN_695 = {{3'd0}, _T_1564}; // @[NV_NVDLA_CSC_dl.scala 548:33:@679.4]
  assign _T_1565 = _T_1539 + _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@679.4]
  assign _T_1566 = _T_1539 + _GEN_695; // @[NV_NVDLA_CSC_dl.scala 548:33:@680.4]
  assign _GEN_696 = {{12'd0}, _T_1290}; // @[NV_NVDLA_CSC_dl.scala 548:51:@681.4]
  assign _T_1567 = _T_1566 + _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@681.4]
  assign _T_1568 = _T_1566 + _GEN_696; // @[NV_NVDLA_CSC_dl.scala 548:51:@682.4]
  assign _GEN_76 = _T_1560 ? _T_1555 : _T_1539; // @[NV_NVDLA_CSC_dl.scala 550:26:@683.4]
  assign _GEN_77 = _T_1387 ? _T_1555 : _T_1542; // @[NV_NVDLA_CSC_dl.scala 551:26:@686.4]
  assign _T_1569 = _T_1442[13]; // @[NV_NVDLA_CSC_dl.scala 554:39:@689.4]
  assign _GEN_697 = {{1'd0}, _T_852}; // @[NV_NVDLA_CSC_dl.scala 554:59:@690.4]
  assign _T_1570 = _T_1442 > _GEN_697; // @[NV_NVDLA_CSC_dl.scala 554:59:@690.4]
  assign _T_1571 = _T_1569 | _T_1570; // @[NV_NVDLA_CSC_dl.scala 554:44:@691.4]
  assign _T_1572 = _T_1568[13]; // @[NV_NVDLA_CSC_dl.scala 554:92:@692.4]
  assign _T_1573 = _T_1571 | _T_1572; // @[NV_NVDLA_CSC_dl.scala 554:78:@693.4]
  assign _GEN_698 = {{1'd0}, _T_859}; // @[NV_NVDLA_CSC_dl.scala 554:112:@694.4]
  assign _T_1574 = _T_1568 > _GEN_698; // @[NV_NVDLA_CSC_dl.scala 554:112:@694.4]
  assign _T_1575 = _T_1573 | _T_1574; // @[NV_NVDLA_CSC_dl.scala 554:97:@695.4]
  assign _T_1588 = _T_1572 | _T_1574; // @[NV_NVDLA_CSC_dl.scala 557:42:@705.4]
  assign _T_1698 = _T_831[10]; // @[NV_NVDLA_CSC_dl.scala 642:33:@791.4]
  assign _T_1699 = ~ _T_1391; // @[NV_NVDLA_CSC_dl.scala 643:24:@792.4]
  assign _T_1701 = _T_1442[12:0]; // @[NV_NVDLA_CSC_dl.scala 643:77:@793.4]
  assign _T_1702 = {2'h0,_T_1701}; // @[Cat.scala 30:58:@794.4]
  assign _T_1704 = _T_1363 > 8'h20; // @[NV_NVDLA_CSC_dl.scala 644:38:@795.4]
  assign _T_1709 = _T_1442[12:1]; // @[NV_NVDLA_CSC_dl.scala 645:54:@798.4]
  assign _T_1710 = {3'h0,_T_1709}; // @[Cat.scala 30:58:@799.4]
  assign _T_1711 = _T_1704 ? _T_1702 : _T_1710; // @[NV_NVDLA_CSC_dl.scala 644:23:@800.4]
  assign _T_1712 = _T_1699 ? _T_1702 : _T_1711; // @[NV_NVDLA_CSC_dl.scala 643:23:@801.4]
  assign _T_1713 = _T_1698 ? _T_1510 : _T_1712; // @[NV_NVDLA_CSC_dl.scala 642:23:@802.4]
  assign _T_1714 = _T_1713[13:0]; // @[NV_NVDLA_CSC_dl.scala 654:24:@804.4]
  assign _T_1591 = _T_1714[13:2]; // @[NV_NVDLA_CSC_dl.scala 561:32:@707.4]
  assign _GEN_700 = {{3'd0}, _T_1591}; // @[NV_NVDLA_CSC_dl.scala 561:40:@708.4]
  assign _T_1592 = _GEN_700 > _T_995; // @[NV_NVDLA_CSC_dl.scala 561:40:@708.4]
  assign _T_1593 = _T_831[5]; // @[NV_NVDLA_CSC_dl.scala 562:34:@709.4]
  assign _T_1594 = _T_1593 ? _T_1588 : _T_1575; // @[NV_NVDLA_CSC_dl.scala 562:24:@710.4]
  assign _T_1595 = _T_831[6]; // @[NV_NVDLA_CSC_dl.scala 563:29:@711.4]
  assign _T_1596 = _T_1595 & _T_1592; // @[NV_NVDLA_CSC_dl.scala 563:33:@712.4]
  assign _T_1597 = ~ _T_1594; // @[NV_NVDLA_CSC_dl.scala 564:39:@713.4]
  assign _T_1598 = _T_1358 & _T_1597; // @[NV_NVDLA_CSC_dl.scala 564:37:@714.4]
  assign _T_1599 = ~ _T_1596; // @[NV_NVDLA_CSC_dl.scala 564:56:@715.4]
  assign _T_1600 = _T_1598 & _T_1599; // @[NV_NVDLA_CSC_dl.scala 564:54:@716.4]
  assign _T_1601 = _T_831[7]; // @[NV_NVDLA_CSC_dl.scala 567:37:@717.4]
  assign _T_1602 = ~ _T_1601; // @[NV_NVDLA_CSC_dl.scala 567:27:@718.4]
  assign _T_1603 = _T_1390[0]; // @[NV_NVDLA_CSC_dl.scala 567:54:@719.4]
  assign _T_1604 = _T_1602 ? _T_1603 : _T_1268; // @[NV_NVDLA_CSC_dl.scala 567:26:@720.4]
  assign _T_1605 = _T_1442[1:0]; // @[NV_NVDLA_CSC_dl.scala 568:35:@721.4]
  assign _T_1607 = _T_1290 == 2'h0; // @[NV_NVDLA_CSC_dl.scala 569:55:@722.4]
  assign _T_1608 = _T_1358 & _T_1607; // @[NV_NVDLA_CSC_dl.scala 569:42:@723.4]
  assign _T_1609 = _T_1315 & _T_1343; // @[NV_NVDLA_CSC_dl.scala 572:42:@725.4]
  assign _T_1613 = {_T_1271,_T_1269,_T_1609,_T_1242,_T_1279}; // @[Cat.scala 30:58:@729.4]
  assign _T_1644 = _T_1272 & _T_1315; // @[NV_NVDLA_CSC_dl.scala 599:38:@749.6]
  assign _T_1645 = _T_1644 & _T_1343; // @[NV_NVDLA_CSC_dl.scala 599:56:@750.6]
  assign _GEN_78 = _T_1358 ? _T_1605 : _T_1619; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_79 = _T_1358 ? _T_1290 : _T_1622; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_80 = _T_1358 ? _T_1604 : _T_1625; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_81 = _T_1358 ? _T_1391 : _T_1628; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_82 = _T_1358 ? _T_1358 : _T_1631; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_83 = _T_1358 ? _T_1267 : _T_1634; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_84 = _T_1358 ? _T_1613 : _T_1640; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_85 = _T_1358 ? _T_1645 : _T_1643; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_86 = _T_1358 ? _T_1532 : _T_1427; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_87 = _T_1358 ? _T_1536 : _T_1424; // @[NV_NVDLA_CSC_dl.scala 591:21:@741.4]
  assign _GEN_88 = _T_1608 ? _T_1242 : _T_1637; // @[NV_NVDLA_CSC_dl.scala 603:26:@755.4]
  assign _T_1667 = _T_831[8]; // @[NV_NVDLA_CSC_dl.scala 620:32:@765.4]
  assign _T_1668 = ~ _T_1667; // @[NV_NVDLA_CSC_dl.scala 620:22:@766.4]
  assign _T_1669 = _T_845[11:0]; // @[NV_NVDLA_CSC_dl.scala 620:49:@767.4]
  assign _T_1671 = _T_1668 ? _T_1669 : 12'h0; // @[NV_NVDLA_CSC_dl.scala 620:21:@768.4]
  assign _T_1673 = _T_1316 & _T_1269; // @[NV_NVDLA_CSC_dl.scala 622:34:@769.4]
  assign _GEN_701 = {{1'd0}, _T_1671}; // @[NV_NVDLA_CSC_dl.scala 622:64:@770.4]
  assign _T_1675 = _T_1648 + _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@770.4]
  assign _T_1676 = _T_1648 + _GEN_701; // @[NV_NVDLA_CSC_dl.scala 622:64:@771.4]
  assign _T_1677 = _T_1673 ? 13'h0 : _T_1676; // @[NV_NVDLA_CSC_dl.scala 622:19:@772.4]
  assign _T_1678 = _T_630 ? 13'h0 : _T_1677; // @[NV_NVDLA_CSC_dl.scala 621:19:@773.4]
  assign _T_1682 = _T_1648 != _T_1651; // @[NV_NVDLA_CSC_dl.scala 624:31:@777.4]
  assign _GEN_702 = {{2'd0}, _T_778}; // @[NV_NVDLA_CSC_dl.scala 627:32:@778.4]
  assign _T_1683 = _T_1539 * _GEN_702; // @[NV_NVDLA_CSC_dl.scala 627:32:@778.4]
  assign _T_1684 = _T_1683[12:0]; // @[NV_NVDLA_CSC_dl.scala 627:50:@779.4]
  assign _GEN_703 = {{7'd0}, _T_1264}; // @[NV_NVDLA_CSC_dl.scala 628:31:@780.4]
  assign _T_1685 = _GEN_703 * _T_785; // @[NV_NVDLA_CSC_dl.scala 628:31:@780.4]
  assign _T_1686 = _T_1685[12:0]; // @[NV_NVDLA_CSC_dl.scala 628:49:@781.4]
  assign _GEN_704 = {{10'd0}, _T_1279}; // @[NV_NVDLA_CSC_dl.scala 629:29:@782.4]
  assign _T_1687 = _GEN_704 * _T_1002; // @[NV_NVDLA_CSC_dl.scala 629:29:@782.4]
  assign _T_1688 = _T_1687[12:0]; // @[NV_NVDLA_CSC_dl.scala 629:47:@783.4]
  assign _GEN_705 = {{13'd0}, _T_1290}; // @[NV_NVDLA_CSC_dl.scala 630:47:@784.4]
  assign _T_1690 = _GEN_705 * _T_1009; // @[NV_NVDLA_CSC_dl.scala 630:47:@784.4]
  assign _T_1691 = _T_630 ? 17'h0 : _T_1690; // @[NV_NVDLA_CSC_dl.scala 630:21:@785.4]
  assign _T_1692 = _T_1691[12:0]; // @[NV_NVDLA_CSC_dl.scala 630:65:@786.4]
  assign _T_1693 = _T_831[9]; // @[NV_NVDLA_CSC_dl.scala 631:45:@787.4]
  assign _T_1694 = _T_630 | _T_1693; // @[NV_NVDLA_CSC_dl.scala 631:34:@788.4]
  assign _T_1695 = {_T_1694,_T_1358}; // @[Cat.scala 30:58:@789.4]
  assign _GEN_89 = _T_1394 ? _T_1678 : _T_1648; // @[NV_NVDLA_CSC_dl.scala 658:20:@806.4]
  assign _GEN_90 = _T_1682 ? _T_1648 : _T_1651; // @[NV_NVDLA_CSC_dl.scala 661:23:@809.4]
  assign _T_1715 = _T_1695[0]; // @[NV_NVDLA_CSC_dl.scala 664:19:@812.4]
  assign _GEN_91 = _T_1715 ? _T_1684 : _T_1654; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  assign _GEN_92 = _T_1715 ? _T_1686 : _T_1657; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  assign _GEN_93 = _T_1715 ? _T_1688 : _T_1660; // @[NV_NVDLA_CSC_dl.scala 664:23:@813.4]
  assign _T_1716 = _T_1695[1]; // @[NV_NVDLA_CSC_dl.scala 669:19:@818.4]
  assign _GEN_94 = _T_1716 ? _T_1692 : _T_1663; // @[NV_NVDLA_CSC_dl.scala 669:23:@819.4]
  assign _GEN_95 = _T_1358 ? _T_1714 : {{1'd0}, _T_1666}; // @[NV_NVDLA_CSC_dl.scala 672:20:@822.4]
  assign _T_1822 = _T_1654 + _T_1657; // @[NV_NVDLA_CSC_dl.scala 696:29:@850.4]
  assign _T_1823 = _T_1654 + _T_1657; // @[NV_NVDLA_CSC_dl.scala 696:29:@851.4]
  assign _T_1824 = _T_1823 + _T_1660; // @[NV_NVDLA_CSC_dl.scala 696:43:@852.4]
  assign _T_1825 = _T_1823 + _T_1660; // @[NV_NVDLA_CSC_dl.scala 696:43:@853.4]
  assign _T_1826 = _T_1825 + _T_1663; // @[NV_NVDLA_CSC_dl.scala 696:57:@854.4]
  assign _T_1827 = _T_1825 + _T_1663; // @[NV_NVDLA_CSC_dl.scala 696:57:@855.4]
  assign _GEN_706 = {{2'd0}, _T_1651}; // @[NV_NVDLA_CSC_dl.scala 697:40:@856.4]
  assign _T_1828 = _T_1076 + _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@856.4]
  assign _T_1829 = _T_1076 + _GEN_706; // @[NV_NVDLA_CSC_dl.scala 697:40:@857.4]
  assign _GEN_707 = {{2'd0}, _T_1827}; // @[NV_NVDLA_CSC_dl.scala 697:52:@858.4]
  assign _T_1830 = _T_1829 + _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@858.4]
  assign _T_1831 = _T_1829 + _GEN_707; // @[NV_NVDLA_CSC_dl.scala 697:52:@859.4]
  assign _GEN_708 = {{2'd0}, _T_1666}; // @[NV_NVDLA_CSC_dl.scala 697:64:@860.4]
  assign _T_1832 = _T_1831 + _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@860.4]
  assign _T_1833 = _T_1831 + _GEN_708; // @[NV_NVDLA_CSC_dl.scala 697:64:@861.4]
  assign _T_1840 = _T_1833 >= _GEN_678; // @[NV_NVDLA_CSC_dl.scala 698:45:@864.4]
  assign _T_1847 = _T_1833 - _GEN_678; // @[NV_NVDLA_CSC_dl.scala 699:42:@867.4]
  assign _T_1848 = $unsigned(_T_1847); // @[NV_NVDLA_CSC_dl.scala 699:42:@868.4]
  assign _T_1849 = _T_1848[14:0]; // @[NV_NVDLA_CSC_dl.scala 699:42:@869.4]
  assign _T_1850 = _T_630 | _T_1631; // @[NV_NVDLA_CSC_dl.scala 700:35:@870.4]
  assign _T_1856 = _T_1840 ? _T_1849 : _T_1833; // @[NV_NVDLA_CSC_dl.scala 701:25:@872.4]
  assign _T_1857 = _T_1850 ? 15'h1fff : _T_1856; // @[NV_NVDLA_CSC_dl.scala 700:25:@873.4]
  assign _T_1881 = 2'h3 == _T_1622; // @[Mux.scala 46:19:@883.4]
  assign _T_1882 = _T_1881 ? _T_1759_3 : 13'h0; // @[Mux.scala 46:16:@884.4]
  assign _T_1883 = 2'h2 == _T_1622; // @[Mux.scala 46:19:@885.4]
  assign _T_1884 = _T_1883 ? _T_1759_2 : _T_1882; // @[Mux.scala 46:16:@886.4]
  assign _T_1885 = 2'h1 == _T_1622; // @[Mux.scala 46:19:@887.4]
  assign _T_1886 = _T_1885 ? _T_1759_1 : _T_1884; // @[Mux.scala 46:16:@888.4]
  assign _T_1887 = 2'h0 == _T_1622; // @[Mux.scala 46:19:@889.4]
  assign _T_1888 = _T_1887 ? _T_1759_0 : _T_1886; // @[Mux.scala 46:16:@890.4]
  assign _GEN_712 = {{2'd0}, _T_1888}; // @[NV_NVDLA_CSC_dl.scala 708:65:@891.4]
  assign _T_1889 = _GEN_712 != _T_1857; // @[NV_NVDLA_CSC_dl.scala 708:65:@891.4]
  assign _T_1890 = _T_1889 | _T_1427; // @[NV_NVDLA_CSC_dl.scala 708:85:@892.4]
  assign _T_1891 = _T_1616 & _T_1890; // @[NV_NVDLA_CSC_dl.scala 708:43:@893.4]
  assign _T_1892 = _T_1616 | _T_1631; // @[NV_NVDLA_CSC_dl.scala 710:38:@894.4]
  assign _T_1894 = _T_1622 == 2'h0; // @[NV_NVDLA_CSC_dl.scala 710:78:@895.4]
  assign _T_1895 = _T_1892 & _T_1894; // @[NV_NVDLA_CSC_dl.scala 710:58:@896.4]
  assign _T_1896 = _T_630 | _T_1895; // @[NV_NVDLA_CSC_dl.scala 710:17:@897.4]
  assign _T_1899 = _T_1622 == 2'h1; // @[NV_NVDLA_CSC_dl.scala 710:78:@899.4]
  assign _T_1900 = _T_1892 & _T_1899; // @[NV_NVDLA_CSC_dl.scala 710:58:@900.4]
  assign _T_1901 = _T_630 | _T_1900; // @[NV_NVDLA_CSC_dl.scala 710:17:@901.4]
  assign _T_1904 = _T_1622 == 2'h2; // @[NV_NVDLA_CSC_dl.scala 710:78:@903.4]
  assign _T_1905 = _T_1892 & _T_1904; // @[NV_NVDLA_CSC_dl.scala 710:58:@904.4]
  assign _T_1906 = _T_630 | _T_1905; // @[NV_NVDLA_CSC_dl.scala 710:17:@905.4]
  assign _T_1909 = _T_1622 == 2'h3; // @[NV_NVDLA_CSC_dl.scala 710:78:@907.4]
  assign _T_1910 = _T_1892 & _T_1909; // @[NV_NVDLA_CSC_dl.scala 710:58:@908.4]
  assign _T_1911 = _T_630 | _T_1910; // @[NV_NVDLA_CSC_dl.scala 710:17:@909.4]
  assign _GEN_96 = _T_1896 ? _T_1857 : {{2'd0}, _T_1759_0}; // @[NV_NVDLA_CSC_dl.scala 717:35:@915.4]
  assign _GEN_97 = _T_1901 ? _T_1857 : {{2'd0}, _T_1759_1}; // @[NV_NVDLA_CSC_dl.scala 717:35:@918.4]
  assign _GEN_98 = _T_1906 ? _T_1857 : {{2'd0}, _T_1759_2}; // @[NV_NVDLA_CSC_dl.scala 717:35:@921.4]
  assign _GEN_99 = _T_1911 ? _T_1857 : {{2'd0}, _T_1759_3}; // @[NV_NVDLA_CSC_dl.scala 717:35:@924.4]
  assign _T_1922 = _T_630 | _T_1891; // @[NV_NVDLA_CSC_dl.scala 723:14:@928.4]
  assign _GEN_100 = _T_1922 ? _T_1857 : _T_1785; // @[NV_NVDLA_CSC_dl.scala 723:34:@929.4]
  assign _GEN_101 = _T_1335 ? _T_1619 : _T_1794; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_102 = _T_1335 ? _T_1622 : _T_1797; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_103 = _T_1335 ? _T_1625 : _T_1800; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_104 = _T_1335 ? _T_1628 : _T_1803; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_105 = _T_1335 ? _T_1361 : _T_1806; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_106 = _T_1335 ? _T_1631 : _T_1809; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_107 = _T_1335 ? _T_1634 : _T_1812; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_108 = _T_1335 ? _T_1637 : _T_1815; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_109 = _T_1335 ? _T_1643 : _T_1818; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _GEN_110 = _T_1335 ? _T_1640 : {{8'd0}, _T_1335}; // @[NV_NVDLA_CSC_dl.scala 730:24:@936.4]
  assign _T_1932 = {1'h0,_T_1803,_T_1800,_T_1797,_T_1794}; // @[Cat.scala 30:58:@956.4]
  assign _T_1938 = {_T_1821,_T_1818,_T_1815,_T_1809,_T_1812,_T_1806,_T_1932}; // @[Cat.scala 30:58:@962.4]
  assign _GEN_111 = _T_1788 ? _T_1938 : _T_1963; // @[NV_NVDLA_CSC_dl.scala 775:33:@1004.4]
  assign _GEN_114 = _T_1943 ? _T_1963 : _T_1966; // @[NV_NVDLA_CSC_dl.scala 775:33:@1013.4]
  assign _GEN_117 = _T_1946 ? _T_1966 : _T_1969; // @[NV_NVDLA_CSC_dl.scala 775:33:@1022.4]
  assign _GEN_120 = _T_1949 ? _T_1969 : _T_1972; // @[NV_NVDLA_CSC_dl.scala 775:33:@1031.4]
  assign _GEN_123 = _T_1952 ? _T_1972 : _T_1975; // @[NV_NVDLA_CSC_dl.scala 775:33:@1040.4]
  assign _GEN_126 = _T_1955 ? _T_1975 : _T_1978; // @[NV_NVDLA_CSC_dl.scala 775:33:@1049.4]
  assign _T_2039 = _T_1978[1:0]; // @[NV_NVDLA_CSC_dl.scala 792:41:@1057.4]
  assign _T_2040 = _T_1978[3:2]; // @[NV_NVDLA_CSC_dl.scala 793:41:@1058.4]
  assign _T_2041 = _T_1978[4]; // @[NV_NVDLA_CSC_dl.scala 794:41:@1059.4]
  assign _T_2042 = _T_1978[5]; // @[NV_NVDLA_CSC_dl.scala 795:42:@1060.4]
  assign _T_2043 = _T_1978[14:7]; // @[NV_NVDLA_CSC_dl.scala 796:41:@1061.4]
  assign _T_2044 = _T_1978[16:15]; // @[NV_NVDLA_CSC_dl.scala 797:45:@1062.4]
  assign _T_2047 = _T_1978[19]; // @[NV_NVDLA_CSC_dl.scala 800:39:@1065.4]
  assign _T_2048 = _T_1978[28:20]; // @[NV_NVDLA_CSC_dl.scala 801:40:@1066.4]
  assign _T_2105 = _T_831[12]; // @[NV_NVDLA_CSC_dl.scala 831:69:@1094.4]
  assign _T_2106 = _T_2105 & io_sc2buf_dat_rd_data_valid; // @[NV_NVDLA_CSC_dl.scala 831:74:@1095.4]
  assign _T_2107 = ~ _T_2051; // @[NV_NVDLA_CSC_dl.scala 831:90:@1096.4]
  assign _T_2108 = _T_2106 & _T_2107; // @[NV_NVDLA_CSC_dl.scala 831:88:@1097.4]
  assign _T_2148 = io_sc2buf_dat_rd_data_valid ? 1'h0 : _T_2051; // @[NV_NVDLA_CSC_dl.scala 846:22:@1131.4]
  assign _T_2162 = io_sc2buf_dat_rd_data_valid ? _T_2051 : _T_2063; // @[NV_NVDLA_CSC_dl.scala 850:48:@1142.4]
  assign _T_2163 = _T_2108 ? 1'h0 : _T_2162; // @[NV_NVDLA_CSC_dl.scala 850:22:@1143.4]
  assign _T_2240 = {_T_2048,_T_2047,_T_2044,_T_2043,1'h0,_T_2042,_T_2041,_T_2040,_T_2039}; // @[Cat.scala 30:58:@1210.4]
  assign _GEN_137 = _T_1958 ? _T_2240 : _T_2222; // @[NV_NVDLA_CSC_dl.scala 889:28:@1213.4]
  assign _GEN_138 = _T_2208 ? _T_2222 : _T_2225; // @[NV_NVDLA_CSC_dl.scala 889:28:@1217.4]
  assign _GEN_139 = _T_2211 ? _T_2225 : _T_2228; // @[NV_NVDLA_CSC_dl.scala 889:28:@1221.4]
  assign _GEN_140 = _T_2214 ? _T_2228 : _T_2231; // @[NV_NVDLA_CSC_dl.scala 889:28:@1225.4]
  assign _T_2269 = _T_2222[4]; // @[NV_NVDLA_CSC_dl.scala 907:39:@1251.4]
  assign _T_2270 = _T_2225[4]; // @[NV_NVDLA_CSC_dl.scala 908:39:@1252.4]
  assign _T_2271 = _T_2228[4]; // @[NV_NVDLA_CSC_dl.scala 909:39:@1253.4]
  assign _T_2272 = _T_2231[4]; // @[NV_NVDLA_CSC_dl.scala 910:39:@1254.4]
  assign _T_2273 = _T_2222[26:18]; // @[NV_NVDLA_CSC_dl.scala 912:38:@1255.4]
  assign _T_2274 = _T_2225[26:18]; // @[NV_NVDLA_CSC_dl.scala 913:38:@1256.4]
  assign _T_2275 = _T_2228[26:18]; // @[NV_NVDLA_CSC_dl.scala 914:38:@1257.4]
  assign _T_2276 = _T_2231[26:18]; // @[NV_NVDLA_CSC_dl.scala 915:38:@1258.4]
  assign _T_2277 = _T_2273[6]; // @[NV_NVDLA_CSC_dl.scala 917:44:@1259.4]
  assign _T_2278 = _T_2274[6]; // @[NV_NVDLA_CSC_dl.scala 918:44:@1260.4]
  assign _T_2279 = _T_2275[6]; // @[NV_NVDLA_CSC_dl.scala 919:44:@1261.4]
  assign _T_2280 = _T_2276[6]; // @[NV_NVDLA_CSC_dl.scala 920:44:@1262.4]
  assign _T_2281 = _T_2268[1:0]; // @[NV_NVDLA_CSC_dl.scala 923:31:@1263.4]
  assign _T_2285 = _T_2268[14:7]; // @[NV_NVDLA_CSC_dl.scala 927:31:@1267.4]
  assign _T_2286 = _T_2268[16:15]; // @[NV_NVDLA_CSC_dl.scala 928:35:@1268.4]
  assign _T_2296 = io_sc2buf_dat_rd_data_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl.scala 939:29:@1277.4]
  assign _T_2307 = _T_960 > 7'h40; // @[NV_NVDLA_CSC_dl.scala 944:50:@1281.4]
  assign _GEN_713 = {{1'd0}, _T_960}; // @[NV_NVDLA_CSC_dl.scala 944:111:@1282.4]
  assign _T_2309 = _T_2182 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@1282.4]
  assign _T_2310 = _T_2182 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 944:111:@1283.4]
  assign _T_2311 = _T_2310 - _T_2296; // @[NV_NVDLA_CSC_dl.scala 944:133:@1284.4]
  assign _T_2312 = $unsigned(_T_2311); // @[NV_NVDLA_CSC_dl.scala 944:133:@1285.4]
  assign _T_2313 = _T_2312[7:0]; // @[NV_NVDLA_CSC_dl.scala 944:133:@1286.4]
  assign _T_2314 = _T_2307 ? 8'h40 : _T_2313; // @[NV_NVDLA_CSC_dl.scala 944:29:@1287.4]
  assign _T_2318 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 945:111:@1289.4]
  assign _T_2319 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 945:111:@1290.4]
  assign _T_2320 = _T_2319 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 945:133:@1291.4]
  assign _T_2321 = $unsigned(_T_2320); // @[NV_NVDLA_CSC_dl.scala 945:133:@1292.4]
  assign _T_2322 = _T_2321[7:0]; // @[NV_NVDLA_CSC_dl.scala 945:133:@1293.4]
  assign _T_2323 = _T_2307 ? 8'h40 : _T_2322; // @[NV_NVDLA_CSC_dl.scala 945:29:@1294.4]
  assign _T_2327 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 946:111:@1296.4]
  assign _T_2328 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 946:111:@1297.4]
  assign _T_2329 = _T_2328 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 946:133:@1298.4]
  assign _T_2330 = $unsigned(_T_2329); // @[NV_NVDLA_CSC_dl.scala 946:133:@1299.4]
  assign _T_2331 = _T_2330[7:0]; // @[NV_NVDLA_CSC_dl.scala 946:133:@1300.4]
  assign _T_2332 = _T_2307 ? 8'h40 : _T_2331; // @[NV_NVDLA_CSC_dl.scala 946:29:@1301.4]
  assign _T_2336 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 947:111:@1303.4]
  assign _T_2337 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl.scala 947:111:@1304.4]
  assign _T_2338 = _T_2337 - 8'h0; // @[NV_NVDLA_CSC_dl.scala 947:133:@1305.4]
  assign _T_2339 = $unsigned(_T_2338); // @[NV_NVDLA_CSC_dl.scala 947:133:@1306.4]
  assign _T_2340 = _T_2339[7:0]; // @[NV_NVDLA_CSC_dl.scala 947:133:@1307.4]
  assign _T_2341 = _T_2307 ? 8'h40 : _T_2340; // @[NV_NVDLA_CSC_dl.scala 947:29:@1308.4]
  assign _T_2343 = ~ _T_2269; // @[NV_NVDLA_CSC_dl.scala 956:52:@1309.4]
  assign _T_2344 = _T_2277 & _T_2343; // @[NV_NVDLA_CSC_dl.scala 956:50:@1310.4]
  assign _T_2345 = _T_2277 & _T_2269; // @[NV_NVDLA_CSC_dl.scala 957:50:@1311.4]
  assign _T_2350 = _T_2345 ? 8'h40 : _T_2314; // @[NV_NVDLA_CSC_dl.scala 957:27:@1314.4]
  assign _T_2351 = _T_2344 ? _T_2194 : _T_2350; // @[NV_NVDLA_CSC_dl.scala 956:27:@1315.4]
  assign _T_2352 = _T_630 ? 8'h40 : _T_2351; // @[NV_NVDLA_CSC_dl.scala 955:27:@1316.4]
  assign _T_2354 = ~ _T_2270; // @[NV_NVDLA_CSC_dl.scala 961:52:@1317.4]
  assign _T_2355 = _T_2278 & _T_2354; // @[NV_NVDLA_CSC_dl.scala 961:50:@1318.4]
  assign _T_2356 = _T_2278 & _T_2270; // @[NV_NVDLA_CSC_dl.scala 962:50:@1319.4]
  assign _T_2361 = _T_2356 ? 8'h40 : _T_2323; // @[NV_NVDLA_CSC_dl.scala 962:27:@1322.4]
  assign _T_2362 = _T_2355 ? _T_2197 : _T_2361; // @[NV_NVDLA_CSC_dl.scala 961:27:@1323.4]
  assign _T_2363 = _T_630 ? 8'h40 : _T_2362; // @[NV_NVDLA_CSC_dl.scala 960:27:@1324.4]
  assign _T_2365 = ~ _T_2271; // @[NV_NVDLA_CSC_dl.scala 966:52:@1325.4]
  assign _T_2366 = _T_2279 & _T_2365; // @[NV_NVDLA_CSC_dl.scala 966:50:@1326.4]
  assign _T_2367 = _T_2279 & _T_2271; // @[NV_NVDLA_CSC_dl.scala 967:50:@1327.4]
  assign _T_2372 = _T_2367 ? 8'h40 : _T_2332; // @[NV_NVDLA_CSC_dl.scala 967:27:@1330.4]
  assign _T_2373 = _T_2366 ? _T_2200 : _T_2372; // @[NV_NVDLA_CSC_dl.scala 966:27:@1331.4]
  assign _T_2374 = _T_630 ? 8'h40 : _T_2373; // @[NV_NVDLA_CSC_dl.scala 965:27:@1332.4]
  assign _T_2376 = ~ _T_2272; // @[NV_NVDLA_CSC_dl.scala 971:52:@1333.4]
  assign _T_2377 = _T_2280 & _T_2376; // @[NV_NVDLA_CSC_dl.scala 971:50:@1334.4]
  assign _T_2378 = _T_2280 & _T_2272; // @[NV_NVDLA_CSC_dl.scala 972:50:@1335.4]
  assign _T_2383 = _T_2378 ? 8'h40 : _T_2341; // @[NV_NVDLA_CSC_dl.scala 972:27:@1338.4]
  assign _T_2384 = _T_2377 ? _T_2203 : _T_2383; // @[NV_NVDLA_CSC_dl.scala 971:27:@1339.4]
  assign _T_2385 = _T_630 ? 8'h40 : _T_2384; // @[NV_NVDLA_CSC_dl.scala 970:27:@1340.4]
  assign _T_2386 = _T_831[17]; // @[NV_NVDLA_CSC_dl.scala 976:46:@1341.4]
  assign _T_2387 = _T_2386 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 976:51:@1342.4]
  assign _T_2388 = _T_630 | _T_2387; // @[NV_NVDLA_CSC_dl.scala 976:34:@1343.4]
  assign _T_2389 = _T_831[18]; // @[NV_NVDLA_CSC_dl.scala 977:46:@1344.4]
  assign _T_2390 = _T_2389 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 977:51:@1345.4]
  assign _T_2392 = _T_884 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 977:87:@1346.4]
  assign _T_2393 = _T_2390 & _T_2392; // @[NV_NVDLA_CSC_dl.scala 977:69:@1347.4]
  assign _T_2394 = _T_630 | _T_2393; // @[NV_NVDLA_CSC_dl.scala 977:34:@1348.4]
  assign _T_2395 = _T_831[19]; // @[NV_NVDLA_CSC_dl.scala 978:46:@1349.4]
  assign _T_2396 = _T_2395 & _T_2214; // @[NV_NVDLA_CSC_dl.scala 978:51:@1350.4]
  assign _T_2398 = _T_884 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 978:87:@1351.4]
  assign _T_2399 = _T_2396 & _T_2398; // @[NV_NVDLA_CSC_dl.scala 978:69:@1352.4]
  assign _T_2400 = _T_630 | _T_2399; // @[NV_NVDLA_CSC_dl.scala 978:34:@1353.4]
  assign _T_2401 = _T_831[20]; // @[NV_NVDLA_CSC_dl.scala 979:46:@1354.4]
  assign _T_2402 = _T_2401 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 979:51:@1355.4]
  assign _T_2405 = _T_2402 & _T_2398; // @[NV_NVDLA_CSC_dl.scala 979:69:@1357.4]
  assign _T_2406 = _T_630 | _T_2405; // @[NV_NVDLA_CSC_dl.scala 979:34:@1358.4]
  assign _T_2407 = _T_831[21]; // @[NV_NVDLA_CSC_dl.scala 981:50:@1359.4]
  assign _T_2408 = _T_2407 & _T_2208; // @[NV_NVDLA_CSC_dl.scala 981:55:@1360.4]
  assign _T_2409 = _T_2408 & _T_2277; // @[NV_NVDLA_CSC_dl.scala 981:73:@1361.4]
  assign _T_2410 = _T_2409 & _T_2269; // @[NV_NVDLA_CSC_dl.scala 981:97:@1362.4]
  assign _T_2411 = _T_630 | _T_2410; // @[NV_NVDLA_CSC_dl.scala 981:38:@1363.4]
  assign _T_2412 = _T_831[22]; // @[NV_NVDLA_CSC_dl.scala 982:50:@1364.4]
  assign _T_2413 = _T_2412 & _T_2211; // @[NV_NVDLA_CSC_dl.scala 982:55:@1365.4]
  assign _T_2414 = _T_2413 & _T_2278; // @[NV_NVDLA_CSC_dl.scala 982:73:@1366.4]
  assign _T_2415 = _T_2414 & _T_2270; // @[NV_NVDLA_CSC_dl.scala 982:97:@1367.4]
  assign _T_2417 = _T_887 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 982:138:@1368.4]
  assign _T_2418 = _T_2415 & _T_2417; // @[NV_NVDLA_CSC_dl.scala 982:120:@1369.4]
  assign _T_2419 = _T_630 | _T_2418; // @[NV_NVDLA_CSC_dl.scala 982:38:@1370.4]
  assign _T_2420 = _T_831[23]; // @[NV_NVDLA_CSC_dl.scala 983:50:@1371.4]
  assign _T_2421 = _T_2420 & _T_2214; // @[NV_NVDLA_CSC_dl.scala 983:55:@1372.4]
  assign _T_2422 = _T_2421 & _T_2279; // @[NV_NVDLA_CSC_dl.scala 983:73:@1373.4]
  assign _T_2423 = _T_2422 & _T_2271; // @[NV_NVDLA_CSC_dl.scala 983:97:@1374.4]
  assign _T_2425 = _T_887 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 983:138:@1375.4]
  assign _T_2426 = _T_2423 & _T_2425; // @[NV_NVDLA_CSC_dl.scala 983:120:@1376.4]
  assign _T_2427 = _T_630 | _T_2426; // @[NV_NVDLA_CSC_dl.scala 983:38:@1377.4]
  assign _T_2428 = _T_831[24]; // @[NV_NVDLA_CSC_dl.scala 984:50:@1378.4]
  assign _T_2429 = _T_2428 & _T_2217; // @[NV_NVDLA_CSC_dl.scala 984:55:@1379.4]
  assign _T_2430 = _T_2429 & _T_2280; // @[NV_NVDLA_CSC_dl.scala 984:73:@1380.4]
  assign _T_2431 = _T_2430 & _T_2272; // @[NV_NVDLA_CSC_dl.scala 984:97:@1381.4]
  assign _T_2434 = _T_2431 & _T_2425; // @[NV_NVDLA_CSC_dl.scala 984:120:@1383.4]
  assign _T_2435 = _T_630 | _T_2434; // @[NV_NVDLA_CSC_dl.scala 984:38:@1384.4]
  assign _GEN_141 = _T_2388 ? _T_2352 : _T_2182; // @[NV_NVDLA_CSC_dl.scala 986:24:@1385.4]
  assign _GEN_142 = _T_2394 ? _T_2363 : _T_2185; // @[NV_NVDLA_CSC_dl.scala 987:24:@1388.4]
  assign _GEN_143 = _T_2400 ? _T_2374 : _T_2188; // @[NV_NVDLA_CSC_dl.scala 988:24:@1391.4]
  assign _GEN_144 = _T_2406 ? _T_2385 : _T_2191; // @[NV_NVDLA_CSC_dl.scala 989:24:@1394.4]
  assign _GEN_145 = _T_2411 ? _T_2352 : _T_2194; // @[NV_NVDLA_CSC_dl.scala 990:28:@1397.4]
  assign _GEN_146 = _T_2419 ? _T_2363 : _T_2197; // @[NV_NVDLA_CSC_dl.scala 991:28:@1400.4]
  assign _GEN_147 = _T_2427 ? _T_2374 : _T_2200; // @[NV_NVDLA_CSC_dl.scala 992:28:@1403.4]
  assign _GEN_148 = _T_2435 ? _T_2385 : _T_2203; // @[NV_NVDLA_CSC_dl.scala 993:28:@1406.4]
  assign _T_2436 = _T_988[7:0]; // @[NV_NVDLA_CSC_dl.scala 1002:55:@1409.4]
  assign _T_2439 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436}; // @[Cat.scala 30:58:@1412.4]
  assign _T_2440 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2439}; // @[Cat.scala 30:58:@1413.4]
  assign _T_2441 = {_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2436,_T_2439,_T_2440}; // @[Cat.scala 30:58:@1414.4]
  assign _T_2442 = {_T_2441,_T_2441}; // @[Cat.scala 30:58:@1415.4]
  assign _T_2443 = _T_2051 ? _T_2442 : _T_2074; // @[NV_NVDLA_CSC_dl.scala 1004:23:@1416.4]
  assign _T_2447 = _T_2063 ? _T_2442 : _T_2082; // @[NV_NVDLA_CSC_dl.scala 1009:23:@1420.4]
  assign _T_2453 = _T_831[26]; // @[NV_NVDLA_CSC_dl.scala 1022:37:@1425.4]
  assign _T_2456 = _T_2285 <= 8'h20; // @[NV_NVDLA_CSC_dl.scala 1023:43:@1426.4]
  assign _T_2457 = _T_2281[0]; // @[NV_NVDLA_CSC_dl.scala 1023:87:@1427.4]
  assign _T_2459 = _T_2457 == 1'h0; // @[NV_NVDLA_CSC_dl.scala 1023:91:@1428.4]
  assign _T_2460 = _T_2456 & _T_2459; // @[NV_NVDLA_CSC_dl.scala 1023:72:@1429.4]
  assign _T_2462 = _T_2443[255:0]; // @[NV_NVDLA_CSC_dl.scala 1023:171:@1430.4]
  assign _T_2463 = {256'h0,_T_2462}; // @[Cat.scala 30:58:@1431.4]
  assign _T_2469 = _T_2456 & _T_2457; // @[NV_NVDLA_CSC_dl.scala 1024:72:@1435.4]
  assign _T_2471 = _T_2443[511:256]; // @[NV_NVDLA_CSC_dl.scala 1024:171:@1436.4]
  assign _T_2472 = {256'h0,_T_2471}; // @[Cat.scala 30:58:@1437.4]
  assign _T_2473 = _T_2469 ? _T_2472 : _T_2443; // @[NV_NVDLA_CSC_dl.scala 1024:27:@1438.4]
  assign _T_2474 = _T_2460 ? _T_2463 : _T_2473; // @[NV_NVDLA_CSC_dl.scala 1023:27:@1439.4]
  assign _T_2475 = _T_2453 ? 512'h0 : _T_2474; // @[NV_NVDLA_CSC_dl.scala 1022:27:@1440.4]
  assign _T_2546 = _T_2475[7:0]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1443.4]
  assign _T_2547 = _T_2475[15:8]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1445.4]
  assign _T_2548 = _T_2475[23:16]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1447.4]
  assign _T_2549 = _T_2475[31:24]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1449.4]
  assign _T_2550 = _T_2475[39:32]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1451.4]
  assign _T_2551 = _T_2475[47:40]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1453.4]
  assign _T_2552 = _T_2475[55:48]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1455.4]
  assign _T_2553 = _T_2475[63:56]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1457.4]
  assign _T_2554 = _T_2475[71:64]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1459.4]
  assign _T_2555 = _T_2475[79:72]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1461.4]
  assign _T_2556 = _T_2475[87:80]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1463.4]
  assign _T_2557 = _T_2475[95:88]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1465.4]
  assign _T_2558 = _T_2475[103:96]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1467.4]
  assign _T_2559 = _T_2475[111:104]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1469.4]
  assign _T_2560 = _T_2475[119:112]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1471.4]
  assign _T_2561 = _T_2475[127:120]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1473.4]
  assign _T_2562 = _T_2475[135:128]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1475.4]
  assign _T_2563 = _T_2475[143:136]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1477.4]
  assign _T_2564 = _T_2475[151:144]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1479.4]
  assign _T_2565 = _T_2475[159:152]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1481.4]
  assign _T_2566 = _T_2475[167:160]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1483.4]
  assign _T_2567 = _T_2475[175:168]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1485.4]
  assign _T_2568 = _T_2475[183:176]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1487.4]
  assign _T_2569 = _T_2475[191:184]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1489.4]
  assign _T_2570 = _T_2475[199:192]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1491.4]
  assign _T_2571 = _T_2475[207:200]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1493.4]
  assign _T_2572 = _T_2475[215:208]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1495.4]
  assign _T_2573 = _T_2475[223:216]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1497.4]
  assign _T_2574 = _T_2475[231:224]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1499.4]
  assign _T_2575 = _T_2475[239:232]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1501.4]
  assign _T_2576 = _T_2475[247:240]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1503.4]
  assign _T_2577 = _T_2475[255:248]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1505.4]
  assign _T_2578 = _T_2475[263:256]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1507.4]
  assign _T_2579 = _T_2475[271:264]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1509.4]
  assign _T_2580 = _T_2475[279:272]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1511.4]
  assign _T_2581 = _T_2475[287:280]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1513.4]
  assign _T_2582 = _T_2475[295:288]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1515.4]
  assign _T_2583 = _T_2475[303:296]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1517.4]
  assign _T_2584 = _T_2475[311:304]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1519.4]
  assign _T_2585 = _T_2475[319:312]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1521.4]
  assign _T_2586 = _T_2475[327:320]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1523.4]
  assign _T_2587 = _T_2475[335:328]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1525.4]
  assign _T_2588 = _T_2475[343:336]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1527.4]
  assign _T_2589 = _T_2475[351:344]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1529.4]
  assign _T_2590 = _T_2475[359:352]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1531.4]
  assign _T_2591 = _T_2475[367:360]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1533.4]
  assign _T_2592 = _T_2475[375:368]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1535.4]
  assign _T_2593 = _T_2475[383:376]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1537.4]
  assign _T_2594 = _T_2475[391:384]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1539.4]
  assign _T_2595 = _T_2475[399:392]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1541.4]
  assign _T_2596 = _T_2475[407:400]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1543.4]
  assign _T_2597 = _T_2475[415:408]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1545.4]
  assign _T_2598 = _T_2475[423:416]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1547.4]
  assign _T_2599 = _T_2475[431:424]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1549.4]
  assign _T_2600 = _T_2475[439:432]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1551.4]
  assign _T_2601 = _T_2475[447:440]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1553.4]
  assign _T_2602 = _T_2475[455:448]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1555.4]
  assign _T_2603 = _T_2475[463:456]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1557.4]
  assign _T_2604 = _T_2475[471:464]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1559.4]
  assign _T_2605 = _T_2475[479:472]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1561.4]
  assign _T_2606 = _T_2475[487:480]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1563.4]
  assign _T_2607 = _T_2475[495:488]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1565.4]
  assign _T_2608 = _T_2475[503:496]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1567.4]
  assign _T_2609 = _T_2475[511:504]; // @[NV_NVDLA_CSC_dl.scala 1040:39:@1569.4]
  assign _T_2622 = _T_831[27]; // @[NV_NVDLA_CSC_dl.scala 1053:39:@1577.4]
  assign _T_2623 = ~ _T_2622; // @[NV_NVDLA_CSC_dl.scala 1053:29:@1578.4]
  assign _T_2625 = {_T_2443,_T_2447}; // @[Cat.scala 30:58:@1579.4]
  assign _T_2626 = _T_2623 ? 1024'h0 : _T_2625; // @[NV_NVDLA_CSC_dl.scala 1053:28:@1580.4]
  assign _T_2627 = _T_831[28]; // @[NV_NVDLA_CSC_dl.scala 1054:39:@1581.4]
  assign _T_2628 = ~ _T_2627; // @[NV_NVDLA_CSC_dl.scala 1054:29:@1582.4]
  assign _T_2630 = {_T_2441,_T_2441,_T_2441,_T_2441}; // @[Cat.scala 30:58:@1583.4]
  assign _T_2631 = _T_2628 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1054:28:@1584.4]
  assign _T_2632 = _T_831[29]; // @[NV_NVDLA_CSC_dl.scala 1055:39:@1585.4]
  assign _T_2633 = ~ _T_2632; // @[NV_NVDLA_CSC_dl.scala 1055:29:@1586.4]
  assign _T_2636 = _T_2633 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1055:28:@1588.4]
  assign _T_2637 = _T_831[30]; // @[NV_NVDLA_CSC_dl.scala 1056:39:@1589.4]
  assign _T_2638 = ~ _T_2637; // @[NV_NVDLA_CSC_dl.scala 1056:29:@1590.4]
  assign _T_2641 = _T_2638 ? 1024'h0 : _T_2630; // @[NV_NVDLA_CSC_dl.scala 1056:28:@1592.4]
  assign _T_2643 = {_T_2182,3'h0}; // @[Cat.scala 30:58:@1593.4]
  assign _T_2644 = _T_2626 >> _T_2643; // @[NV_NVDLA_CSC_dl.scala 1058:41:@1594.4]
  assign _T_2645 = _T_2644[511:0]; // @[NV_NVDLA_CSC_dl.scala 1058:82:@1595.4]
  assign _T_2647 = {_T_2185,3'h0}; // @[Cat.scala 30:58:@1596.4]
  assign _T_2648 = _T_2631 >> _T_2647; // @[NV_NVDLA_CSC_dl.scala 1059:41:@1597.4]
  assign _T_2649 = _T_2648[511:0]; // @[NV_NVDLA_CSC_dl.scala 1059:82:@1598.4]
  assign _T_2651 = {_T_2188,3'h0}; // @[Cat.scala 30:58:@1599.4]
  assign _T_2652 = _T_2636 >> _T_2651; // @[NV_NVDLA_CSC_dl.scala 1060:41:@1600.4]
  assign _T_2653 = _T_2652[511:0]; // @[NV_NVDLA_CSC_dl.scala 1060:82:@1601.4]
  assign _T_2655 = {_T_2191,3'h0}; // @[Cat.scala 30:58:@1602.4]
  assign _T_2656 = _T_2641 >> _T_2655; // @[NV_NVDLA_CSC_dl.scala 1061:41:@1603.4]
  assign _T_2657 = _T_2656[511:0]; // @[NV_NVDLA_CSC_dl.scala 1061:82:@1604.4]
  assign _T_2658 = _T_831[32]; // @[NV_NVDLA_CSC_dl.scala 1063:36:@1605.4]
  assign _T_2659 = ~ _T_2658; // @[NV_NVDLA_CSC_dl.scala 1063:26:@1606.4]
  assign _T_2662 = _T_893 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1064:41:@1607.4]
  assign _T_2663 = _T_2657[127:0]; // @[NV_NVDLA_CSC_dl.scala 1064:81:@1608.4]
  assign _T_2669 = {_T_2663,_T_2621,_T_2619,_T_2615}; // @[Cat.scala 30:58:@1614.4]
  assign _T_2671 = _T_893 == 3'h2; // @[NV_NVDLA_CSC_dl.scala 1065:41:@1615.4]
  assign _T_2672 = _T_2649[255:0]; // @[NV_NVDLA_CSC_dl.scala 1065:81:@1616.4]
  assign _T_2674 = {_T_2672,_T_2611}; // @[Cat.scala 30:58:@1618.4]
  assign _T_2676 = _T_2671 ? _T_2674 : _T_2645; // @[NV_NVDLA_CSC_dl.scala 1065:25:@1620.4]
  assign _T_2677 = _T_2662 ? _T_2669 : _T_2676; // @[NV_NVDLA_CSC_dl.scala 1064:25:@1621.4]
  assign _T_2678 = _T_2659 ? 512'h0 : _T_2677; // @[NV_NVDLA_CSC_dl.scala 1063:25:@1622.4]
  assign _T_2749 = _T_2678[7:0]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1624.4]
  assign _T_2750 = _T_2678[15:8]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1626.4]
  assign _T_2751 = _T_2678[23:16]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1628.4]
  assign _T_2752 = _T_2678[31:24]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1630.4]
  assign _T_2753 = _T_2678[39:32]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1632.4]
  assign _T_2754 = _T_2678[47:40]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1634.4]
  assign _T_2755 = _T_2678[55:48]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1636.4]
  assign _T_2756 = _T_2678[63:56]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1638.4]
  assign _T_2757 = _T_2678[71:64]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1640.4]
  assign _T_2758 = _T_2678[79:72]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1642.4]
  assign _T_2759 = _T_2678[87:80]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1644.4]
  assign _T_2760 = _T_2678[95:88]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1646.4]
  assign _T_2761 = _T_2678[103:96]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1648.4]
  assign _T_2762 = _T_2678[111:104]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1650.4]
  assign _T_2763 = _T_2678[119:112]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1652.4]
  assign _T_2764 = _T_2678[127:120]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1654.4]
  assign _T_2765 = _T_2678[135:128]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1656.4]
  assign _T_2766 = _T_2678[143:136]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1658.4]
  assign _T_2767 = _T_2678[151:144]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1660.4]
  assign _T_2768 = _T_2678[159:152]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1662.4]
  assign _T_2769 = _T_2678[167:160]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1664.4]
  assign _T_2770 = _T_2678[175:168]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1666.4]
  assign _T_2771 = _T_2678[183:176]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1668.4]
  assign _T_2772 = _T_2678[191:184]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1670.4]
  assign _T_2773 = _T_2678[199:192]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1672.4]
  assign _T_2774 = _T_2678[207:200]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1674.4]
  assign _T_2775 = _T_2678[215:208]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1676.4]
  assign _T_2776 = _T_2678[223:216]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1678.4]
  assign _T_2777 = _T_2678[231:224]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1680.4]
  assign _T_2778 = _T_2678[239:232]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1682.4]
  assign _T_2779 = _T_2678[247:240]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1684.4]
  assign _T_2780 = _T_2678[255:248]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1686.4]
  assign _T_2781 = _T_2678[263:256]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1688.4]
  assign _T_2782 = _T_2678[271:264]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1690.4]
  assign _T_2783 = _T_2678[279:272]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1692.4]
  assign _T_2784 = _T_2678[287:280]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1694.4]
  assign _T_2785 = _T_2678[295:288]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1696.4]
  assign _T_2786 = _T_2678[303:296]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1698.4]
  assign _T_2787 = _T_2678[311:304]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1700.4]
  assign _T_2788 = _T_2678[319:312]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1702.4]
  assign _T_2789 = _T_2678[327:320]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1704.4]
  assign _T_2790 = _T_2678[335:328]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1706.4]
  assign _T_2791 = _T_2678[343:336]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1708.4]
  assign _T_2792 = _T_2678[351:344]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1710.4]
  assign _T_2793 = _T_2678[359:352]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1712.4]
  assign _T_2794 = _T_2678[367:360]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1714.4]
  assign _T_2795 = _T_2678[375:368]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1716.4]
  assign _T_2796 = _T_2678[383:376]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1718.4]
  assign _T_2797 = _T_2678[391:384]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1720.4]
  assign _T_2798 = _T_2678[399:392]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1722.4]
  assign _T_2799 = _T_2678[407:400]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1724.4]
  assign _T_2800 = _T_2678[415:408]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1726.4]
  assign _T_2801 = _T_2678[423:416]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1728.4]
  assign _T_2802 = _T_2678[431:424]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1730.4]
  assign _T_2803 = _T_2678[439:432]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1732.4]
  assign _T_2804 = _T_2678[447:440]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1734.4]
  assign _T_2805 = _T_2678[455:448]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1736.4]
  assign _T_2806 = _T_2678[463:456]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1738.4]
  assign _T_2807 = _T_2678[471:464]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1740.4]
  assign _T_2808 = _T_2678[479:472]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1742.4]
  assign _T_2809 = _T_2678[487:480]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1744.4]
  assign _T_2810 = _T_2678[495:488]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1746.4]
  assign _T_2811 = _T_2678[503:496]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1748.4]
  assign _T_2812 = _T_2678[511:504]; // @[NV_NVDLA_CSC_dl.scala 1071:37:@1750.4]
  assign _T_2814 = _T_896 != 3'h1; // @[NV_NVDLA_CSC_dl.scala 1074:59:@1752.4]
  assign _T_2815 = _T_2208 & _T_2814; // @[NV_NVDLA_CSC_dl.scala 1074:41:@1753.4]
  assign _T_2817 = _T_896 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1075:59:@1754.4]
  assign _T_2818 = _T_2211 & _T_2817; // @[NV_NVDLA_CSC_dl.scala 1075:41:@1755.4]
  assign _T_2821 = _T_2214 & _T_2817; // @[NV_NVDLA_CSC_dl.scala 1076:41:@1757.4]
  assign _GEN_149 = _T_2815 ? _T_2645 : {{256'd0}, _T_2611}; // @[NV_NVDLA_CSC_dl.scala 1078:24:@1758.4]
  assign _GEN_150 = _T_2818 ? _T_2611 : {{128'd0}, _T_2613}; // @[NV_NVDLA_CSC_dl.scala 1081:24:@1761.4]
  assign _GEN_151 = _T_2818 ? _T_2649 : {{384'd0}, _T_2617}; // @[NV_NVDLA_CSC_dl.scala 1081:24:@1761.4]
  assign _GEN_154 = _T_2821 ? _T_2653 : {{384'd0}, _T_2621}; // @[NV_NVDLA_CSC_dl.scala 1085:24:@1765.4]
  assign _T_2827 = 319'hffffffffffffffff << _T_2285; // @[NV_NVDLA_CSC_dl.scala 1094:56:@1771.4]
  assign _T_2828 = _T_2827[63:0]; // @[NV_NVDLA_CSC_dl.scala 1094:73:@1772.4]
  assign _T_2829 = ~ _T_2828; // @[NV_NVDLA_CSC_dl.scala 1094:24:@1773.4]
  assign _T_2831 = _T_2286 >= 2'h1; // @[NV_NVDLA_CSC_dl.scala 1096:51:@1774.4]
  assign _T_2838 = _T_2831 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl.scala 1096:32:@1776.4]
  assign _T_2840 = _T_2286 >= 2'h2; // @[NV_NVDLA_CSC_dl.scala 1097:51:@1777.4]
  assign _T_2847 = _T_2840 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl.scala 1097:32:@1779.4]
  assign _T_2849 = _T_2286 == 2'h3; // @[NV_NVDLA_CSC_dl.scala 1098:51:@1780.4]
  assign _T_2856 = _T_2849 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl.scala 1098:32:@1782.4]
  assign _T_2857 = _T_2838[31:0]; // @[NV_NVDLA_CSC_dl.scala 1100:57:@1783.4]
  assign _T_2863 = {_T_2857,32'hffffffff}; // @[Cat.scala 30:58:@1785.4]
  assign _T_2864 = _T_2856[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:57:@1786.4]
  assign _T_2865 = _T_2847[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:106:@1787.4]
  assign _T_2866 = _T_2838[15:0]; // @[NV_NVDLA_CSC_dl.scala 1101:155:@1788.4]
  assign _T_2874 = {_T_2864,_T_2865,_T_2866,16'hffff}; // @[Cat.scala 30:58:@1792.4]
  assign _T_2876 = _T_902 == 3'h4; // @[NV_NVDLA_CSC_dl.scala 1103:43:@1793.4]
  assign _T_2877 = _T_2829[15:0]; // @[NV_NVDLA_CSC_dl.scala 1103:89:@1794.4]
  assign _T_2879 = {_T_2877,_T_2877,_T_2877,_T_2877}; // @[Cat.scala 30:58:@1796.4]
  assign _T_2880 = _T_2879 & _T_2874; // @[NV_NVDLA_CSC_dl.scala 1103:116:@1797.4]
  assign _T_2882 = _T_902 == 3'h2; // @[NV_NVDLA_CSC_dl.scala 1104:43:@1798.4]
  assign _T_2883 = _T_2829[31:0]; // @[NV_NVDLA_CSC_dl.scala 1104:89:@1799.4]
  assign _T_2884 = {_T_2883,_T_2883}; // @[Cat.scala 30:58:@1800.4]
  assign _T_2885 = _T_2884 & _T_2863; // @[NV_NVDLA_CSC_dl.scala 1104:116:@1801.4]
  assign _T_2886 = _T_2882 ? _T_2885 : _T_2829; // @[NV_NVDLA_CSC_dl.scala 1104:26:@1802.4]
  assign _T_2887 = _T_2876 ? _T_2880 : _T_2886; // @[NV_NVDLA_CSC_dl.scala 1103:26:@1803.4]
  assign _T_2888 = _T_831[33]; // @[NV_NVDLA_CSC_dl.scala 1108:35:@1804.4]
  assign _T_2889_0 = _T_2888 ? _T_2749 : _T_2546; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_1 = _T_2888 ? _T_2750 : _T_2547; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_2 = _T_2888 ? _T_2751 : _T_2548; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_3 = _T_2888 ? _T_2752 : _T_2549; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_4 = _T_2888 ? _T_2753 : _T_2550; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_5 = _T_2888 ? _T_2754 : _T_2551; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_6 = _T_2888 ? _T_2755 : _T_2552; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_7 = _T_2888 ? _T_2756 : _T_2553; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_8 = _T_2888 ? _T_2757 : _T_2554; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_9 = _T_2888 ? _T_2758 : _T_2555; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_10 = _T_2888 ? _T_2759 : _T_2556; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_11 = _T_2888 ? _T_2760 : _T_2557; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_12 = _T_2888 ? _T_2761 : _T_2558; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_13 = _T_2888 ? _T_2762 : _T_2559; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_14 = _T_2888 ? _T_2763 : _T_2560; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_15 = _T_2888 ? _T_2764 : _T_2561; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_16 = _T_2888 ? _T_2765 : _T_2562; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_17 = _T_2888 ? _T_2766 : _T_2563; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_18 = _T_2888 ? _T_2767 : _T_2564; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_19 = _T_2888 ? _T_2768 : _T_2565; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_20 = _T_2888 ? _T_2769 : _T_2566; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_21 = _T_2888 ? _T_2770 : _T_2567; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_22 = _T_2888 ? _T_2771 : _T_2568; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_23 = _T_2888 ? _T_2772 : _T_2569; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_24 = _T_2888 ? _T_2773 : _T_2570; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_25 = _T_2888 ? _T_2774 : _T_2571; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_26 = _T_2888 ? _T_2775 : _T_2572; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_27 = _T_2888 ? _T_2776 : _T_2573; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_28 = _T_2888 ? _T_2777 : _T_2574; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_29 = _T_2888 ? _T_2778 : _T_2575; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_30 = _T_2888 ? _T_2779 : _T_2576; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_31 = _T_2888 ? _T_2780 : _T_2577; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_32 = _T_2888 ? _T_2781 : _T_2578; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_33 = _T_2888 ? _T_2782 : _T_2579; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_34 = _T_2888 ? _T_2783 : _T_2580; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_35 = _T_2888 ? _T_2784 : _T_2581; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_36 = _T_2888 ? _T_2785 : _T_2582; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_37 = _T_2888 ? _T_2786 : _T_2583; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_38 = _T_2888 ? _T_2787 : _T_2584; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_39 = _T_2888 ? _T_2788 : _T_2585; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_40 = _T_2888 ? _T_2789 : _T_2586; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_41 = _T_2888 ? _T_2790 : _T_2587; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_42 = _T_2888 ? _T_2791 : _T_2588; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_43 = _T_2888 ? _T_2792 : _T_2589; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_44 = _T_2888 ? _T_2793 : _T_2590; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_45 = _T_2888 ? _T_2794 : _T_2591; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_46 = _T_2888 ? _T_2795 : _T_2592; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_47 = _T_2888 ? _T_2796 : _T_2593; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_48 = _T_2888 ? _T_2797 : _T_2594; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_49 = _T_2888 ? _T_2798 : _T_2595; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_50 = _T_2888 ? _T_2799 : _T_2596; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_51 = _T_2888 ? _T_2800 : _T_2597; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_52 = _T_2888 ? _T_2801 : _T_2598; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_53 = _T_2888 ? _T_2802 : _T_2599; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_54 = _T_2888 ? _T_2803 : _T_2600; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_55 = _T_2888 ? _T_2804 : _T_2601; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_56 = _T_2888 ? _T_2805 : _T_2602; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_57 = _T_2888 ? _T_2806 : _T_2603; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_58 = _T_2888 ? _T_2807 : _T_2604; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_59 = _T_2888 ? _T_2808 : _T_2605; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_60 = _T_2888 ? _T_2809 : _T_2606; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_61 = _T_2888 ? _T_2810 : _T_2607; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_62 = _T_2888 ? _T_2811 : _T_2608; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_2889_63 = _T_2888 ? _T_2812 : _T_2609; // @[NV_NVDLA_CSC_dl.scala 1108:25:@1805.4]
  assign _T_3022 = _T_2889_0 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1806.4]
  assign _T_3024 = _T_2889_1 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1807.4]
  assign _T_3026 = _T_2889_2 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1808.4]
  assign _T_3028 = _T_2889_3 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1809.4]
  assign _T_3030 = _T_2889_4 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1810.4]
  assign _T_3032 = _T_2889_5 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1811.4]
  assign _T_3034 = _T_2889_6 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1812.4]
  assign _T_3036 = _T_2889_7 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1813.4]
  assign _T_3038 = _T_2889_8 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1814.4]
  assign _T_3040 = _T_2889_9 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1815.4]
  assign _T_3042 = _T_2889_10 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1816.4]
  assign _T_3044 = _T_2889_11 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1817.4]
  assign _T_3046 = _T_2889_12 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1818.4]
  assign _T_3048 = _T_2889_13 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1819.4]
  assign _T_3050 = _T_2889_14 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1820.4]
  assign _T_3052 = _T_2889_15 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1821.4]
  assign _T_3054 = _T_2889_16 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1822.4]
  assign _T_3056 = _T_2889_17 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1823.4]
  assign _T_3058 = _T_2889_18 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1824.4]
  assign _T_3060 = _T_2889_19 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1825.4]
  assign _T_3062 = _T_2889_20 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1826.4]
  assign _T_3064 = _T_2889_21 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1827.4]
  assign _T_3066 = _T_2889_22 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1828.4]
  assign _T_3068 = _T_2889_23 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1829.4]
  assign _T_3070 = _T_2889_24 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1830.4]
  assign _T_3072 = _T_2889_25 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1831.4]
  assign _T_3074 = _T_2889_26 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1832.4]
  assign _T_3076 = _T_2889_27 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1833.4]
  assign _T_3078 = _T_2889_28 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1834.4]
  assign _T_3080 = _T_2889_29 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1835.4]
  assign _T_3082 = _T_2889_30 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1836.4]
  assign _T_3084 = _T_2889_31 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1837.4]
  assign _T_3086 = _T_2889_32 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1838.4]
  assign _T_3088 = _T_2889_33 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1839.4]
  assign _T_3090 = _T_2889_34 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1840.4]
  assign _T_3092 = _T_2889_35 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1841.4]
  assign _T_3094 = _T_2889_36 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1842.4]
  assign _T_3096 = _T_2889_37 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1843.4]
  assign _T_3098 = _T_2889_38 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1844.4]
  assign _T_3100 = _T_2889_39 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1845.4]
  assign _T_3102 = _T_2889_40 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1846.4]
  assign _T_3104 = _T_2889_41 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1847.4]
  assign _T_3106 = _T_2889_42 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1848.4]
  assign _T_3108 = _T_2889_43 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1849.4]
  assign _T_3110 = _T_2889_44 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1850.4]
  assign _T_3112 = _T_2889_45 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1851.4]
  assign _T_3114 = _T_2889_46 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1852.4]
  assign _T_3116 = _T_2889_47 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1853.4]
  assign _T_3118 = _T_2889_48 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1854.4]
  assign _T_3120 = _T_2889_49 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1855.4]
  assign _T_3122 = _T_2889_50 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1856.4]
  assign _T_3124 = _T_2889_51 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1857.4]
  assign _T_3126 = _T_2889_52 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1858.4]
  assign _T_3128 = _T_2889_53 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1859.4]
  assign _T_3130 = _T_2889_54 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1860.4]
  assign _T_3132 = _T_2889_55 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1861.4]
  assign _T_3134 = _T_2889_56 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1862.4]
  assign _T_3136 = _T_2889_57 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1863.4]
  assign _T_3138 = _T_2889_58 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1864.4]
  assign _T_3140 = _T_2889_59 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1865.4]
  assign _T_3142 = _T_2889_60 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1866.4]
  assign _T_3144 = _T_2889_61 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1867.4]
  assign _T_3146 = _T_2889_62 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1868.4]
  assign _T_3148 = _T_2889_63 != 8'h0; // @[NV_NVDLA_CSC_dl.scala 1109:97:@1869.4]
  assign _T_3219 = _T_2887[0]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1935.4]
  assign _T_3220 = _T_3219 & _T_3022; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1936.4]
  assign _T_3221 = _T_2887[1]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1937.4]
  assign _T_3222 = _T_3221 & _T_3024; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1938.4]
  assign _T_3223 = _T_2887[2]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1939.4]
  assign _T_3224 = _T_3223 & _T_3026; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1940.4]
  assign _T_3225 = _T_2887[3]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1941.4]
  assign _T_3226 = _T_3225 & _T_3028; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1942.4]
  assign _T_3227 = _T_2887[4]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1943.4]
  assign _T_3228 = _T_3227 & _T_3030; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1944.4]
  assign _T_3229 = _T_2887[5]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1945.4]
  assign _T_3230 = _T_3229 & _T_3032; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1946.4]
  assign _T_3231 = _T_2887[6]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1947.4]
  assign _T_3232 = _T_3231 & _T_3034; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1948.4]
  assign _T_3233 = _T_2887[7]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1949.4]
  assign _T_3234 = _T_3233 & _T_3036; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1950.4]
  assign _T_3235 = _T_2887[8]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1951.4]
  assign _T_3236 = _T_3235 & _T_3038; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1952.4]
  assign _T_3237 = _T_2887[9]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1953.4]
  assign _T_3238 = _T_3237 & _T_3040; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1954.4]
  assign _T_3239 = _T_2887[10]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1955.4]
  assign _T_3240 = _T_3239 & _T_3042; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1956.4]
  assign _T_3241 = _T_2887[11]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1957.4]
  assign _T_3242 = _T_3241 & _T_3044; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1958.4]
  assign _T_3243 = _T_2887[12]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1959.4]
  assign _T_3244 = _T_3243 & _T_3046; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1960.4]
  assign _T_3245 = _T_2887[13]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1961.4]
  assign _T_3246 = _T_3245 & _T_3048; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1962.4]
  assign _T_3247 = _T_2887[14]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1963.4]
  assign _T_3248 = _T_3247 & _T_3050; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1964.4]
  assign _T_3249 = _T_2887[15]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1965.4]
  assign _T_3250 = _T_3249 & _T_3052; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1966.4]
  assign _T_3251 = _T_2887[16]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1967.4]
  assign _T_3252 = _T_3251 & _T_3054; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1968.4]
  assign _T_3253 = _T_2887[17]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1969.4]
  assign _T_3254 = _T_3253 & _T_3056; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1970.4]
  assign _T_3255 = _T_2887[18]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1971.4]
  assign _T_3256 = _T_3255 & _T_3058; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1972.4]
  assign _T_3257 = _T_2887[19]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1973.4]
  assign _T_3258 = _T_3257 & _T_3060; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1974.4]
  assign _T_3259 = _T_2887[20]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1975.4]
  assign _T_3260 = _T_3259 & _T_3062; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1976.4]
  assign _T_3261 = _T_2887[21]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1977.4]
  assign _T_3262 = _T_3261 & _T_3064; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1978.4]
  assign _T_3263 = _T_2887[22]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1979.4]
  assign _T_3264 = _T_3263 & _T_3066; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1980.4]
  assign _T_3265 = _T_2887[23]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1981.4]
  assign _T_3266 = _T_3265 & _T_3068; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1982.4]
  assign _T_3267 = _T_2887[24]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1983.4]
  assign _T_3268 = _T_3267 & _T_3070; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1984.4]
  assign _T_3269 = _T_2887[25]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1985.4]
  assign _T_3270 = _T_3269 & _T_3072; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1986.4]
  assign _T_3271 = _T_2887[26]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1987.4]
  assign _T_3272 = _T_3271 & _T_3074; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1988.4]
  assign _T_3273 = _T_2887[27]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1989.4]
  assign _T_3274 = _T_3273 & _T_3076; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1990.4]
  assign _T_3275 = _T_2887[28]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1991.4]
  assign _T_3276 = _T_3275 & _T_3078; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1992.4]
  assign _T_3277 = _T_2887[29]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1993.4]
  assign _T_3278 = _T_3277 & _T_3080; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1994.4]
  assign _T_3279 = _T_2887[30]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1995.4]
  assign _T_3280 = _T_3279 & _T_3082; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1996.4]
  assign _T_3281 = _T_2887[31]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1997.4]
  assign _T_3282 = _T_3281 & _T_3084; // @[NV_NVDLA_CSC_dl.scala 1110:83:@1998.4]
  assign _T_3283 = _T_2887[32]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@1999.4]
  assign _T_3284 = _T_3283 & _T_3086; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2000.4]
  assign _T_3285 = _T_2887[33]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2001.4]
  assign _T_3286 = _T_3285 & _T_3088; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2002.4]
  assign _T_3287 = _T_2887[34]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2003.4]
  assign _T_3288 = _T_3287 & _T_3090; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2004.4]
  assign _T_3289 = _T_2887[35]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2005.4]
  assign _T_3290 = _T_3289 & _T_3092; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2006.4]
  assign _T_3291 = _T_2887[36]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2007.4]
  assign _T_3292 = _T_3291 & _T_3094; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2008.4]
  assign _T_3293 = _T_2887[37]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2009.4]
  assign _T_3294 = _T_3293 & _T_3096; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2010.4]
  assign _T_3295 = _T_2887[38]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2011.4]
  assign _T_3296 = _T_3295 & _T_3098; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2012.4]
  assign _T_3297 = _T_2887[39]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2013.4]
  assign _T_3298 = _T_3297 & _T_3100; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2014.4]
  assign _T_3299 = _T_2887[40]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2015.4]
  assign _T_3300 = _T_3299 & _T_3102; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2016.4]
  assign _T_3301 = _T_2887[41]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2017.4]
  assign _T_3302 = _T_3301 & _T_3104; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2018.4]
  assign _T_3303 = _T_2887[42]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2019.4]
  assign _T_3304 = _T_3303 & _T_3106; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2020.4]
  assign _T_3305 = _T_2887[43]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2021.4]
  assign _T_3306 = _T_3305 & _T_3108; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2022.4]
  assign _T_3307 = _T_2887[44]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2023.4]
  assign _T_3308 = _T_3307 & _T_3110; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2024.4]
  assign _T_3309 = _T_2887[45]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2025.4]
  assign _T_3310 = _T_3309 & _T_3112; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2026.4]
  assign _T_3311 = _T_2887[46]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2027.4]
  assign _T_3312 = _T_3311 & _T_3114; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2028.4]
  assign _T_3313 = _T_2887[47]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2029.4]
  assign _T_3314 = _T_3313 & _T_3116; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2030.4]
  assign _T_3315 = _T_2887[48]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2031.4]
  assign _T_3316 = _T_3315 & _T_3118; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2032.4]
  assign _T_3317 = _T_2887[49]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2033.4]
  assign _T_3318 = _T_3317 & _T_3120; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2034.4]
  assign _T_3319 = _T_2887[50]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2035.4]
  assign _T_3320 = _T_3319 & _T_3122; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2036.4]
  assign _T_3321 = _T_2887[51]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2037.4]
  assign _T_3322 = _T_3321 & _T_3124; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2038.4]
  assign _T_3323 = _T_2887[52]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2039.4]
  assign _T_3324 = _T_3323 & _T_3126; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2040.4]
  assign _T_3325 = _T_2887[53]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2041.4]
  assign _T_3326 = _T_3325 & _T_3128; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2042.4]
  assign _T_3327 = _T_2887[54]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2043.4]
  assign _T_3328 = _T_3327 & _T_3130; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2044.4]
  assign _T_3329 = _T_2887[55]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2045.4]
  assign _T_3330 = _T_3329 & _T_3132; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2046.4]
  assign _T_3331 = _T_2887[56]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2047.4]
  assign _T_3332 = _T_3331 & _T_3134; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2048.4]
  assign _T_3333 = _T_2887[57]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2049.4]
  assign _T_3334 = _T_3333 & _T_3136; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2050.4]
  assign _T_3335 = _T_2887[58]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2051.4]
  assign _T_3336 = _T_3335 & _T_3138; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2052.4]
  assign _T_3337 = _T_2887[59]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2053.4]
  assign _T_3338 = _T_3337 & _T_3140; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2054.4]
  assign _T_3339 = _T_2887[60]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2055.4]
  assign _T_3340 = _T_3339 & _T_3142; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2056.4]
  assign _T_3341 = _T_2887[61]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2057.4]
  assign _T_3342 = _T_3341 & _T_3144; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2058.4]
  assign _T_3343 = _T_2887[62]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2059.4]
  assign _T_3344 = _T_3343 & _T_3146; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2060.4]
  assign _T_3345 = _T_2887[63]; // @[NV_NVDLA_CSC_dl.scala 1110:80:@2061.4]
  assign _T_3346 = _T_3345 & _T_3148; // @[NV_NVDLA_CSC_dl.scala 1110:83:@2062.4]
  assign _GEN_156 = _T_2248 ? _T_3220 : _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_157 = _T_2248 ? _T_3222 : _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_158 = _T_2248 ? _T_3224 : _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_159 = _T_2248 ? _T_3226 : _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_160 = _T_2248 ? _T_3228 : _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_161 = _T_2248 ? _T_3230 : _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_162 = _T_2248 ? _T_3232 : _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_163 = _T_2248 ? _T_3234 : _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_164 = _T_2248 ? _T_3236 : _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_165 = _T_2248 ? _T_3238 : _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_166 = _T_2248 ? _T_3240 : _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_167 = _T_2248 ? _T_3242 : _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_168 = _T_2248 ? _T_3244 : _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_169 = _T_2248 ? _T_3246 : _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_170 = _T_2248 ? _T_3248 : _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_171 = _T_2248 ? _T_3250 : _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_172 = _T_2248 ? _T_3252 : _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_173 = _T_2248 ? _T_3254 : _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_174 = _T_2248 ? _T_3256 : _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_175 = _T_2248 ? _T_3258 : _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_176 = _T_2248 ? _T_3260 : _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_177 = _T_2248 ? _T_3262 : _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_178 = _T_2248 ? _T_3264 : _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_179 = _T_2248 ? _T_3266 : _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_180 = _T_2248 ? _T_3268 : _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_181 = _T_2248 ? _T_3270 : _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_182 = _T_2248 ? _T_3272 : _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_183 = _T_2248 ? _T_3274 : _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_184 = _T_2248 ? _T_3276 : _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_185 = _T_2248 ? _T_3278 : _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_186 = _T_2248 ? _T_3280 : _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_187 = _T_2248 ? _T_3282 : _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_188 = _T_2248 ? _T_3284 : _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_189 = _T_2248 ? _T_3286 : _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_190 = _T_2248 ? _T_3288 : _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_191 = _T_2248 ? _T_3290 : _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_192 = _T_2248 ? _T_3292 : _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_193 = _T_2248 ? _T_3294 : _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_194 = _T_2248 ? _T_3296 : _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_195 = _T_2248 ? _T_3298 : _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_196 = _T_2248 ? _T_3300 : _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_197 = _T_2248 ? _T_3302 : _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_198 = _T_2248 ? _T_3304 : _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_199 = _T_2248 ? _T_3306 : _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_200 = _T_2248 ? _T_3308 : _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_201 = _T_2248 ? _T_3310 : _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_202 = _T_2248 ? _T_3312 : _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_203 = _T_2248 ? _T_3314 : _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_204 = _T_2248 ? _T_3316 : _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_205 = _T_2248 ? _T_3318 : _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_206 = _T_2248 ? _T_3320 : _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_207 = _T_2248 ? _T_3322 : _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_208 = _T_2248 ? _T_3324 : _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_209 = _T_2248 ? _T_3326 : _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_210 = _T_2248 ? _T_3328 : _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_211 = _T_2248 ? _T_3330 : _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_212 = _T_2248 ? _T_3332 : _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_213 = _T_2248 ? _T_3334 : _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_214 = _T_2248 ? _T_3336 : _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_215 = _T_2248 ? _T_3338 : _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_216 = _T_2248 ? _T_3340 : _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_217 = _T_2248 ? _T_3342 : _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_218 = _T_2248 ? _T_3344 : _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _GEN_219 = _T_2248 ? _T_3346 : _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1133:30:@2201.4]
  assign _T_3956 = _T_2248 & _T_3220; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2267.4]
  assign _T_3957 = _T_2248 & _T_3222; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2271.4]
  assign _T_3958 = _T_2248 & _T_3224; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2275.4]
  assign _T_3959 = _T_2248 & _T_3226; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2279.4]
  assign _T_3960 = _T_2248 & _T_3228; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2283.4]
  assign _T_3961 = _T_2248 & _T_3230; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2287.4]
  assign _T_3962 = _T_2248 & _T_3232; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2291.4]
  assign _T_3963 = _T_2248 & _T_3234; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2295.4]
  assign _T_3964 = _T_2248 & _T_3236; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2299.4]
  assign _T_3965 = _T_2248 & _T_3238; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2303.4]
  assign _T_3966 = _T_2248 & _T_3240; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2307.4]
  assign _T_3967 = _T_2248 & _T_3242; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2311.4]
  assign _T_3968 = _T_2248 & _T_3244; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2315.4]
  assign _T_3969 = _T_2248 & _T_3246; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2319.4]
  assign _T_3970 = _T_2248 & _T_3248; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2323.4]
  assign _T_3971 = _T_2248 & _T_3250; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2327.4]
  assign _T_3972 = _T_2248 & _T_3252; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2331.4]
  assign _T_3973 = _T_2248 & _T_3254; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2335.4]
  assign _T_3974 = _T_2248 & _T_3256; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2339.4]
  assign _T_3975 = _T_2248 & _T_3258; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2343.4]
  assign _T_3976 = _T_2248 & _T_3260; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2347.4]
  assign _T_3977 = _T_2248 & _T_3262; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2351.4]
  assign _T_3978 = _T_2248 & _T_3264; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2355.4]
  assign _T_3979 = _T_2248 & _T_3266; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2359.4]
  assign _T_3980 = _T_2248 & _T_3268; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2363.4]
  assign _T_3981 = _T_2248 & _T_3270; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2367.4]
  assign _T_3982 = _T_2248 & _T_3272; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2371.4]
  assign _T_3983 = _T_2248 & _T_3274; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2375.4]
  assign _T_3984 = _T_2248 & _T_3276; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2379.4]
  assign _T_3985 = _T_2248 & _T_3278; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2383.4]
  assign _T_3986 = _T_2248 & _T_3280; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2387.4]
  assign _T_3987 = _T_2248 & _T_3282; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2391.4]
  assign _T_3988 = _T_2248 & _T_3284; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2395.4]
  assign _T_3989 = _T_2248 & _T_3286; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2399.4]
  assign _T_3990 = _T_2248 & _T_3288; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2403.4]
  assign _T_3991 = _T_2248 & _T_3290; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2407.4]
  assign _T_3992 = _T_2248 & _T_3292; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2411.4]
  assign _T_3993 = _T_2248 & _T_3294; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2415.4]
  assign _T_3994 = _T_2248 & _T_3296; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2419.4]
  assign _T_3995 = _T_2248 & _T_3298; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2423.4]
  assign _T_3996 = _T_2248 & _T_3300; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2427.4]
  assign _T_3997 = _T_2248 & _T_3302; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2431.4]
  assign _T_3998 = _T_2248 & _T_3304; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2435.4]
  assign _T_3999 = _T_2248 & _T_3306; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2439.4]
  assign _T_4000 = _T_2248 & _T_3308; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2443.4]
  assign _T_4001 = _T_2248 & _T_3310; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2447.4]
  assign _T_4002 = _T_2248 & _T_3312; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2451.4]
  assign _T_4003 = _T_2248 & _T_3314; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2455.4]
  assign _T_4004 = _T_2248 & _T_3316; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2459.4]
  assign _T_4005 = _T_2248 & _T_3318; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2463.4]
  assign _T_4006 = _T_2248 & _T_3320; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2467.4]
  assign _T_4007 = _T_2248 & _T_3322; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2471.4]
  assign _T_4008 = _T_2248 & _T_3324; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2475.4]
  assign _T_4009 = _T_2248 & _T_3326; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2479.4]
  assign _T_4010 = _T_2248 & _T_3328; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2483.4]
  assign _T_4011 = _T_2248 & _T_3330; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2487.4]
  assign _T_4012 = _T_2248 & _T_3332; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2491.4]
  assign _T_4013 = _T_2248 & _T_3334; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2495.4]
  assign _T_4014 = _T_2248 & _T_3336; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2499.4]
  assign _T_4015 = _T_2248 & _T_3338; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2503.4]
  assign _T_4016 = _T_2248 & _T_3340; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2507.4]
  assign _T_4017 = _T_2248 & _T_3342; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2511.4]
  assign _T_4018 = _T_2248 & _T_3344; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2515.4]
  assign _T_4019 = _T_2248 & _T_3346; // @[NV_NVDLA_CSC_dl.scala 1137:34:@2519.4]
  assign _T_4559 = ~ _T_3419; // @[NV_NVDLA_CSC_dl.scala 1151:24:@2592.4]
  assign _T_4694_0 = _T_4559 ? 1'h0 : _T_3689_0; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_1 = _T_4559 ? 1'h0 : _T_3689_1; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_2 = _T_4559 ? 1'h0 : _T_3689_2; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_3 = _T_4559 ? 1'h0 : _T_3689_3; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_4 = _T_4559 ? 1'h0 : _T_3689_4; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_5 = _T_4559 ? 1'h0 : _T_3689_5; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_6 = _T_4559 ? 1'h0 : _T_3689_6; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_7 = _T_4559 ? 1'h0 : _T_3689_7; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_8 = _T_4559 ? 1'h0 : _T_3689_8; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_9 = _T_4559 ? 1'h0 : _T_3689_9; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_10 = _T_4559 ? 1'h0 : _T_3689_10; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_11 = _T_4559 ? 1'h0 : _T_3689_11; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_12 = _T_4559 ? 1'h0 : _T_3689_12; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_13 = _T_4559 ? 1'h0 : _T_3689_13; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_14 = _T_4559 ? 1'h0 : _T_3689_14; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_15 = _T_4559 ? 1'h0 : _T_3689_15; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_16 = _T_4559 ? 1'h0 : _T_3689_16; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_17 = _T_4559 ? 1'h0 : _T_3689_17; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_18 = _T_4559 ? 1'h0 : _T_3689_18; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_19 = _T_4559 ? 1'h0 : _T_3689_19; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_20 = _T_4559 ? 1'h0 : _T_3689_20; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_21 = _T_4559 ? 1'h0 : _T_3689_21; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_22 = _T_4559 ? 1'h0 : _T_3689_22; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_23 = _T_4559 ? 1'h0 : _T_3689_23; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_24 = _T_4559 ? 1'h0 : _T_3689_24; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_25 = _T_4559 ? 1'h0 : _T_3689_25; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_26 = _T_4559 ? 1'h0 : _T_3689_26; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_27 = _T_4559 ? 1'h0 : _T_3689_27; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_28 = _T_4559 ? 1'h0 : _T_3689_28; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_29 = _T_4559 ? 1'h0 : _T_3689_29; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_30 = _T_4559 ? 1'h0 : _T_3689_30; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_31 = _T_4559 ? 1'h0 : _T_3689_31; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_32 = _T_4559 ? 1'h0 : _T_3689_32; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_33 = _T_4559 ? 1'h0 : _T_3689_33; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_34 = _T_4559 ? 1'h0 : _T_3689_34; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_35 = _T_4559 ? 1'h0 : _T_3689_35; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_36 = _T_4559 ? 1'h0 : _T_3689_36; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_37 = _T_4559 ? 1'h0 : _T_3689_37; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_38 = _T_4559 ? 1'h0 : _T_3689_38; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_39 = _T_4559 ? 1'h0 : _T_3689_39; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_40 = _T_4559 ? 1'h0 : _T_3689_40; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_41 = _T_4559 ? 1'h0 : _T_3689_41; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_42 = _T_4559 ? 1'h0 : _T_3689_42; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_43 = _T_4559 ? 1'h0 : _T_3689_43; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_44 = _T_4559 ? 1'h0 : _T_3689_44; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_45 = _T_4559 ? 1'h0 : _T_3689_45; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_46 = _T_4559 ? 1'h0 : _T_3689_46; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_47 = _T_4559 ? 1'h0 : _T_3689_47; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_48 = _T_4559 ? 1'h0 : _T_3689_48; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_49 = _T_4559 ? 1'h0 : _T_3689_49; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_50 = _T_4559 ? 1'h0 : _T_3689_50; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_51 = _T_4559 ? 1'h0 : _T_3689_51; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_52 = _T_4559 ? 1'h0 : _T_3689_52; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_53 = _T_4559 ? 1'h0 : _T_3689_53; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_54 = _T_4559 ? 1'h0 : _T_3689_54; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_55 = _T_4559 ? 1'h0 : _T_3689_55; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_56 = _T_4559 ? 1'h0 : _T_3689_56; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_57 = _T_4559 ? 1'h0 : _T_3689_57; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_58 = _T_4559 ? 1'h0 : _T_3689_58; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_59 = _T_4559 ? 1'h0 : _T_3689_59; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_60 = _T_4559 ? 1'h0 : _T_3689_60; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_61 = _T_4559 ? 1'h0 : _T_3689_61; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_62 = _T_4559 ? 1'h0 : _T_3689_62; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4694_63 = _T_4559 ? 1'h0 : _T_3689_63; // @[NV_NVDLA_CSC_dl.scala 1151:23:@2658.4]
  assign _T_4826 = _T_3419 | _T_4022; // @[NV_NVDLA_CSC_dl.scala 1155:19:@2660.4]
  assign _GEN_284 = _T_4826 ? _T_4694_0 : _T_4289_0; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_285 = _T_4826 ? _T_4694_1 : _T_4289_1; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_286 = _T_4826 ? _T_4694_2 : _T_4289_2; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_287 = _T_4826 ? _T_4694_3 : _T_4289_3; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_288 = _T_4826 ? _T_4694_4 : _T_4289_4; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_289 = _T_4826 ? _T_4694_5 : _T_4289_5; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_290 = _T_4826 ? _T_4694_6 : _T_4289_6; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_291 = _T_4826 ? _T_4694_7 : _T_4289_7; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_292 = _T_4826 ? _T_4694_8 : _T_4289_8; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_293 = _T_4826 ? _T_4694_9 : _T_4289_9; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_294 = _T_4826 ? _T_4694_10 : _T_4289_10; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_295 = _T_4826 ? _T_4694_11 : _T_4289_11; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_296 = _T_4826 ? _T_4694_12 : _T_4289_12; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_297 = _T_4826 ? _T_4694_13 : _T_4289_13; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_298 = _T_4826 ? _T_4694_14 : _T_4289_14; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_299 = _T_4826 ? _T_4694_15 : _T_4289_15; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_300 = _T_4826 ? _T_4694_16 : _T_4289_16; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_301 = _T_4826 ? _T_4694_17 : _T_4289_17; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_302 = _T_4826 ? _T_4694_18 : _T_4289_18; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_303 = _T_4826 ? _T_4694_19 : _T_4289_19; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_304 = _T_4826 ? _T_4694_20 : _T_4289_20; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_305 = _T_4826 ? _T_4694_21 : _T_4289_21; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_306 = _T_4826 ? _T_4694_22 : _T_4289_22; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_307 = _T_4826 ? _T_4694_23 : _T_4289_23; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_308 = _T_4826 ? _T_4694_24 : _T_4289_24; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_309 = _T_4826 ? _T_4694_25 : _T_4289_25; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_310 = _T_4826 ? _T_4694_26 : _T_4289_26; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_311 = _T_4826 ? _T_4694_27 : _T_4289_27; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_312 = _T_4826 ? _T_4694_28 : _T_4289_28; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_313 = _T_4826 ? _T_4694_29 : _T_4289_29; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_314 = _T_4826 ? _T_4694_30 : _T_4289_30; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_315 = _T_4826 ? _T_4694_31 : _T_4289_31; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_316 = _T_4826 ? _T_4694_32 : _T_4289_32; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_317 = _T_4826 ? _T_4694_33 : _T_4289_33; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_318 = _T_4826 ? _T_4694_34 : _T_4289_34; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_319 = _T_4826 ? _T_4694_35 : _T_4289_35; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_320 = _T_4826 ? _T_4694_36 : _T_4289_36; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_321 = _T_4826 ? _T_4694_37 : _T_4289_37; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_322 = _T_4826 ? _T_4694_38 : _T_4289_38; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_323 = _T_4826 ? _T_4694_39 : _T_4289_39; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_324 = _T_4826 ? _T_4694_40 : _T_4289_40; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_325 = _T_4826 ? _T_4694_41 : _T_4289_41; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_326 = _T_4826 ? _T_4694_42 : _T_4289_42; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_327 = _T_4826 ? _T_4694_43 : _T_4289_43; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_328 = _T_4826 ? _T_4694_44 : _T_4289_44; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_329 = _T_4826 ? _T_4694_45 : _T_4289_45; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_330 = _T_4826 ? _T_4694_46 : _T_4289_46; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_331 = _T_4826 ? _T_4694_47 : _T_4289_47; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_332 = _T_4826 ? _T_4694_48 : _T_4289_48; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_333 = _T_4826 ? _T_4694_49 : _T_4289_49; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_334 = _T_4826 ? _T_4694_50 : _T_4289_50; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_335 = _T_4826 ? _T_4694_51 : _T_4289_51; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_336 = _T_4826 ? _T_4694_52 : _T_4289_52; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_337 = _T_4826 ? _T_4694_53 : _T_4289_53; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_338 = _T_4826 ? _T_4694_54 : _T_4289_54; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_339 = _T_4826 ? _T_4694_55 : _T_4289_55; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_340 = _T_4826 ? _T_4694_56 : _T_4289_56; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_341 = _T_4826 ? _T_4694_57 : _T_4289_57; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_342 = _T_4826 ? _T_4694_58 : _T_4289_58; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_343 = _T_4826 ? _T_4694_59 : _T_4289_59; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_344 = _T_4826 ? _T_4694_60 : _T_4289_60; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_345 = _T_4826 ? _T_4694_61 : _T_4289_61; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_346 = _T_4826 ? _T_4694_62 : _T_4289_62; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_347 = _T_4826 ? _T_4694_63 : _T_4289_63; // @[NV_NVDLA_CSC_dl.scala 1155:33:@2661.4]
  assign _GEN_348 = _T_3419 ? {{8'd0}, _T_3419} : _T_4488; // @[NV_NVDLA_CSC_dl.scala 1158:19:@2727.4]
  assign _T_4830 = ~ _T_4022; // @[NV_NVDLA_CSC_dl.scala 1172:27:@2924.4]
  assign _T_4832 = _T_4830 ? 9'h0 : _T_4488; // @[NV_NVDLA_CSC_dl.scala 1172:26:@2925.4]
  assign _T_4840 = _T_4022 | _T_4829; // @[NV_NVDLA_CSC_dl.scala 1176:85:@2932.4]
  assign _GEN_413 = _T_4840 ? _T_4832 : _T_4842; // @[Reg.scala 20:19:@2934.4]
  assign _GEN_414 = _T_4840 ? _T_4832 : _T_4846; // @[Reg.scala 20:19:@2940.4]
  assign _GEN_415 = _T_4840 ? _T_4289_0 : _T_5114_0; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_416 = _T_4840 ? _T_4289_1 : _T_5114_1; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_417 = _T_4840 ? _T_4289_2 : _T_5114_2; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_418 = _T_4840 ? _T_4289_3 : _T_5114_3; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_419 = _T_4840 ? _T_4289_4 : _T_5114_4; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_420 = _T_4840 ? _T_4289_5 : _T_5114_5; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_421 = _T_4840 ? _T_4289_6 : _T_5114_6; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_422 = _T_4840 ? _T_4289_7 : _T_5114_7; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_423 = _T_4840 ? _T_4289_8 : _T_5114_8; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_424 = _T_4840 ? _T_4289_9 : _T_5114_9; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_425 = _T_4840 ? _T_4289_10 : _T_5114_10; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_426 = _T_4840 ? _T_4289_11 : _T_5114_11; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_427 = _T_4840 ? _T_4289_12 : _T_5114_12; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_428 = _T_4840 ? _T_4289_13 : _T_5114_13; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_429 = _T_4840 ? _T_4289_14 : _T_5114_14; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_430 = _T_4840 ? _T_4289_15 : _T_5114_15; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_431 = _T_4840 ? _T_4289_16 : _T_5114_16; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_432 = _T_4840 ? _T_4289_17 : _T_5114_17; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_433 = _T_4840 ? _T_4289_18 : _T_5114_18; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_434 = _T_4840 ? _T_4289_19 : _T_5114_19; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_435 = _T_4840 ? _T_4289_20 : _T_5114_20; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_436 = _T_4840 ? _T_4289_21 : _T_5114_21; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_437 = _T_4840 ? _T_4289_22 : _T_5114_22; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_438 = _T_4840 ? _T_4289_23 : _T_5114_23; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_439 = _T_4840 ? _T_4289_24 : _T_5114_24; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_440 = _T_4840 ? _T_4289_25 : _T_5114_25; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_441 = _T_4840 ? _T_4289_26 : _T_5114_26; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_442 = _T_4840 ? _T_4289_27 : _T_5114_27; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_443 = _T_4840 ? _T_4289_28 : _T_5114_28; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_444 = _T_4840 ? _T_4289_29 : _T_5114_29; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_445 = _T_4840 ? _T_4289_30 : _T_5114_30; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_446 = _T_4840 ? _T_4289_31 : _T_5114_31; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_447 = _T_4840 ? _T_4289_32 : _T_5114_32; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_448 = _T_4840 ? _T_4289_33 : _T_5114_33; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_449 = _T_4840 ? _T_4289_34 : _T_5114_34; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_450 = _T_4840 ? _T_4289_35 : _T_5114_35; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_451 = _T_4840 ? _T_4289_36 : _T_5114_36; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_452 = _T_4840 ? _T_4289_37 : _T_5114_37; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_453 = _T_4840 ? _T_4289_38 : _T_5114_38; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_454 = _T_4840 ? _T_4289_39 : _T_5114_39; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_455 = _T_4840 ? _T_4289_40 : _T_5114_40; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_456 = _T_4840 ? _T_4289_41 : _T_5114_41; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_457 = _T_4840 ? _T_4289_42 : _T_5114_42; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_458 = _T_4840 ? _T_4289_43 : _T_5114_43; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_459 = _T_4840 ? _T_4289_44 : _T_5114_44; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_460 = _T_4840 ? _T_4289_45 : _T_5114_45; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_461 = _T_4840 ? _T_4289_46 : _T_5114_46; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_462 = _T_4840 ? _T_4289_47 : _T_5114_47; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_463 = _T_4840 ? _T_4289_48 : _T_5114_48; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_464 = _T_4840 ? _T_4289_49 : _T_5114_49; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_465 = _T_4840 ? _T_4289_50 : _T_5114_50; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_466 = _T_4840 ? _T_4289_51 : _T_5114_51; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_467 = _T_4840 ? _T_4289_52 : _T_5114_52; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_468 = _T_4840 ? _T_4289_53 : _T_5114_53; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_469 = _T_4840 ? _T_4289_54 : _T_5114_54; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_470 = _T_4840 ? _T_4289_55 : _T_5114_55; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_471 = _T_4840 ? _T_4289_56 : _T_5114_56; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_472 = _T_4840 ? _T_4289_57 : _T_5114_57; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_473 = _T_4840 ? _T_4289_58 : _T_5114_58; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_474 = _T_4840 ? _T_4289_59 : _T_5114_59; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_475 = _T_4840 ? _T_4289_60 : _T_5114_60; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_476 = _T_4840 ? _T_4289_61 : _T_5114_61; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_477 = _T_4840 ? _T_4289_62 : _T_5114_62; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_478 = _T_4840 ? _T_4289_63 : _T_5114_63; // @[Reg.scala 20:19:@3011.4]
  assign _GEN_479 = _T_4840 ? _T_4289_0 : _T_5578_0; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_480 = _T_4840 ? _T_4289_1 : _T_5578_1; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_481 = _T_4840 ? _T_4289_2 : _T_5578_2; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_482 = _T_4840 ? _T_4289_3 : _T_5578_3; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_483 = _T_4840 ? _T_4289_4 : _T_5578_4; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_484 = _T_4840 ? _T_4289_5 : _T_5578_5; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_485 = _T_4840 ? _T_4289_6 : _T_5578_6; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_486 = _T_4840 ? _T_4289_7 : _T_5578_7; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_487 = _T_4840 ? _T_4289_8 : _T_5578_8; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_488 = _T_4840 ? _T_4289_9 : _T_5578_9; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_489 = _T_4840 ? _T_4289_10 : _T_5578_10; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_490 = _T_4840 ? _T_4289_11 : _T_5578_11; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_491 = _T_4840 ? _T_4289_12 : _T_5578_12; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_492 = _T_4840 ? _T_4289_13 : _T_5578_13; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_493 = _T_4840 ? _T_4289_14 : _T_5578_14; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_494 = _T_4840 ? _T_4289_15 : _T_5578_15; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_495 = _T_4840 ? _T_4289_16 : _T_5578_16; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_496 = _T_4840 ? _T_4289_17 : _T_5578_17; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_497 = _T_4840 ? _T_4289_18 : _T_5578_18; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_498 = _T_4840 ? _T_4289_19 : _T_5578_19; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_499 = _T_4840 ? _T_4289_20 : _T_5578_20; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_500 = _T_4840 ? _T_4289_21 : _T_5578_21; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_501 = _T_4840 ? _T_4289_22 : _T_5578_22; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_502 = _T_4840 ? _T_4289_23 : _T_5578_23; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_503 = _T_4840 ? _T_4289_24 : _T_5578_24; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_504 = _T_4840 ? _T_4289_25 : _T_5578_25; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_505 = _T_4840 ? _T_4289_26 : _T_5578_26; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_506 = _T_4840 ? _T_4289_27 : _T_5578_27; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_507 = _T_4840 ? _T_4289_28 : _T_5578_28; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_508 = _T_4840 ? _T_4289_29 : _T_5578_29; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_509 = _T_4840 ? _T_4289_30 : _T_5578_30; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_510 = _T_4840 ? _T_4289_31 : _T_5578_31; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_511 = _T_4840 ? _T_4289_32 : _T_5578_32; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_512 = _T_4840 ? _T_4289_33 : _T_5578_33; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_513 = _T_4840 ? _T_4289_34 : _T_5578_34; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_514 = _T_4840 ? _T_4289_35 : _T_5578_35; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_515 = _T_4840 ? _T_4289_36 : _T_5578_36; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_516 = _T_4840 ? _T_4289_37 : _T_5578_37; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_517 = _T_4840 ? _T_4289_38 : _T_5578_38; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_518 = _T_4840 ? _T_4289_39 : _T_5578_39; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_519 = _T_4840 ? _T_4289_40 : _T_5578_40; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_520 = _T_4840 ? _T_4289_41 : _T_5578_41; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_521 = _T_4840 ? _T_4289_42 : _T_5578_42; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_522 = _T_4840 ? _T_4289_43 : _T_5578_43; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_523 = _T_4840 ? _T_4289_44 : _T_5578_44; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_524 = _T_4840 ? _T_4289_45 : _T_5578_45; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_525 = _T_4840 ? _T_4289_46 : _T_5578_46; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_526 = _T_4840 ? _T_4289_47 : _T_5578_47; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_527 = _T_4840 ? _T_4289_48 : _T_5578_48; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_528 = _T_4840 ? _T_4289_49 : _T_5578_49; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_529 = _T_4840 ? _T_4289_50 : _T_5578_50; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_530 = _T_4840 ? _T_4289_51 : _T_5578_51; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_531 = _T_4840 ? _T_4289_52 : _T_5578_52; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_532 = _T_4840 ? _T_4289_53 : _T_5578_53; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_533 = _T_4840 ? _T_4289_54 : _T_5578_54; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_534 = _T_4840 ? _T_4289_55 : _T_5578_55; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_535 = _T_4840 ? _T_4289_56 : _T_5578_56; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_536 = _T_4840 ? _T_4289_57 : _T_5578_57; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_537 = _T_4840 ? _T_4289_58 : _T_5578_58; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_538 = _T_4840 ? _T_4289_59 : _T_5578_59; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_539 = _T_4840 ? _T_4289_60 : _T_5578_60; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_540 = _T_4840 ? _T_4289_61 : _T_5578_61; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_541 = _T_4840 ? _T_4289_62 : _T_5578_62; // @[Reg.scala 20:19:@3208.4]
  assign _GEN_542 = _T_4840 ? _T_4289_63 : _T_5578_63; // @[Reg.scala 20:19:@3208.4]
  assign io_sc2cdma_dat_updt_valid = _T_1166; // @[NV_NVDLA_CSC_dl.scala 308:27:@325.4]
  assign io_sc2cdma_dat_updt_bits_entries = _T_1172; // @[NV_NVDLA_CSC_dl.scala 310:34:@335.4]
  assign io_sc2cdma_dat_updt_bits_slices = _T_1169; // @[NV_NVDLA_CSC_dl.scala 309:33:@330.4]
  assign io_sc2buf_dat_rd_addr_valid = _T_1778; // @[NV_NVDLA_CSC_dl.scala 725:29:@932.4]
  assign io_sc2buf_dat_rd_addr_bits = _T_1785[12:0]; // @[NV_NVDLA_CSC_dl.scala 726:28:@933.4]
  assign io_sc2mac_dat_a_valid = _T_4835; // @[NV_NVDLA_CSC_dl.scala 1174:23:@2928.4]
  assign io_sc2mac_dat_a_bits_mask_0 = _T_5114_0; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3077.4]
  assign io_sc2mac_dat_a_bits_mask_1 = _T_5114_1; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3078.4]
  assign io_sc2mac_dat_a_bits_mask_2 = _T_5114_2; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3079.4]
  assign io_sc2mac_dat_a_bits_mask_3 = _T_5114_3; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3080.4]
  assign io_sc2mac_dat_a_bits_mask_4 = _T_5114_4; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3081.4]
  assign io_sc2mac_dat_a_bits_mask_5 = _T_5114_5; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3082.4]
  assign io_sc2mac_dat_a_bits_mask_6 = _T_5114_6; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3083.4]
  assign io_sc2mac_dat_a_bits_mask_7 = _T_5114_7; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3084.4]
  assign io_sc2mac_dat_a_bits_mask_8 = _T_5114_8; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3085.4]
  assign io_sc2mac_dat_a_bits_mask_9 = _T_5114_9; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3086.4]
  assign io_sc2mac_dat_a_bits_mask_10 = _T_5114_10; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3087.4]
  assign io_sc2mac_dat_a_bits_mask_11 = _T_5114_11; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3088.4]
  assign io_sc2mac_dat_a_bits_mask_12 = _T_5114_12; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3089.4]
  assign io_sc2mac_dat_a_bits_mask_13 = _T_5114_13; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3090.4]
  assign io_sc2mac_dat_a_bits_mask_14 = _T_5114_14; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3091.4]
  assign io_sc2mac_dat_a_bits_mask_15 = _T_5114_15; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3092.4]
  assign io_sc2mac_dat_a_bits_mask_16 = _T_5114_16; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3093.4]
  assign io_sc2mac_dat_a_bits_mask_17 = _T_5114_17; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3094.4]
  assign io_sc2mac_dat_a_bits_mask_18 = _T_5114_18; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3095.4]
  assign io_sc2mac_dat_a_bits_mask_19 = _T_5114_19; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3096.4]
  assign io_sc2mac_dat_a_bits_mask_20 = _T_5114_20; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3097.4]
  assign io_sc2mac_dat_a_bits_mask_21 = _T_5114_21; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3098.4]
  assign io_sc2mac_dat_a_bits_mask_22 = _T_5114_22; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3099.4]
  assign io_sc2mac_dat_a_bits_mask_23 = _T_5114_23; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3100.4]
  assign io_sc2mac_dat_a_bits_mask_24 = _T_5114_24; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3101.4]
  assign io_sc2mac_dat_a_bits_mask_25 = _T_5114_25; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3102.4]
  assign io_sc2mac_dat_a_bits_mask_26 = _T_5114_26; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3103.4]
  assign io_sc2mac_dat_a_bits_mask_27 = _T_5114_27; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3104.4]
  assign io_sc2mac_dat_a_bits_mask_28 = _T_5114_28; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3105.4]
  assign io_sc2mac_dat_a_bits_mask_29 = _T_5114_29; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3106.4]
  assign io_sc2mac_dat_a_bits_mask_30 = _T_5114_30; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3107.4]
  assign io_sc2mac_dat_a_bits_mask_31 = _T_5114_31; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3108.4]
  assign io_sc2mac_dat_a_bits_mask_32 = _T_5114_32; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3109.4]
  assign io_sc2mac_dat_a_bits_mask_33 = _T_5114_33; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3110.4]
  assign io_sc2mac_dat_a_bits_mask_34 = _T_5114_34; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3111.4]
  assign io_sc2mac_dat_a_bits_mask_35 = _T_5114_35; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3112.4]
  assign io_sc2mac_dat_a_bits_mask_36 = _T_5114_36; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3113.4]
  assign io_sc2mac_dat_a_bits_mask_37 = _T_5114_37; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3114.4]
  assign io_sc2mac_dat_a_bits_mask_38 = _T_5114_38; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3115.4]
  assign io_sc2mac_dat_a_bits_mask_39 = _T_5114_39; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3116.4]
  assign io_sc2mac_dat_a_bits_mask_40 = _T_5114_40; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3117.4]
  assign io_sc2mac_dat_a_bits_mask_41 = _T_5114_41; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3118.4]
  assign io_sc2mac_dat_a_bits_mask_42 = _T_5114_42; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3119.4]
  assign io_sc2mac_dat_a_bits_mask_43 = _T_5114_43; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3120.4]
  assign io_sc2mac_dat_a_bits_mask_44 = _T_5114_44; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3121.4]
  assign io_sc2mac_dat_a_bits_mask_45 = _T_5114_45; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3122.4]
  assign io_sc2mac_dat_a_bits_mask_46 = _T_5114_46; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3123.4]
  assign io_sc2mac_dat_a_bits_mask_47 = _T_5114_47; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3124.4]
  assign io_sc2mac_dat_a_bits_mask_48 = _T_5114_48; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3125.4]
  assign io_sc2mac_dat_a_bits_mask_49 = _T_5114_49; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3126.4]
  assign io_sc2mac_dat_a_bits_mask_50 = _T_5114_50; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3127.4]
  assign io_sc2mac_dat_a_bits_mask_51 = _T_5114_51; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3128.4]
  assign io_sc2mac_dat_a_bits_mask_52 = _T_5114_52; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3129.4]
  assign io_sc2mac_dat_a_bits_mask_53 = _T_5114_53; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3130.4]
  assign io_sc2mac_dat_a_bits_mask_54 = _T_5114_54; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3131.4]
  assign io_sc2mac_dat_a_bits_mask_55 = _T_5114_55; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3132.4]
  assign io_sc2mac_dat_a_bits_mask_56 = _T_5114_56; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3133.4]
  assign io_sc2mac_dat_a_bits_mask_57 = _T_5114_57; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3134.4]
  assign io_sc2mac_dat_a_bits_mask_58 = _T_5114_58; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3135.4]
  assign io_sc2mac_dat_a_bits_mask_59 = _T_5114_59; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3136.4]
  assign io_sc2mac_dat_a_bits_mask_60 = _T_5114_60; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3137.4]
  assign io_sc2mac_dat_a_bits_mask_61 = _T_5114_61; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3138.4]
  assign io_sc2mac_dat_a_bits_mask_62 = _T_5114_62; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3139.4]
  assign io_sc2mac_dat_a_bits_mask_63 = _T_5114_63; // @[NV_NVDLA_CSC_dl.scala 1178:27:@3140.4]
  assign io_sc2mac_dat_a_bits_data_0 = _T_5776; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3342.4]
  assign io_sc2mac_dat_a_bits_data_1 = _T_5780; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3352.4]
  assign io_sc2mac_dat_a_bits_data_2 = _T_5784; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3362.4]
  assign io_sc2mac_dat_a_bits_data_3 = _T_5788; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3372.4]
  assign io_sc2mac_dat_a_bits_data_4 = _T_5792; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3382.4]
  assign io_sc2mac_dat_a_bits_data_5 = _T_5796; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3392.4]
  assign io_sc2mac_dat_a_bits_data_6 = _T_5800; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3402.4]
  assign io_sc2mac_dat_a_bits_data_7 = _T_5804; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3412.4]
  assign io_sc2mac_dat_a_bits_data_8 = _T_5808; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3422.4]
  assign io_sc2mac_dat_a_bits_data_9 = _T_5812; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3432.4]
  assign io_sc2mac_dat_a_bits_data_10 = _T_5816; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3442.4]
  assign io_sc2mac_dat_a_bits_data_11 = _T_5820; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3452.4]
  assign io_sc2mac_dat_a_bits_data_12 = _T_5824; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3462.4]
  assign io_sc2mac_dat_a_bits_data_13 = _T_5828; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3472.4]
  assign io_sc2mac_dat_a_bits_data_14 = _T_5832; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3482.4]
  assign io_sc2mac_dat_a_bits_data_15 = _T_5836; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3492.4]
  assign io_sc2mac_dat_a_bits_data_16 = _T_5840; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3502.4]
  assign io_sc2mac_dat_a_bits_data_17 = _T_5844; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3512.4]
  assign io_sc2mac_dat_a_bits_data_18 = _T_5848; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3522.4]
  assign io_sc2mac_dat_a_bits_data_19 = _T_5852; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3532.4]
  assign io_sc2mac_dat_a_bits_data_20 = _T_5856; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3542.4]
  assign io_sc2mac_dat_a_bits_data_21 = _T_5860; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3552.4]
  assign io_sc2mac_dat_a_bits_data_22 = _T_5864; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3562.4]
  assign io_sc2mac_dat_a_bits_data_23 = _T_5868; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3572.4]
  assign io_sc2mac_dat_a_bits_data_24 = _T_5872; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3582.4]
  assign io_sc2mac_dat_a_bits_data_25 = _T_5876; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3592.4]
  assign io_sc2mac_dat_a_bits_data_26 = _T_5880; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3602.4]
  assign io_sc2mac_dat_a_bits_data_27 = _T_5884; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3612.4]
  assign io_sc2mac_dat_a_bits_data_28 = _T_5888; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3622.4]
  assign io_sc2mac_dat_a_bits_data_29 = _T_5892; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3632.4]
  assign io_sc2mac_dat_a_bits_data_30 = _T_5896; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3642.4]
  assign io_sc2mac_dat_a_bits_data_31 = _T_5900; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3652.4]
  assign io_sc2mac_dat_a_bits_data_32 = _T_5904; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3662.4]
  assign io_sc2mac_dat_a_bits_data_33 = _T_5908; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3672.4]
  assign io_sc2mac_dat_a_bits_data_34 = _T_5912; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3682.4]
  assign io_sc2mac_dat_a_bits_data_35 = _T_5916; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3692.4]
  assign io_sc2mac_dat_a_bits_data_36 = _T_5920; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3702.4]
  assign io_sc2mac_dat_a_bits_data_37 = _T_5924; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3712.4]
  assign io_sc2mac_dat_a_bits_data_38 = _T_5928; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3722.4]
  assign io_sc2mac_dat_a_bits_data_39 = _T_5932; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3732.4]
  assign io_sc2mac_dat_a_bits_data_40 = _T_5936; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3742.4]
  assign io_sc2mac_dat_a_bits_data_41 = _T_5940; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3752.4]
  assign io_sc2mac_dat_a_bits_data_42 = _T_5944; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3762.4]
  assign io_sc2mac_dat_a_bits_data_43 = _T_5948; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3772.4]
  assign io_sc2mac_dat_a_bits_data_44 = _T_5952; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3782.4]
  assign io_sc2mac_dat_a_bits_data_45 = _T_5956; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3792.4]
  assign io_sc2mac_dat_a_bits_data_46 = _T_5960; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3802.4]
  assign io_sc2mac_dat_a_bits_data_47 = _T_5964; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3812.4]
  assign io_sc2mac_dat_a_bits_data_48 = _T_5968; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3822.4]
  assign io_sc2mac_dat_a_bits_data_49 = _T_5972; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3832.4]
  assign io_sc2mac_dat_a_bits_data_50 = _T_5976; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3842.4]
  assign io_sc2mac_dat_a_bits_data_51 = _T_5980; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3852.4]
  assign io_sc2mac_dat_a_bits_data_52 = _T_5984; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3862.4]
  assign io_sc2mac_dat_a_bits_data_53 = _T_5988; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3872.4]
  assign io_sc2mac_dat_a_bits_data_54 = _T_5992; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3882.4]
  assign io_sc2mac_dat_a_bits_data_55 = _T_5996; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3892.4]
  assign io_sc2mac_dat_a_bits_data_56 = _T_6000; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3902.4]
  assign io_sc2mac_dat_a_bits_data_57 = _T_6004; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3912.4]
  assign io_sc2mac_dat_a_bits_data_58 = _T_6008; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3922.4]
  assign io_sc2mac_dat_a_bits_data_59 = _T_6012; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3932.4]
  assign io_sc2mac_dat_a_bits_data_60 = _T_6016; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3942.4]
  assign io_sc2mac_dat_a_bits_data_61 = _T_6020; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3952.4]
  assign io_sc2mac_dat_a_bits_data_62 = _T_6024; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3962.4]
  assign io_sc2mac_dat_a_bits_data_63 = _T_6028; // @[NV_NVDLA_CSC_dl.scala 1181:34:@3972.4]
  assign io_sc2mac_dat_a_bits_pd = _T_4842; // @[NV_NVDLA_CSC_dl.scala 1176:25:@2937.4]
  assign io_sc2mac_dat_b_valid = _T_4838; // @[NV_NVDLA_CSC_dl.scala 1175:23:@2931.4]
  assign io_sc2mac_dat_b_bits_mask_0 = _T_5578_0; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3274.4]
  assign io_sc2mac_dat_b_bits_mask_1 = _T_5578_1; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3275.4]
  assign io_sc2mac_dat_b_bits_mask_2 = _T_5578_2; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3276.4]
  assign io_sc2mac_dat_b_bits_mask_3 = _T_5578_3; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3277.4]
  assign io_sc2mac_dat_b_bits_mask_4 = _T_5578_4; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3278.4]
  assign io_sc2mac_dat_b_bits_mask_5 = _T_5578_5; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3279.4]
  assign io_sc2mac_dat_b_bits_mask_6 = _T_5578_6; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3280.4]
  assign io_sc2mac_dat_b_bits_mask_7 = _T_5578_7; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3281.4]
  assign io_sc2mac_dat_b_bits_mask_8 = _T_5578_8; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3282.4]
  assign io_sc2mac_dat_b_bits_mask_9 = _T_5578_9; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3283.4]
  assign io_sc2mac_dat_b_bits_mask_10 = _T_5578_10; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3284.4]
  assign io_sc2mac_dat_b_bits_mask_11 = _T_5578_11; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3285.4]
  assign io_sc2mac_dat_b_bits_mask_12 = _T_5578_12; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3286.4]
  assign io_sc2mac_dat_b_bits_mask_13 = _T_5578_13; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3287.4]
  assign io_sc2mac_dat_b_bits_mask_14 = _T_5578_14; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3288.4]
  assign io_sc2mac_dat_b_bits_mask_15 = _T_5578_15; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3289.4]
  assign io_sc2mac_dat_b_bits_mask_16 = _T_5578_16; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3290.4]
  assign io_sc2mac_dat_b_bits_mask_17 = _T_5578_17; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3291.4]
  assign io_sc2mac_dat_b_bits_mask_18 = _T_5578_18; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3292.4]
  assign io_sc2mac_dat_b_bits_mask_19 = _T_5578_19; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3293.4]
  assign io_sc2mac_dat_b_bits_mask_20 = _T_5578_20; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3294.4]
  assign io_sc2mac_dat_b_bits_mask_21 = _T_5578_21; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3295.4]
  assign io_sc2mac_dat_b_bits_mask_22 = _T_5578_22; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3296.4]
  assign io_sc2mac_dat_b_bits_mask_23 = _T_5578_23; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3297.4]
  assign io_sc2mac_dat_b_bits_mask_24 = _T_5578_24; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3298.4]
  assign io_sc2mac_dat_b_bits_mask_25 = _T_5578_25; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3299.4]
  assign io_sc2mac_dat_b_bits_mask_26 = _T_5578_26; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3300.4]
  assign io_sc2mac_dat_b_bits_mask_27 = _T_5578_27; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3301.4]
  assign io_sc2mac_dat_b_bits_mask_28 = _T_5578_28; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3302.4]
  assign io_sc2mac_dat_b_bits_mask_29 = _T_5578_29; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3303.4]
  assign io_sc2mac_dat_b_bits_mask_30 = _T_5578_30; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3304.4]
  assign io_sc2mac_dat_b_bits_mask_31 = _T_5578_31; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3305.4]
  assign io_sc2mac_dat_b_bits_mask_32 = _T_5578_32; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3306.4]
  assign io_sc2mac_dat_b_bits_mask_33 = _T_5578_33; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3307.4]
  assign io_sc2mac_dat_b_bits_mask_34 = _T_5578_34; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3308.4]
  assign io_sc2mac_dat_b_bits_mask_35 = _T_5578_35; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3309.4]
  assign io_sc2mac_dat_b_bits_mask_36 = _T_5578_36; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3310.4]
  assign io_sc2mac_dat_b_bits_mask_37 = _T_5578_37; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3311.4]
  assign io_sc2mac_dat_b_bits_mask_38 = _T_5578_38; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3312.4]
  assign io_sc2mac_dat_b_bits_mask_39 = _T_5578_39; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3313.4]
  assign io_sc2mac_dat_b_bits_mask_40 = _T_5578_40; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3314.4]
  assign io_sc2mac_dat_b_bits_mask_41 = _T_5578_41; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3315.4]
  assign io_sc2mac_dat_b_bits_mask_42 = _T_5578_42; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3316.4]
  assign io_sc2mac_dat_b_bits_mask_43 = _T_5578_43; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3317.4]
  assign io_sc2mac_dat_b_bits_mask_44 = _T_5578_44; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3318.4]
  assign io_sc2mac_dat_b_bits_mask_45 = _T_5578_45; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3319.4]
  assign io_sc2mac_dat_b_bits_mask_46 = _T_5578_46; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3320.4]
  assign io_sc2mac_dat_b_bits_mask_47 = _T_5578_47; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3321.4]
  assign io_sc2mac_dat_b_bits_mask_48 = _T_5578_48; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3322.4]
  assign io_sc2mac_dat_b_bits_mask_49 = _T_5578_49; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3323.4]
  assign io_sc2mac_dat_b_bits_mask_50 = _T_5578_50; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3324.4]
  assign io_sc2mac_dat_b_bits_mask_51 = _T_5578_51; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3325.4]
  assign io_sc2mac_dat_b_bits_mask_52 = _T_5578_52; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3326.4]
  assign io_sc2mac_dat_b_bits_mask_53 = _T_5578_53; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3327.4]
  assign io_sc2mac_dat_b_bits_mask_54 = _T_5578_54; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3328.4]
  assign io_sc2mac_dat_b_bits_mask_55 = _T_5578_55; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3329.4]
  assign io_sc2mac_dat_b_bits_mask_56 = _T_5578_56; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3330.4]
  assign io_sc2mac_dat_b_bits_mask_57 = _T_5578_57; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3331.4]
  assign io_sc2mac_dat_b_bits_mask_58 = _T_5578_58; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3332.4]
  assign io_sc2mac_dat_b_bits_mask_59 = _T_5578_59; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3333.4]
  assign io_sc2mac_dat_b_bits_mask_60 = _T_5578_60; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3334.4]
  assign io_sc2mac_dat_b_bits_mask_61 = _T_5578_61; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3335.4]
  assign io_sc2mac_dat_b_bits_mask_62 = _T_5578_62; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3336.4]
  assign io_sc2mac_dat_b_bits_mask_63 = _T_5578_63; // @[NV_NVDLA_CSC_dl.scala 1179:27:@3337.4]
  assign io_sc2mac_dat_b_bits_data_0 = _T_5778; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3347.4]
  assign io_sc2mac_dat_b_bits_data_1 = _T_5782; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3357.4]
  assign io_sc2mac_dat_b_bits_data_2 = _T_5786; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3367.4]
  assign io_sc2mac_dat_b_bits_data_3 = _T_5790; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3377.4]
  assign io_sc2mac_dat_b_bits_data_4 = _T_5794; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3387.4]
  assign io_sc2mac_dat_b_bits_data_5 = _T_5798; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3397.4]
  assign io_sc2mac_dat_b_bits_data_6 = _T_5802; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3407.4]
  assign io_sc2mac_dat_b_bits_data_7 = _T_5806; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3417.4]
  assign io_sc2mac_dat_b_bits_data_8 = _T_5810; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3427.4]
  assign io_sc2mac_dat_b_bits_data_9 = _T_5814; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3437.4]
  assign io_sc2mac_dat_b_bits_data_10 = _T_5818; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3447.4]
  assign io_sc2mac_dat_b_bits_data_11 = _T_5822; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3457.4]
  assign io_sc2mac_dat_b_bits_data_12 = _T_5826; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3467.4]
  assign io_sc2mac_dat_b_bits_data_13 = _T_5830; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3477.4]
  assign io_sc2mac_dat_b_bits_data_14 = _T_5834; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3487.4]
  assign io_sc2mac_dat_b_bits_data_15 = _T_5838; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3497.4]
  assign io_sc2mac_dat_b_bits_data_16 = _T_5842; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3507.4]
  assign io_sc2mac_dat_b_bits_data_17 = _T_5846; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3517.4]
  assign io_sc2mac_dat_b_bits_data_18 = _T_5850; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3527.4]
  assign io_sc2mac_dat_b_bits_data_19 = _T_5854; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3537.4]
  assign io_sc2mac_dat_b_bits_data_20 = _T_5858; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3547.4]
  assign io_sc2mac_dat_b_bits_data_21 = _T_5862; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3557.4]
  assign io_sc2mac_dat_b_bits_data_22 = _T_5866; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3567.4]
  assign io_sc2mac_dat_b_bits_data_23 = _T_5870; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3577.4]
  assign io_sc2mac_dat_b_bits_data_24 = _T_5874; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3587.4]
  assign io_sc2mac_dat_b_bits_data_25 = _T_5878; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3597.4]
  assign io_sc2mac_dat_b_bits_data_26 = _T_5882; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3607.4]
  assign io_sc2mac_dat_b_bits_data_27 = _T_5886; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3617.4]
  assign io_sc2mac_dat_b_bits_data_28 = _T_5890; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3627.4]
  assign io_sc2mac_dat_b_bits_data_29 = _T_5894; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3637.4]
  assign io_sc2mac_dat_b_bits_data_30 = _T_5898; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3647.4]
  assign io_sc2mac_dat_b_bits_data_31 = _T_5902; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3657.4]
  assign io_sc2mac_dat_b_bits_data_32 = _T_5906; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3667.4]
  assign io_sc2mac_dat_b_bits_data_33 = _T_5910; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3677.4]
  assign io_sc2mac_dat_b_bits_data_34 = _T_5914; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3687.4]
  assign io_sc2mac_dat_b_bits_data_35 = _T_5918; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3697.4]
  assign io_sc2mac_dat_b_bits_data_36 = _T_5922; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3707.4]
  assign io_sc2mac_dat_b_bits_data_37 = _T_5926; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3717.4]
  assign io_sc2mac_dat_b_bits_data_38 = _T_5930; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3727.4]
  assign io_sc2mac_dat_b_bits_data_39 = _T_5934; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3737.4]
  assign io_sc2mac_dat_b_bits_data_40 = _T_5938; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3747.4]
  assign io_sc2mac_dat_b_bits_data_41 = _T_5942; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3757.4]
  assign io_sc2mac_dat_b_bits_data_42 = _T_5946; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3767.4]
  assign io_sc2mac_dat_b_bits_data_43 = _T_5950; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3777.4]
  assign io_sc2mac_dat_b_bits_data_44 = _T_5954; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3787.4]
  assign io_sc2mac_dat_b_bits_data_45 = _T_5958; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3797.4]
  assign io_sc2mac_dat_b_bits_data_46 = _T_5962; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3807.4]
  assign io_sc2mac_dat_b_bits_data_47 = _T_5966; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3817.4]
  assign io_sc2mac_dat_b_bits_data_48 = _T_5970; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3827.4]
  assign io_sc2mac_dat_b_bits_data_49 = _T_5974; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3837.4]
  assign io_sc2mac_dat_b_bits_data_50 = _T_5978; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3847.4]
  assign io_sc2mac_dat_b_bits_data_51 = _T_5982; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3857.4]
  assign io_sc2mac_dat_b_bits_data_52 = _T_5986; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3867.4]
  assign io_sc2mac_dat_b_bits_data_53 = _T_5990; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3877.4]
  assign io_sc2mac_dat_b_bits_data_54 = _T_5994; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3887.4]
  assign io_sc2mac_dat_b_bits_data_55 = _T_5998; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3897.4]
  assign io_sc2mac_dat_b_bits_data_56 = _T_6002; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3907.4]
  assign io_sc2mac_dat_b_bits_data_57 = _T_6006; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3917.4]
  assign io_sc2mac_dat_b_bits_data_58 = _T_6010; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3927.4]
  assign io_sc2mac_dat_b_bits_data_59 = _T_6014; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3937.4]
  assign io_sc2mac_dat_b_bits_data_60 = _T_6018; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3947.4]
  assign io_sc2mac_dat_b_bits_data_61 = _T_6022; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3957.4]
  assign io_sc2mac_dat_b_bits_data_62 = _T_6026; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3967.4]
  assign io_sc2mac_dat_b_bits_data_63 = _T_6030; // @[NV_NVDLA_CSC_dl.scala 1182:34:@3977.4]
  assign io_sc2mac_dat_b_bits_pd = _T_4846; // @[NV_NVDLA_CSC_dl.scala 1177:25:@2943.4]
  assign io_slcg_wg_en = 1'h0; // @[NV_NVDLA_CSC_dl.scala 249:15:@242.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_715 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_722 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_729 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_736 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_743 = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_750 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_757 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_771 = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_778 = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_785 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_792 = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_831 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_838 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_845 = _RAND_13[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_852 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_859 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_866 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_869 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_872 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_878 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_881 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_884 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_887 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_893 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_896 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_902 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_905 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_908 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_915 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_922 = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_932 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_939 = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_946 = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_953 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_960 = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_967 = _RAND_35[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_974 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_981 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_988 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_995 = _RAND_39[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1002 = _RAND_40[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1009 = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1016 = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1023 = _RAND_43[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1076 = _RAND_44[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_2217 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2211 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2208 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2231 = _RAND_48[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2225 = _RAND_49[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_2222 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1166 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1169 = _RAND_52[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1172 = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1177 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1180 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1183 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1186 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1189 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1211 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1214 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1217 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1220 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1225 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1228 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1231 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1234 = _RAND_66[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1279 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1290 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1306 = _RAND_69[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1335 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1329 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1332 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1361 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1366 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1369 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1390 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1404 = _RAND_77[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1407 = _RAND_78[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1410 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1413 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1416 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1419 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1424 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1427 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1539 = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1542 = _RAND_86[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1616 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1619 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1622 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1625 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1628 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1631 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1634 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1637 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1640 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1643 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1648 = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1651 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1654 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1657 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1660 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1663 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1666 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1759_0 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1759_1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1759_2 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1759_3 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1778 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1785 = _RAND_109[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1788 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1794 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1797 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1800 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1803 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1806 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1809 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1812 = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1815 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1818 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1821 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1943 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1946 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1949 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1952 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1955 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1958 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1963 = _RAND_127[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1966 = _RAND_128[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1969 = _RAND_129[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1972 = _RAND_130[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1975 = _RAND_131[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1978 = _RAND_132[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_2051 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_2063 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {16{`RANDOM}};
  _T_2074 = _RAND_135[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {16{`RANDOM}};
  _T_2082 = _RAND_136[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_2182 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_2185 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_2188 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_2191 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_2194 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_2197 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_2200 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_2203 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2214 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2228 = _RAND_146[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {8{`RANDOM}};
  _T_2611 = _RAND_147[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {4{`RANDOM}};
  _T_2613 = _RAND_148[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {4{`RANDOM}};
  _T_2615 = _RAND_149[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {4{`RANDOM}};
  _T_2617 = _RAND_150[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {4{`RANDOM}};
  _T_2619 = _RAND_151[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {4{`RANDOM}};
  _T_2621 = _RAND_152[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_3419 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_3689_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_3689_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_3689_2 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_3689_3 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_3689_4 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_3689_5 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_3689_6 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_3689_7 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_3689_8 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_3689_9 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_3689_10 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_3689_11 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_3689_12 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_3689_13 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_3689_14 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_3689_15 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_3689_16 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_3689_17 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_3689_18 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_3689_19 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_3689_20 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_3689_21 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_3689_22 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_3689_23 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_3689_24 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_3689_25 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_3689_26 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_3689_27 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_3689_28 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_3689_29 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_3689_30 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_3689_31 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_3689_32 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_3689_33 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_3689_34 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_3689_35 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_3689_36 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_3689_37 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_3689_38 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_3689_39 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_3689_40 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_3689_41 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_3689_42 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_3689_43 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_3689_44 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_3689_45 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_3689_46 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_3689_47 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_3689_48 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_3689_49 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_3689_50 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_3689_51 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_3689_52 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_3689_53 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_3689_54 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_3689_55 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_3689_56 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_3689_57 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_3689_58 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_3689_59 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_3689_60 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_3689_61 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_3689_62 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_3689_63 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_3889_0 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_3889_1 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_3889_2 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_3889_3 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_3889_4 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_3889_5 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_3889_6 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_3889_7 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_3889_8 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_3889_9 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3889_10 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3889_11 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3889_12 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3889_13 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3889_14 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3889_15 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3889_16 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3889_17 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3889_18 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3889_19 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3889_20 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3889_21 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3889_22 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3889_23 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3889_24 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3889_25 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3889_26 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3889_27 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3889_28 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3889_29 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3889_30 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3889_31 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3889_32 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3889_33 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3889_34 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3889_35 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3889_36 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3889_37 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3889_38 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3889_39 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3889_40 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3889_41 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3889_42 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3889_43 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3889_44 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3889_45 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3889_46 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3889_47 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3889_48 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3889_49 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3889_50 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3889_51 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3889_52 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3889_53 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3889_54 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3889_55 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3889_56 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3889_57 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3889_58 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3889_59 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3889_60 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3889_61 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3889_62 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3889_63 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_4022 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_4289_0 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_4289_1 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_4289_2 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_4289_3 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_4289_4 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_4289_5 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_4289_6 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_4289_7 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_4289_8 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_4289_9 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_4289_10 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_4289_11 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_4289_12 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_4289_13 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_4289_14 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_4289_15 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_4289_16 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_4289_17 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_4289_18 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_4289_19 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_4289_20 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_4289_21 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_4289_22 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_4289_23 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_4289_24 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_4289_25 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_4289_26 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_4289_27 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_4289_28 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_4289_29 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_4289_30 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_4289_31 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_4289_32 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_4289_33 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_4289_34 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_4289_35 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_4289_36 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_4289_37 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_4289_38 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_4289_39 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_4289_40 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_4289_41 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_4289_42 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_4289_43 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_4289_44 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_4289_45 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_4289_46 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_4289_47 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_4289_48 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_4289_49 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_4289_50 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_4289_51 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_4289_52 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_4289_53 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_4289_54 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_4289_55 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_4289_56 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_4289_57 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_4289_58 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_4289_59 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_4289_60 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_4289_61 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_4289_62 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_4289_63 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_4488 = _RAND_347[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_4492_0 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_4492_1 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_4492_2 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_4492_3 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_4492_4 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_4492_5 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_4492_6 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_4492_7 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_4492_8 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_4492_9 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_4492_10 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4492_11 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4492_12 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4492_13 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4492_14 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4492_15 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4492_16 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4492_17 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4492_18 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4492_19 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4492_20 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4492_21 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4492_22 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4492_23 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4492_24 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4492_25 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4492_26 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4492_27 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4492_28 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4492_29 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4492_30 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4492_31 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4492_32 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4492_33 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4492_34 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4492_35 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4492_36 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4492_37 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4492_38 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4492_39 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4492_40 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4492_41 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4492_42 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4492_43 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4492_44 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4492_45 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4492_46 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4492_47 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4492_48 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4492_49 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4492_50 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4492_51 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4492_52 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4492_53 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4492_54 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4492_55 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4492_56 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4492_57 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4492_58 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4492_59 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4492_60 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4492_61 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4492_62 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4492_63 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4829 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4835 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4838 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4842 = _RAND_415[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4846 = _RAND_416[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_5114_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_5114_1 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_5114_2 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_5114_3 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_5114_4 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_5114_5 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_5114_6 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_5114_7 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_5114_8 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_5114_9 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_5114_10 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_5114_11 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_5114_12 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_5114_13 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_5114_14 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_5114_15 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_5114_16 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_5114_17 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_5114_18 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_5114_19 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_5114_20 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_5114_21 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_5114_22 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_5114_23 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_5114_24 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_5114_25 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_5114_26 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_5114_27 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_5114_28 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_5114_29 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_5114_30 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_5114_31 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_5114_32 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_5114_33 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_5114_34 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_5114_35 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_5114_36 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_5114_37 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_5114_38 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_5114_39 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_5114_40 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_5114_41 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_5114_42 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_5114_43 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_5114_44 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_5114_45 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_5114_46 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_5114_47 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_5114_48 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_5114_49 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_5114_50 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_5114_51 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_5114_52 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_5114_53 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_5114_54 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_5114_55 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_5114_56 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_5114_57 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_5114_58 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_5114_59 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_5114_60 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_5114_61 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_5114_62 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_5114_63 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_5578_0 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_5578_1 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_5578_2 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_5578_3 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_5578_4 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_5578_5 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_5578_6 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_5578_7 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_5578_8 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_5578_9 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_5578_10 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_5578_11 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_5578_12 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_5578_13 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_5578_14 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_5578_15 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_5578_16 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_5578_17 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_5578_18 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_5578_19 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_5578_20 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_5578_21 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_5578_22 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_5578_23 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_5578_24 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_5578_25 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_5578_26 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_5578_27 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_5578_28 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_5578_29 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_5578_30 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_5578_31 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_5578_32 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_5578_33 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_5578_34 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_5578_35 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_5578_36 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_5578_37 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_5578_38 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_5578_39 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_5578_40 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_5578_41 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_5578_42 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_5578_43 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_5578_44 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_5578_45 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_5578_46 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_5578_47 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_5578_48 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_5578_49 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5578_50 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5578_51 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5578_52 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5578_53 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5578_54 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5578_55 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5578_56 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5578_57 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5578_58 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5578_59 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5578_60 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5578_61 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5578_62 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5578_63 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5776 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5778 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5780 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5782 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5784 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5786 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5788 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5790 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5792 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5794 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5796 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5798 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5800 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5802 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5804 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5806 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5808 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5810 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5812 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5814 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5816 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5818 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5820 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5822 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5824 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5826 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5828 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5830 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5832 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5834 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5836 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5838 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5840 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5842 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5844 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5846 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5848 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5850 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5852 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5854 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5856 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5858 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5860 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5862 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5864 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5866 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5868 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5870 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5872 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5874 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5876 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5878 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5880 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5882 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5884 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5886 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5888 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5890 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5892 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5894 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5896 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5898 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5900 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5902 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5904 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5906 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5908 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5910 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5912 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5914 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5916 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5918 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5920 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5922 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5924 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5926 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5928 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5930 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5932 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5934 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5936 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5938 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5940 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5942 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5944 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5946 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5948 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5950 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5952 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5954 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5956 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5958 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5960 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5962 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5964 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5966 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5968 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5970 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5972 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5974 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5976 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5978 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5980 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5982 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5984 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5986 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5988 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5990 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5992 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5994 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5996 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_5998 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_6000 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_6002 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_6004 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_6006 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_6008 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_6010 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_6012 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_6014 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_6016 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_6018 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_6020 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_6022 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_6024 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_6026 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_6028 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_6030 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (reset) begin
      _T_715 <= 1'h0;
    end else begin
      _T_715 <= _T_630;
    end
    if (reset) begin
      _T_722 <= 6'h0;
    end else begin
      if (_T_630) begin
        _T_722 <= 6'h1;
      end
    end
    if (reset) begin
      _T_729 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_729 <= {{2'd0}, _T_805};
      end
    end
    if (reset) begin
      _T_736 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_736 <= {{2'd0}, _T_798};
      end
    end
    if (reset) begin
      _T_743 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_743 <= _T_794;
      end
    end
    if (reset) begin
      _T_750 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_750 <= _T_797;
      end
    end
    if (reset) begin
      _T_757 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_757 <= io_reg2dp_dataout_width;
      end
    end
    if (reset) begin
      _T_771 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_771 <= _T_813;
      end
    end
    if (reset) begin
      _T_778 <= 12'h0;
    end else begin
      if (_T_715) begin
        _T_778 <= _T_800;
      end
    end
    if (reset) begin
      _T_785 <= 12'h0;
    end else begin
      if (_T_715) begin
        _T_785 <= _T_802;
      end
    end
    if (reset) begin
      _T_792 <= 14'h0;
    end else begin
      if (_T_630) begin
        if (io_reg2dp_skip_data_rls) begin
          _T_792 <= _T_807;
        end else begin
          _T_792 <= _T_809;
        end
      end
    end
    if (reset) begin
      _T_831 <= 34'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_831 <= 34'h3ffffffff;
        end else begin
          _T_831 <= 34'h0;
        end
      end
    end
    if (reset) begin
      _T_838 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_838 <= _T_1041;
      end
    end
    if (reset) begin
      _T_845 <= 14'h0;
    end else begin
      if (_T_630) begin
        _T_845 <= _T_1043;
      end
    end
    if (reset) begin
      _T_852 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_852 <= io_reg2dp_datain_width_ext;
      end
    end
    if (reset) begin
      _T_859 <= 13'h0;
    end else begin
      if (_T_630) begin
        _T_859 <= io_reg2dp_datain_height_ext;
      end
    end
    if (reset) begin
      _T_866 <= 11'h0;
    end else begin
      if (_T_630) begin
        _T_866 <= _T_1050;
      end
    end
    if (reset) begin
      _T_869 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_869 <= _T_643;
      end
    end
    if (reset) begin
      _T_872 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_872 <= _T_643;
      end
    end
    if (reset) begin
      _T_878 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_878 <= _T_643;
      end
    end
    if (reset) begin
      _T_881 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_881 <= _T_643;
      end
    end
    if (reset) begin
      _T_884 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_884 <= _T_643;
      end
    end
    if (reset) begin
      _T_887 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_887 <= _T_643;
      end
    end
    if (reset) begin
      _T_893 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_893 <= _T_643;
      end
    end
    if (reset) begin
      _T_896 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_896 <= _T_643;
      end
    end
    if (reset) begin
      _T_902 <= 3'h1;
    end else begin
      if (_T_630) begin
        _T_902 <= _T_643;
      end
    end
    if (reset) begin
      _T_905 <= 3'h1;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_905 <= _T_643;
        end else begin
          _T_905 <= 3'h1;
        end
      end
    end
    if (reset) begin
      _T_908 <= 3'h1;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_908 <= _T_643;
        end else begin
          _T_908 <= 3'h1;
        end
      end
    end
    if (reset) begin
      _T_915 <= 4'h0;
    end else begin
      if (_T_630) begin
        _T_915 <= _T_650;
      end
    end
    if (reset) begin
      _T_922 <= 4'h0;
    end else begin
      if (_T_630) begin
        _T_922 <= _T_704;
      end
    end
    if (reset) begin
      _T_932 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_932 <= 5'h0;
      end
    end
    if (reset) begin
      _T_939 <= 7'h0;
    end else begin
      if (_T_630) begin
        if (_T_686) begin
          _T_939 <= _T_679;
        end else begin
          _T_939 <= {{1'd0}, _T_685};
        end
      end
    end
    if (reset) begin
      _T_946 <= 7'h0;
    end else begin
      if (_T_630) begin
        _T_946 <= _T_690;
      end
    end
    if (reset) begin
      _T_953 <= 8'h0;
    end else begin
      if (_T_630) begin
        if (_T_686) begin
          _T_953 <= _T_693;
        end else begin
          _T_953 <= {{1'd0}, _T_698};
        end
      end
    end
    if (reset) begin
      _T_960 <= 7'h0;
    end else begin
      if (_T_630) begin
        _T_960 <= {{1'd0}, _T_662};
      end
    end
    if (reset) begin
      _T_967 <= 12'h0;
    end else begin
      if (_T_630) begin
        _T_967 <= _T_702;
      end
    end
    if (reset) begin
      _T_974 <= 6'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_974 <= 6'h1;
        end else begin
          _T_974 <= _T_707;
        end
      end
    end
    if (reset) begin
      _T_981 <= 6'h0;
    end else begin
      if (_T_630) begin
        if (_T_635) begin
          _T_981 <= 6'h1;
        end else begin
          _T_981 <= _T_711;
        end
      end
    end
    if (reset) begin
      _T_988 <= 16'h0;
    end else begin
      if (_T_630) begin
        _T_988 <= io_reg2dp_pad_value;
      end
    end
    if (reset) begin
      _T_995 <= 15'h0;
    end else begin
      if (_T_630) begin
        _T_995 <= _T_1054;
      end
    end
    if (reset) begin
      _T_1002 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_1002 <= _T_743;
      end
    end
    if (reset) begin
      _T_1009 <= 15'h0;
    end else begin
      if (_T_715) begin
        _T_1009 <= _T_743;
      end
    end
    if (reset) begin
      _T_1016 <= 14'h0;
    end else begin
      if (_T_626) begin
        _T_1016 <= _T_792;
      end
    end
    if (reset) begin
      _T_1023 <= 15'h0;
    end else begin
      if (_T_626) begin
        _T_1023 <= _T_813;
      end
    end
    if (reset) begin
      _T_2217 <= 1'h0;
    end else begin
      _T_2217 <= _T_2214;
    end
    if (reset) begin
      _T_2211 <= 1'h0;
    end else begin
      _T_2211 <= _T_2208;
    end
    if (reset) begin
      _T_2208 <= 1'h0;
    end else begin
      _T_2208 <= _T_1958;
    end
    if (reset) begin
      _T_2231 <= 27'h0;
    end else begin
      if (_T_2214) begin
        _T_2231 <= _T_2228;
      end
    end
    if (reset) begin
      _T_2225 <= 27'h0;
    end else begin
      if (_T_2208) begin
        _T_2225 <= _T_2222;
      end
    end
    if (reset) begin
      _T_2222 <= 27'h0;
    end else begin
      if (_T_1958) begin
        _T_2222 <= _T_2240;
      end
    end
    if (reset) begin
      _T_1166 <= 1'h0;
    end else begin
      _T_1166 <= _T_1161;
    end
    if (reset) begin
      _T_1169 <= 14'h0;
    end else begin
      if (_T_1161) begin
        if (_T_1154) begin
          _T_1169 <= _T_729;
        end else begin
          _T_1169 <= _T_1016;
        end
      end
    end
    if (reset) begin
      _T_1172 <= 15'h0;
    end else begin
      if (_T_1161) begin
        if (_T_1154) begin
          _T_1172 <= _T_771;
        end else begin
          _T_1172 <= _T_1023;
        end
      end
    end
    if (reset) begin
      _T_1177 <= 1'h0;
    end else begin
      _T_1177 <= io_sg2dl_pd_valid;
    end
    if (reset) begin
      _T_1180 <= 1'h0;
    end else begin
      _T_1180 <= _T_1177;
    end
    if (reset) begin
      _T_1183 <= 1'h0;
    end else begin
      _T_1183 <= _T_1180;
    end
    if (reset) begin
      _T_1186 <= 1'h0;
    end else begin
      _T_1186 <= _T_1183;
    end
    if (reset) begin
      _T_1189 <= 1'h0;
    end else begin
      _T_1189 <= _T_1186;
    end
    if (reset) begin
      _T_1211 <= 1'h0;
    end else begin
      _T_1211 <= _T_1189;
    end
    if (reset) begin
      _T_1214 <= 1'h0;
    end else begin
      _T_1214 <= _T_1211;
    end
    if (reset) begin
      _T_1217 <= 1'h0;
    end else begin
      _T_1217 <= _T_1214;
    end
    if (reset) begin
      _T_1220 <= 1'h0;
    end else begin
      _T_1220 <= _T_1217;
    end
    if (reset) begin
      _T_1225 <= 31'h0;
    end else begin
      if (_T_1189) begin
        _T_1225 <= _T_1222;
      end
    end
    if (reset) begin
      _T_1228 <= 31'h0;
    end else begin
      if (_T_1211) begin
        _T_1228 <= _T_1225;
      end
    end
    if (reset) begin
      _T_1231 <= 31'h0;
    end else begin
      if (_T_1214) begin
        _T_1231 <= _T_1228;
      end
    end
    if (reset) begin
      _T_1234 <= 31'h0;
    end else begin
      if (_T_1217) begin
        _T_1234 <= _T_1231;
      end
    end
    if (reset) begin
      _T_1279 <= 5'h0;
    end else begin
      if (_T_630) begin
        _T_1279 <= 5'h0;
      end else begin
        if (_T_1287) begin
          _T_1279 <= 5'h0;
        end else begin
          _T_1279 <= _T_1284;
        end
      end
    end
    if (reset) begin
      _T_1290 <= 2'h0;
    end else begin
      if (_T_1300) begin
        if (_T_1301) begin
          _T_1290 <= 2'h0;
        end else begin
          _T_1290 <= _T_1295;
        end
      end
    end
    if (reset) begin
      _T_1306 <= 7'h0;
    end else begin
      if (_T_1318) begin
        if (_T_630) begin
          _T_1306 <= 7'h0;
        end else begin
          if (_T_1321) begin
            _T_1306 <= 7'h0;
          end else begin
            if (_T_1316) begin
              _T_1306 <= 7'h0;
            end else begin
              _T_1306 <= _T_1313;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1335 <= 1'h0;
    end else begin
      if (_T_1242) begin
        _T_1335 <= 1'h1;
      end else begin
        if (_T_1355) begin
          _T_1335 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_1329 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1329 <= 1'h0;
      end else begin
        if (_T_1242) begin
          _T_1329 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_1332 <= 1'h0;
    end else begin
      _T_1332 <= _T_1343;
    end
    if (reset) begin
      _T_1361 <= 8'h0;
    end else begin
      if (_T_1358) begin
        _T_1361 <= _T_1363;
      end
    end
    if (reset) begin
      _T_1366 <= 13'h0;
    end else begin
      if (_T_1384) begin
        if (_T_630) begin
          _T_1366 <= {{9'd0}, _T_648};
        end else begin
          if (_T_1378) begin
            _T_1366 <= _T_1369;
          end else begin
            if (_T_1374) begin
              _T_1366 <= {{9'd0}, _T_648};
            end else begin
              _T_1366 <= _T_1371;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1369 <= 13'h0;
    end else begin
      if (_T_1387) begin
        if (_T_630) begin
          _T_1369 <= {{9'd0}, _T_648};
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              _T_1369 <= {{9'd0}, _T_648};
            end else begin
              _T_1369 <= _T_1371;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1390 <= 11'h0;
    end else begin
      if (_T_1394) begin
        if (_T_630) begin
          _T_1390 <= 11'h0;
        end else begin
          if (_T_1269) begin
            _T_1390 <= 11'h0;
          end else begin
            _T_1390 <= _T_1399;
          end
        end
      end
    end
    if (reset) begin
      _T_1404 <= 14'h0;
    end else begin
      if (_T_1448) begin
        if (_T_630) begin
          if (_T_635) begin
            _T_1404 <= 14'h0;
          end else begin
            _T_1404 <= _T_1431;
          end
        end else begin
          if (_T_1378) begin
            _T_1404 <= _T_1407;
          end else begin
            if (_T_1374) begin
              if (_T_635) begin
                _T_1404 <= 14'h0;
              end else begin
                _T_1404 <= _T_1431;
              end
            end else begin
              _T_1404 <= _T_1434;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1407 <= 14'h0;
    end else begin
      if (_T_1454) begin
        if (_T_630) begin
          if (_T_635) begin
            _T_1407 <= 14'h0;
          end else begin
            _T_1407 <= _T_1431;
          end
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              if (_T_635) begin
                _T_1407 <= 14'h0;
              end else begin
                _T_1407 <= _T_1431;
              end
            end else begin
              _T_1407 <= _T_1434;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1410 <= 16'h0;
    end else begin
      if (_T_1448) begin
        if (_T_715) begin
          _T_1410 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1410 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1410 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1410 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1410 <= _T_1493;
                end else begin
                  if (_T_1495) begin
                    _T_1410 <= _T_1413;
                  end else begin
                    _T_1410 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1413 <= 16'h0;
    end else begin
      if (_T_1454) begin
        if (_T_715) begin
          _T_1413 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1413 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1413 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1413 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1413 <= _T_1493;
                end else begin
                  if (!(_T_1495)) begin
                    _T_1413 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1416 <= 16'h0;
    end else begin
      if (_T_1526) begin
        if (_T_715) begin
          _T_1416 <= {{9'd0}, _T_939};
        end else begin
          if (_T_1477) begin
            _T_1416 <= {{9'd0}, _T_939};
          end else begin
            if (_T_1481) begin
              _T_1416 <= _T_1483;
            end else begin
              if (_T_1485) begin
                _T_1416 <= _T_1487;
              end else begin
                if (_T_1490) begin
                  _T_1416 <= _T_1493;
                end else begin
                  if (_T_1495) begin
                    _T_1416 <= _T_1413;
                  end else begin
                    _T_1416 <= _T_1497;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1419 <= 13'h2;
    end else begin
      if (_T_1466) begin
        _T_1419 <= 13'h2;
      end else begin
        if (_T_1468) begin
          _T_1419 <= _T_1471;
        end
      end
    end
    if (reset) begin
      _T_1424 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1424 <= _T_1536;
      end
    end
    if (reset) begin
      _T_1427 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1528) begin
          _T_1427 <= 1'h1;
        end else begin
          if (_T_1424) begin
            _T_1427 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_1539 <= 14'h0;
    end else begin
      if (_T_1560) begin
        if (_T_1550) begin
          _T_1539 <= _T_1546;
        end else begin
          if (_T_1378) begin
            _T_1539 <= _T_1542;
          end else begin
            if (_T_1374) begin
              _T_1539 <= _T_1548;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1542 <= 14'h0;
    end else begin
      if (_T_1387) begin
        if (_T_1550) begin
          _T_1542 <= _T_1546;
        end else begin
          if (!(_T_1378)) begin
            if (_T_1374) begin
              _T_1542 <= _T_1548;
            end else begin
              _T_1542 <= _T_1539;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_1616 <= 1'h0;
    end else begin
      _T_1616 <= _T_1600;
    end
    if (reset) begin
      _T_1619 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1619 <= _T_1605;
      end
    end
    if (reset) begin
      _T_1622 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1622 <= _T_1290;
      end
    end
    if (reset) begin
      _T_1625 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1602) begin
          _T_1625 <= _T_1603;
        end else begin
          _T_1625 <= _T_1268;
        end
      end
    end
    if (reset) begin
      _T_1628 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1628 <= _T_1391;
      end
    end
    if (reset) begin
      _T_1631 <= 1'h0;
    end else begin
      if (_T_1358) begin
        if (_T_1242) begin
          _T_1631 <= 1'h1;
        end else begin
          if (_T_1355) begin
            _T_1631 <= 1'h0;
          end else begin
            _T_1631 <= _T_1335;
          end
        end
      end
    end
    if (reset) begin
      _T_1634 <= 2'h0;
    end else begin
      if (_T_1358) begin
        _T_1634 <= _T_1267;
      end
    end
    if (reset) begin
      _T_1637 <= 1'h0;
    end else begin
      if (_T_1608) begin
        _T_1637 <= _T_1242;
      end
    end
    if (reset) begin
      _T_1640 <= 9'h0;
    end else begin
      if (_T_1358) begin
        _T_1640 <= _T_1613;
      end
    end
    if (reset) begin
      _T_1643 <= 1'h0;
    end else begin
      if (_T_1358) begin
        _T_1643 <= _T_1645;
      end
    end
    if (reset) begin
      _T_1648 <= 13'h0;
    end else begin
      if (_T_1394) begin
        if (_T_630) begin
          _T_1648 <= 13'h0;
        end else begin
          if (_T_1673) begin
            _T_1648 <= 13'h0;
          end else begin
            _T_1648 <= _T_1676;
          end
        end
      end
    end
    if (reset) begin
      _T_1651 <= 13'h0;
    end else begin
      if (_T_1682) begin
        _T_1651 <= _T_1648;
      end
    end
    if (reset) begin
      _T_1654 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1654 <= _T_1684;
      end
    end
    if (reset) begin
      _T_1657 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1657 <= _T_1686;
      end
    end
    if (reset) begin
      _T_1660 <= 13'h0;
    end else begin
      if (_T_1715) begin
        _T_1660 <= _T_1688;
      end
    end
    if (reset) begin
      _T_1663 <= 13'h0;
    end else begin
      if (_T_1716) begin
        _T_1663 <= _T_1692;
      end
    end
    if (reset) begin
      _T_1666 <= 13'h0;
    end else begin
      _T_1666 <= _GEN_95[12:0];
    end
    if (reset) begin
      _T_1759_0 <= 13'h1fff;
    end else begin
      _T_1759_0 <= _GEN_96[12:0];
    end
    if (reset) begin
      _T_1759_1 <= 13'h1fff;
    end else begin
      _T_1759_1 <= _GEN_97[12:0];
    end
    if (reset) begin
      _T_1759_2 <= 13'h1fff;
    end else begin
      _T_1759_2 <= _GEN_98[12:0];
    end
    if (reset) begin
      _T_1759_3 <= 13'h1fff;
    end else begin
      _T_1759_3 <= _GEN_99[12:0];
    end
    if (reset) begin
      _T_1778 <= 1'h0;
    end else begin
      _T_1778 <= _T_1891;
    end
    if (reset) begin
      _T_1785 <= 15'h1fff;
    end else begin
      if (_T_1922) begin
        if (_T_1850) begin
          _T_1785 <= 15'h1fff;
        end else begin
          if (_T_1840) begin
            _T_1785 <= _T_1849;
          end else begin
            _T_1785 <= _T_1833;
          end
        end
      end
    end
    if (reset) begin
      _T_1788 <= 1'h0;
    end else begin
      _T_1788 <= _T_1332;
    end
    if (reset) begin
      _T_1794 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1794 <= _T_1619;
      end
    end
    if (reset) begin
      _T_1797 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1797 <= _T_1622;
      end
    end
    if (reset) begin
      _T_1800 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1800 <= _T_1625;
      end
    end
    if (reset) begin
      _T_1803 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1803 <= _T_1628;
      end
    end
    if (reset) begin
      _T_1806 <= 8'h0;
    end else begin
      if (_T_1335) begin
        _T_1806 <= _T_1361;
      end
    end
    if (reset) begin
      _T_1809 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1809 <= _T_1631;
      end
    end
    if (reset) begin
      _T_1812 <= 2'h0;
    end else begin
      if (_T_1335) begin
        _T_1812 <= _T_1634;
      end
    end
    if (reset) begin
      _T_1815 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1815 <= _T_1637;
      end
    end
    if (reset) begin
      _T_1818 <= 1'h0;
    end else begin
      if (_T_1335) begin
        _T_1818 <= _T_1643;
      end
    end
    if (reset) begin
      _T_1821 <= 9'h0;
    end else begin
      if (_T_1335) begin
        _T_1821 <= _T_1640;
      end else begin
        _T_1821 <= {{8'd0}, _T_1335};
      end
    end
    if (reset) begin
      _T_1943 <= 1'h0;
    end else begin
      _T_1943 <= _T_1788;
    end
    if (reset) begin
      _T_1946 <= 1'h0;
    end else begin
      _T_1946 <= _T_1943;
    end
    if (reset) begin
      _T_1949 <= 1'h0;
    end else begin
      _T_1949 <= _T_1946;
    end
    if (reset) begin
      _T_1952 <= 1'h0;
    end else begin
      _T_1952 <= _T_1949;
    end
    if (reset) begin
      _T_1955 <= 1'h0;
    end else begin
      _T_1955 <= _T_1952;
    end
    if (reset) begin
      _T_1958 <= 1'h0;
    end else begin
      _T_1958 <= _T_1955;
    end
    if (reset) begin
      _T_1963 <= 29'h0;
    end else begin
      if (_T_1788) begin
        _T_1963 <= _T_1938;
      end
    end
    if (reset) begin
      _T_1966 <= 29'h0;
    end else begin
      if (_T_1943) begin
        _T_1966 <= _T_1963;
      end
    end
    if (reset) begin
      _T_1969 <= 29'h0;
    end else begin
      if (_T_1946) begin
        _T_1969 <= _T_1966;
      end
    end
    if (reset) begin
      _T_1972 <= 29'h0;
    end else begin
      if (_T_1949) begin
        _T_1972 <= _T_1969;
      end
    end
    if (reset) begin
      _T_1975 <= 29'h0;
    end else begin
      if (_T_1952) begin
        _T_1975 <= _T_1972;
      end
    end
    if (reset) begin
      _T_1978 <= 29'h0;
    end else begin
      if (_T_1955) begin
        _T_1978 <= _T_1975;
      end
    end
    if (reset) begin
      _T_2051 <= 1'h1;
    end else begin
      if (io_sc2buf_dat_rd_data_valid) begin
        _T_2051 <= 1'h0;
      end
    end
    if (reset) begin
      _T_2063 <= 1'h1;
    end else begin
      if (_T_2108) begin
        _T_2063 <= 1'h0;
      end else begin
        if (io_sc2buf_dat_rd_data_valid) begin
          _T_2063 <= _T_2051;
        end
      end
    end
    if (io_sc2buf_dat_rd_data_valid) begin
      _T_2074 <= io_sc2buf_dat_rd_data_bits;
    end
    if (_T_2108) begin
      _T_2082 <= _T_2074;
    end
    if (reset) begin
      _T_2182 <= 8'h0;
    end else begin
      if (_T_2388) begin
        if (_T_630) begin
          _T_2182 <= 8'h40;
        end else begin
          if (_T_2344) begin
            _T_2182 <= _T_2194;
          end else begin
            if (_T_2345) begin
              _T_2182 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2182 <= 8'h40;
              end else begin
                _T_2182 <= _T_2313;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2185 <= 8'h0;
    end else begin
      if (_T_2394) begin
        if (_T_630) begin
          _T_2185 <= 8'h40;
        end else begin
          if (_T_2355) begin
            _T_2185 <= _T_2197;
          end else begin
            if (_T_2356) begin
              _T_2185 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2185 <= 8'h40;
              end else begin
                _T_2185 <= _T_2322;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2188 <= 8'h0;
    end else begin
      if (_T_2400) begin
        if (_T_630) begin
          _T_2188 <= 8'h40;
        end else begin
          if (_T_2366) begin
            _T_2188 <= _T_2200;
          end else begin
            if (_T_2367) begin
              _T_2188 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2188 <= 8'h40;
              end else begin
                _T_2188 <= _T_2331;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2191 <= 8'h0;
    end else begin
      if (_T_2406) begin
        if (_T_630) begin
          _T_2191 <= 8'h40;
        end else begin
          if (_T_2377) begin
            _T_2191 <= _T_2203;
          end else begin
            if (_T_2378) begin
              _T_2191 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2191 <= 8'h40;
              end else begin
                _T_2191 <= _T_2340;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2194 <= 8'h0;
    end else begin
      if (_T_2411) begin
        if (_T_630) begin
          _T_2194 <= 8'h40;
        end else begin
          if (!(_T_2344)) begin
            if (_T_2345) begin
              _T_2194 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2194 <= 8'h40;
              end else begin
                _T_2194 <= _T_2313;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2197 <= 8'h0;
    end else begin
      if (_T_2419) begin
        if (_T_630) begin
          _T_2197 <= 8'h40;
        end else begin
          if (!(_T_2355)) begin
            if (_T_2356) begin
              _T_2197 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2197 <= 8'h40;
              end else begin
                _T_2197 <= _T_2322;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2200 <= 8'h0;
    end else begin
      if (_T_2427) begin
        if (_T_630) begin
          _T_2200 <= 8'h40;
        end else begin
          if (!(_T_2366)) begin
            if (_T_2367) begin
              _T_2200 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2200 <= 8'h40;
              end else begin
                _T_2200 <= _T_2331;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2203 <= 8'h0;
    end else begin
      if (_T_2435) begin
        if (_T_630) begin
          _T_2203 <= 8'h40;
        end else begin
          if (!(_T_2377)) begin
            if (_T_2378) begin
              _T_2203 <= 8'h40;
            end else begin
              if (_T_2307) begin
                _T_2203 <= 8'h40;
              end else begin
                _T_2203 <= _T_2340;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_2214 <= 1'h0;
    end else begin
      _T_2214 <= _T_2211;
    end
    if (reset) begin
      _T_2228 <= 27'h0;
    end else begin
      if (_T_2211) begin
        _T_2228 <= _T_2225;
      end
    end
    _T_2611 <= _GEN_149[255:0];
    _T_2613 <= _GEN_150[127:0];
    if (_T_2821) begin
      _T_2615 <= _T_2613;
    end
    _T_2617 <= _GEN_151[127:0];
    if (_T_2821) begin
      _T_2619 <= _T_2617;
    end
    _T_2621 <= _GEN_154[127:0];
    if (reset) begin
      _T_3419 <= 1'h0;
    end else begin
      _T_3419 <= _T_2248;
    end
    if (reset) begin
      _T_3689_0 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_0 <= _T_3220;
      end
    end
    if (reset) begin
      _T_3689_1 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_1 <= _T_3222;
      end
    end
    if (reset) begin
      _T_3689_2 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_2 <= _T_3224;
      end
    end
    if (reset) begin
      _T_3689_3 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_3 <= _T_3226;
      end
    end
    if (reset) begin
      _T_3689_4 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_4 <= _T_3228;
      end
    end
    if (reset) begin
      _T_3689_5 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_5 <= _T_3230;
      end
    end
    if (reset) begin
      _T_3689_6 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_6 <= _T_3232;
      end
    end
    if (reset) begin
      _T_3689_7 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_7 <= _T_3234;
      end
    end
    if (reset) begin
      _T_3689_8 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_8 <= _T_3236;
      end
    end
    if (reset) begin
      _T_3689_9 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_9 <= _T_3238;
      end
    end
    if (reset) begin
      _T_3689_10 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_10 <= _T_3240;
      end
    end
    if (reset) begin
      _T_3689_11 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_11 <= _T_3242;
      end
    end
    if (reset) begin
      _T_3689_12 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_12 <= _T_3244;
      end
    end
    if (reset) begin
      _T_3689_13 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_13 <= _T_3246;
      end
    end
    if (reset) begin
      _T_3689_14 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_14 <= _T_3248;
      end
    end
    if (reset) begin
      _T_3689_15 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_15 <= _T_3250;
      end
    end
    if (reset) begin
      _T_3689_16 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_16 <= _T_3252;
      end
    end
    if (reset) begin
      _T_3689_17 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_17 <= _T_3254;
      end
    end
    if (reset) begin
      _T_3689_18 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_18 <= _T_3256;
      end
    end
    if (reset) begin
      _T_3689_19 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_19 <= _T_3258;
      end
    end
    if (reset) begin
      _T_3689_20 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_20 <= _T_3260;
      end
    end
    if (reset) begin
      _T_3689_21 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_21 <= _T_3262;
      end
    end
    if (reset) begin
      _T_3689_22 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_22 <= _T_3264;
      end
    end
    if (reset) begin
      _T_3689_23 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_23 <= _T_3266;
      end
    end
    if (reset) begin
      _T_3689_24 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_24 <= _T_3268;
      end
    end
    if (reset) begin
      _T_3689_25 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_25 <= _T_3270;
      end
    end
    if (reset) begin
      _T_3689_26 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_26 <= _T_3272;
      end
    end
    if (reset) begin
      _T_3689_27 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_27 <= _T_3274;
      end
    end
    if (reset) begin
      _T_3689_28 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_28 <= _T_3276;
      end
    end
    if (reset) begin
      _T_3689_29 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_29 <= _T_3278;
      end
    end
    if (reset) begin
      _T_3689_30 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_30 <= _T_3280;
      end
    end
    if (reset) begin
      _T_3689_31 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_31 <= _T_3282;
      end
    end
    if (reset) begin
      _T_3689_32 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_32 <= _T_3284;
      end
    end
    if (reset) begin
      _T_3689_33 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_33 <= _T_3286;
      end
    end
    if (reset) begin
      _T_3689_34 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_34 <= _T_3288;
      end
    end
    if (reset) begin
      _T_3689_35 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_35 <= _T_3290;
      end
    end
    if (reset) begin
      _T_3689_36 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_36 <= _T_3292;
      end
    end
    if (reset) begin
      _T_3689_37 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_37 <= _T_3294;
      end
    end
    if (reset) begin
      _T_3689_38 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_38 <= _T_3296;
      end
    end
    if (reset) begin
      _T_3689_39 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_39 <= _T_3298;
      end
    end
    if (reset) begin
      _T_3689_40 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_40 <= _T_3300;
      end
    end
    if (reset) begin
      _T_3689_41 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_41 <= _T_3302;
      end
    end
    if (reset) begin
      _T_3689_42 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_42 <= _T_3304;
      end
    end
    if (reset) begin
      _T_3689_43 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_43 <= _T_3306;
      end
    end
    if (reset) begin
      _T_3689_44 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_44 <= _T_3308;
      end
    end
    if (reset) begin
      _T_3689_45 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_45 <= _T_3310;
      end
    end
    if (reset) begin
      _T_3689_46 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_46 <= _T_3312;
      end
    end
    if (reset) begin
      _T_3689_47 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_47 <= _T_3314;
      end
    end
    if (reset) begin
      _T_3689_48 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_48 <= _T_3316;
      end
    end
    if (reset) begin
      _T_3689_49 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_49 <= _T_3318;
      end
    end
    if (reset) begin
      _T_3689_50 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_50 <= _T_3320;
      end
    end
    if (reset) begin
      _T_3689_51 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_51 <= _T_3322;
      end
    end
    if (reset) begin
      _T_3689_52 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_52 <= _T_3324;
      end
    end
    if (reset) begin
      _T_3689_53 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_53 <= _T_3326;
      end
    end
    if (reset) begin
      _T_3689_54 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_54 <= _T_3328;
      end
    end
    if (reset) begin
      _T_3689_55 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_55 <= _T_3330;
      end
    end
    if (reset) begin
      _T_3689_56 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_56 <= _T_3332;
      end
    end
    if (reset) begin
      _T_3689_57 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_57 <= _T_3334;
      end
    end
    if (reset) begin
      _T_3689_58 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_58 <= _T_3336;
      end
    end
    if (reset) begin
      _T_3689_59 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_59 <= _T_3338;
      end
    end
    if (reset) begin
      _T_3689_60 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_60 <= _T_3340;
      end
    end
    if (reset) begin
      _T_3689_61 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_61 <= _T_3342;
      end
    end
    if (reset) begin
      _T_3689_62 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_62 <= _T_3344;
      end
    end
    if (reset) begin
      _T_3689_63 <= 1'h0;
    end else begin
      if (_T_2248) begin
        _T_3689_63 <= _T_3346;
      end
    end
    if (_T_3956) begin
      if (_T_2888) begin
        _T_3889_0 <= _T_2749;
      end else begin
        _T_3889_0 <= _T_2546;
      end
    end
    if (_T_3957) begin
      if (_T_2888) begin
        _T_3889_1 <= _T_2750;
      end else begin
        _T_3889_1 <= _T_2547;
      end
    end
    if (_T_3958) begin
      if (_T_2888) begin
        _T_3889_2 <= _T_2751;
      end else begin
        _T_3889_2 <= _T_2548;
      end
    end
    if (_T_3959) begin
      if (_T_2888) begin
        _T_3889_3 <= _T_2752;
      end else begin
        _T_3889_3 <= _T_2549;
      end
    end
    if (_T_3960) begin
      if (_T_2888) begin
        _T_3889_4 <= _T_2753;
      end else begin
        _T_3889_4 <= _T_2550;
      end
    end
    if (_T_3961) begin
      if (_T_2888) begin
        _T_3889_5 <= _T_2754;
      end else begin
        _T_3889_5 <= _T_2551;
      end
    end
    if (_T_3962) begin
      if (_T_2888) begin
        _T_3889_6 <= _T_2755;
      end else begin
        _T_3889_6 <= _T_2552;
      end
    end
    if (_T_3963) begin
      if (_T_2888) begin
        _T_3889_7 <= _T_2756;
      end else begin
        _T_3889_7 <= _T_2553;
      end
    end
    if (_T_3964) begin
      if (_T_2888) begin
        _T_3889_8 <= _T_2757;
      end else begin
        _T_3889_8 <= _T_2554;
      end
    end
    if (_T_3965) begin
      if (_T_2888) begin
        _T_3889_9 <= _T_2758;
      end else begin
        _T_3889_9 <= _T_2555;
      end
    end
    if (_T_3966) begin
      if (_T_2888) begin
        _T_3889_10 <= _T_2759;
      end else begin
        _T_3889_10 <= _T_2556;
      end
    end
    if (_T_3967) begin
      if (_T_2888) begin
        _T_3889_11 <= _T_2760;
      end else begin
        _T_3889_11 <= _T_2557;
      end
    end
    if (_T_3968) begin
      if (_T_2888) begin
        _T_3889_12 <= _T_2761;
      end else begin
        _T_3889_12 <= _T_2558;
      end
    end
    if (_T_3969) begin
      if (_T_2888) begin
        _T_3889_13 <= _T_2762;
      end else begin
        _T_3889_13 <= _T_2559;
      end
    end
    if (_T_3970) begin
      if (_T_2888) begin
        _T_3889_14 <= _T_2763;
      end else begin
        _T_3889_14 <= _T_2560;
      end
    end
    if (_T_3971) begin
      if (_T_2888) begin
        _T_3889_15 <= _T_2764;
      end else begin
        _T_3889_15 <= _T_2561;
      end
    end
    if (_T_3972) begin
      if (_T_2888) begin
        _T_3889_16 <= _T_2765;
      end else begin
        _T_3889_16 <= _T_2562;
      end
    end
    if (_T_3973) begin
      if (_T_2888) begin
        _T_3889_17 <= _T_2766;
      end else begin
        _T_3889_17 <= _T_2563;
      end
    end
    if (_T_3974) begin
      if (_T_2888) begin
        _T_3889_18 <= _T_2767;
      end else begin
        _T_3889_18 <= _T_2564;
      end
    end
    if (_T_3975) begin
      if (_T_2888) begin
        _T_3889_19 <= _T_2768;
      end else begin
        _T_3889_19 <= _T_2565;
      end
    end
    if (_T_3976) begin
      if (_T_2888) begin
        _T_3889_20 <= _T_2769;
      end else begin
        _T_3889_20 <= _T_2566;
      end
    end
    if (_T_3977) begin
      if (_T_2888) begin
        _T_3889_21 <= _T_2770;
      end else begin
        _T_3889_21 <= _T_2567;
      end
    end
    if (_T_3978) begin
      if (_T_2888) begin
        _T_3889_22 <= _T_2771;
      end else begin
        _T_3889_22 <= _T_2568;
      end
    end
    if (_T_3979) begin
      if (_T_2888) begin
        _T_3889_23 <= _T_2772;
      end else begin
        _T_3889_23 <= _T_2569;
      end
    end
    if (_T_3980) begin
      if (_T_2888) begin
        _T_3889_24 <= _T_2773;
      end else begin
        _T_3889_24 <= _T_2570;
      end
    end
    if (_T_3981) begin
      if (_T_2888) begin
        _T_3889_25 <= _T_2774;
      end else begin
        _T_3889_25 <= _T_2571;
      end
    end
    if (_T_3982) begin
      if (_T_2888) begin
        _T_3889_26 <= _T_2775;
      end else begin
        _T_3889_26 <= _T_2572;
      end
    end
    if (_T_3983) begin
      if (_T_2888) begin
        _T_3889_27 <= _T_2776;
      end else begin
        _T_3889_27 <= _T_2573;
      end
    end
    if (_T_3984) begin
      if (_T_2888) begin
        _T_3889_28 <= _T_2777;
      end else begin
        _T_3889_28 <= _T_2574;
      end
    end
    if (_T_3985) begin
      if (_T_2888) begin
        _T_3889_29 <= _T_2778;
      end else begin
        _T_3889_29 <= _T_2575;
      end
    end
    if (_T_3986) begin
      if (_T_2888) begin
        _T_3889_30 <= _T_2779;
      end else begin
        _T_3889_30 <= _T_2576;
      end
    end
    if (_T_3987) begin
      if (_T_2888) begin
        _T_3889_31 <= _T_2780;
      end else begin
        _T_3889_31 <= _T_2577;
      end
    end
    if (_T_3988) begin
      if (_T_2888) begin
        _T_3889_32 <= _T_2781;
      end else begin
        _T_3889_32 <= _T_2578;
      end
    end
    if (_T_3989) begin
      if (_T_2888) begin
        _T_3889_33 <= _T_2782;
      end else begin
        _T_3889_33 <= _T_2579;
      end
    end
    if (_T_3990) begin
      if (_T_2888) begin
        _T_3889_34 <= _T_2783;
      end else begin
        _T_3889_34 <= _T_2580;
      end
    end
    if (_T_3991) begin
      if (_T_2888) begin
        _T_3889_35 <= _T_2784;
      end else begin
        _T_3889_35 <= _T_2581;
      end
    end
    if (_T_3992) begin
      if (_T_2888) begin
        _T_3889_36 <= _T_2785;
      end else begin
        _T_3889_36 <= _T_2582;
      end
    end
    if (_T_3993) begin
      if (_T_2888) begin
        _T_3889_37 <= _T_2786;
      end else begin
        _T_3889_37 <= _T_2583;
      end
    end
    if (_T_3994) begin
      if (_T_2888) begin
        _T_3889_38 <= _T_2787;
      end else begin
        _T_3889_38 <= _T_2584;
      end
    end
    if (_T_3995) begin
      if (_T_2888) begin
        _T_3889_39 <= _T_2788;
      end else begin
        _T_3889_39 <= _T_2585;
      end
    end
    if (_T_3996) begin
      if (_T_2888) begin
        _T_3889_40 <= _T_2789;
      end else begin
        _T_3889_40 <= _T_2586;
      end
    end
    if (_T_3997) begin
      if (_T_2888) begin
        _T_3889_41 <= _T_2790;
      end else begin
        _T_3889_41 <= _T_2587;
      end
    end
    if (_T_3998) begin
      if (_T_2888) begin
        _T_3889_42 <= _T_2791;
      end else begin
        _T_3889_42 <= _T_2588;
      end
    end
    if (_T_3999) begin
      if (_T_2888) begin
        _T_3889_43 <= _T_2792;
      end else begin
        _T_3889_43 <= _T_2589;
      end
    end
    if (_T_4000) begin
      if (_T_2888) begin
        _T_3889_44 <= _T_2793;
      end else begin
        _T_3889_44 <= _T_2590;
      end
    end
    if (_T_4001) begin
      if (_T_2888) begin
        _T_3889_45 <= _T_2794;
      end else begin
        _T_3889_45 <= _T_2591;
      end
    end
    if (_T_4002) begin
      if (_T_2888) begin
        _T_3889_46 <= _T_2795;
      end else begin
        _T_3889_46 <= _T_2592;
      end
    end
    if (_T_4003) begin
      if (_T_2888) begin
        _T_3889_47 <= _T_2796;
      end else begin
        _T_3889_47 <= _T_2593;
      end
    end
    if (_T_4004) begin
      if (_T_2888) begin
        _T_3889_48 <= _T_2797;
      end else begin
        _T_3889_48 <= _T_2594;
      end
    end
    if (_T_4005) begin
      if (_T_2888) begin
        _T_3889_49 <= _T_2798;
      end else begin
        _T_3889_49 <= _T_2595;
      end
    end
    if (_T_4006) begin
      if (_T_2888) begin
        _T_3889_50 <= _T_2799;
      end else begin
        _T_3889_50 <= _T_2596;
      end
    end
    if (_T_4007) begin
      if (_T_2888) begin
        _T_3889_51 <= _T_2800;
      end else begin
        _T_3889_51 <= _T_2597;
      end
    end
    if (_T_4008) begin
      if (_T_2888) begin
        _T_3889_52 <= _T_2801;
      end else begin
        _T_3889_52 <= _T_2598;
      end
    end
    if (_T_4009) begin
      if (_T_2888) begin
        _T_3889_53 <= _T_2802;
      end else begin
        _T_3889_53 <= _T_2599;
      end
    end
    if (_T_4010) begin
      if (_T_2888) begin
        _T_3889_54 <= _T_2803;
      end else begin
        _T_3889_54 <= _T_2600;
      end
    end
    if (_T_4011) begin
      if (_T_2888) begin
        _T_3889_55 <= _T_2804;
      end else begin
        _T_3889_55 <= _T_2601;
      end
    end
    if (_T_4012) begin
      if (_T_2888) begin
        _T_3889_56 <= _T_2805;
      end else begin
        _T_3889_56 <= _T_2602;
      end
    end
    if (_T_4013) begin
      if (_T_2888) begin
        _T_3889_57 <= _T_2806;
      end else begin
        _T_3889_57 <= _T_2603;
      end
    end
    if (_T_4014) begin
      if (_T_2888) begin
        _T_3889_58 <= _T_2807;
      end else begin
        _T_3889_58 <= _T_2604;
      end
    end
    if (_T_4015) begin
      if (_T_2888) begin
        _T_3889_59 <= _T_2808;
      end else begin
        _T_3889_59 <= _T_2605;
      end
    end
    if (_T_4016) begin
      if (_T_2888) begin
        _T_3889_60 <= _T_2809;
      end else begin
        _T_3889_60 <= _T_2606;
      end
    end
    if (_T_4017) begin
      if (_T_2888) begin
        _T_3889_61 <= _T_2810;
      end else begin
        _T_3889_61 <= _T_2607;
      end
    end
    if (_T_4018) begin
      if (_T_2888) begin
        _T_3889_62 <= _T_2811;
      end else begin
        _T_3889_62 <= _T_2608;
      end
    end
    if (_T_4019) begin
      if (_T_2888) begin
        _T_3889_63 <= _T_2812;
      end else begin
        _T_3889_63 <= _T_2609;
      end
    end
    if (reset) begin
      _T_4022 <= 1'h0;
    end else begin
      _T_4022 <= _T_3419;
    end
    if (reset) begin
      _T_4289_0 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_0 <= 1'h0;
        end else begin
          _T_4289_0 <= _T_3689_0;
        end
      end
    end
    if (reset) begin
      _T_4289_1 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_1 <= 1'h0;
        end else begin
          _T_4289_1 <= _T_3689_1;
        end
      end
    end
    if (reset) begin
      _T_4289_2 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_2 <= 1'h0;
        end else begin
          _T_4289_2 <= _T_3689_2;
        end
      end
    end
    if (reset) begin
      _T_4289_3 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_3 <= 1'h0;
        end else begin
          _T_4289_3 <= _T_3689_3;
        end
      end
    end
    if (reset) begin
      _T_4289_4 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_4 <= 1'h0;
        end else begin
          _T_4289_4 <= _T_3689_4;
        end
      end
    end
    if (reset) begin
      _T_4289_5 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_5 <= 1'h0;
        end else begin
          _T_4289_5 <= _T_3689_5;
        end
      end
    end
    if (reset) begin
      _T_4289_6 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_6 <= 1'h0;
        end else begin
          _T_4289_6 <= _T_3689_6;
        end
      end
    end
    if (reset) begin
      _T_4289_7 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_7 <= 1'h0;
        end else begin
          _T_4289_7 <= _T_3689_7;
        end
      end
    end
    if (reset) begin
      _T_4289_8 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_8 <= 1'h0;
        end else begin
          _T_4289_8 <= _T_3689_8;
        end
      end
    end
    if (reset) begin
      _T_4289_9 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_9 <= 1'h0;
        end else begin
          _T_4289_9 <= _T_3689_9;
        end
      end
    end
    if (reset) begin
      _T_4289_10 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_10 <= 1'h0;
        end else begin
          _T_4289_10 <= _T_3689_10;
        end
      end
    end
    if (reset) begin
      _T_4289_11 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_11 <= 1'h0;
        end else begin
          _T_4289_11 <= _T_3689_11;
        end
      end
    end
    if (reset) begin
      _T_4289_12 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_12 <= 1'h0;
        end else begin
          _T_4289_12 <= _T_3689_12;
        end
      end
    end
    if (reset) begin
      _T_4289_13 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_13 <= 1'h0;
        end else begin
          _T_4289_13 <= _T_3689_13;
        end
      end
    end
    if (reset) begin
      _T_4289_14 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_14 <= 1'h0;
        end else begin
          _T_4289_14 <= _T_3689_14;
        end
      end
    end
    if (reset) begin
      _T_4289_15 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_15 <= 1'h0;
        end else begin
          _T_4289_15 <= _T_3689_15;
        end
      end
    end
    if (reset) begin
      _T_4289_16 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_16 <= 1'h0;
        end else begin
          _T_4289_16 <= _T_3689_16;
        end
      end
    end
    if (reset) begin
      _T_4289_17 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_17 <= 1'h0;
        end else begin
          _T_4289_17 <= _T_3689_17;
        end
      end
    end
    if (reset) begin
      _T_4289_18 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_18 <= 1'h0;
        end else begin
          _T_4289_18 <= _T_3689_18;
        end
      end
    end
    if (reset) begin
      _T_4289_19 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_19 <= 1'h0;
        end else begin
          _T_4289_19 <= _T_3689_19;
        end
      end
    end
    if (reset) begin
      _T_4289_20 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_20 <= 1'h0;
        end else begin
          _T_4289_20 <= _T_3689_20;
        end
      end
    end
    if (reset) begin
      _T_4289_21 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_21 <= 1'h0;
        end else begin
          _T_4289_21 <= _T_3689_21;
        end
      end
    end
    if (reset) begin
      _T_4289_22 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_22 <= 1'h0;
        end else begin
          _T_4289_22 <= _T_3689_22;
        end
      end
    end
    if (reset) begin
      _T_4289_23 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_23 <= 1'h0;
        end else begin
          _T_4289_23 <= _T_3689_23;
        end
      end
    end
    if (reset) begin
      _T_4289_24 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_24 <= 1'h0;
        end else begin
          _T_4289_24 <= _T_3689_24;
        end
      end
    end
    if (reset) begin
      _T_4289_25 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_25 <= 1'h0;
        end else begin
          _T_4289_25 <= _T_3689_25;
        end
      end
    end
    if (reset) begin
      _T_4289_26 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_26 <= 1'h0;
        end else begin
          _T_4289_26 <= _T_3689_26;
        end
      end
    end
    if (reset) begin
      _T_4289_27 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_27 <= 1'h0;
        end else begin
          _T_4289_27 <= _T_3689_27;
        end
      end
    end
    if (reset) begin
      _T_4289_28 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_28 <= 1'h0;
        end else begin
          _T_4289_28 <= _T_3689_28;
        end
      end
    end
    if (reset) begin
      _T_4289_29 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_29 <= 1'h0;
        end else begin
          _T_4289_29 <= _T_3689_29;
        end
      end
    end
    if (reset) begin
      _T_4289_30 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_30 <= 1'h0;
        end else begin
          _T_4289_30 <= _T_3689_30;
        end
      end
    end
    if (reset) begin
      _T_4289_31 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_31 <= 1'h0;
        end else begin
          _T_4289_31 <= _T_3689_31;
        end
      end
    end
    if (reset) begin
      _T_4289_32 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_32 <= 1'h0;
        end else begin
          _T_4289_32 <= _T_3689_32;
        end
      end
    end
    if (reset) begin
      _T_4289_33 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_33 <= 1'h0;
        end else begin
          _T_4289_33 <= _T_3689_33;
        end
      end
    end
    if (reset) begin
      _T_4289_34 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_34 <= 1'h0;
        end else begin
          _T_4289_34 <= _T_3689_34;
        end
      end
    end
    if (reset) begin
      _T_4289_35 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_35 <= 1'h0;
        end else begin
          _T_4289_35 <= _T_3689_35;
        end
      end
    end
    if (reset) begin
      _T_4289_36 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_36 <= 1'h0;
        end else begin
          _T_4289_36 <= _T_3689_36;
        end
      end
    end
    if (reset) begin
      _T_4289_37 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_37 <= 1'h0;
        end else begin
          _T_4289_37 <= _T_3689_37;
        end
      end
    end
    if (reset) begin
      _T_4289_38 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_38 <= 1'h0;
        end else begin
          _T_4289_38 <= _T_3689_38;
        end
      end
    end
    if (reset) begin
      _T_4289_39 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_39 <= 1'h0;
        end else begin
          _T_4289_39 <= _T_3689_39;
        end
      end
    end
    if (reset) begin
      _T_4289_40 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_40 <= 1'h0;
        end else begin
          _T_4289_40 <= _T_3689_40;
        end
      end
    end
    if (reset) begin
      _T_4289_41 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_41 <= 1'h0;
        end else begin
          _T_4289_41 <= _T_3689_41;
        end
      end
    end
    if (reset) begin
      _T_4289_42 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_42 <= 1'h0;
        end else begin
          _T_4289_42 <= _T_3689_42;
        end
      end
    end
    if (reset) begin
      _T_4289_43 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_43 <= 1'h0;
        end else begin
          _T_4289_43 <= _T_3689_43;
        end
      end
    end
    if (reset) begin
      _T_4289_44 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_44 <= 1'h0;
        end else begin
          _T_4289_44 <= _T_3689_44;
        end
      end
    end
    if (reset) begin
      _T_4289_45 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_45 <= 1'h0;
        end else begin
          _T_4289_45 <= _T_3689_45;
        end
      end
    end
    if (reset) begin
      _T_4289_46 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_46 <= 1'h0;
        end else begin
          _T_4289_46 <= _T_3689_46;
        end
      end
    end
    if (reset) begin
      _T_4289_47 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_47 <= 1'h0;
        end else begin
          _T_4289_47 <= _T_3689_47;
        end
      end
    end
    if (reset) begin
      _T_4289_48 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_48 <= 1'h0;
        end else begin
          _T_4289_48 <= _T_3689_48;
        end
      end
    end
    if (reset) begin
      _T_4289_49 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_49 <= 1'h0;
        end else begin
          _T_4289_49 <= _T_3689_49;
        end
      end
    end
    if (reset) begin
      _T_4289_50 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_50 <= 1'h0;
        end else begin
          _T_4289_50 <= _T_3689_50;
        end
      end
    end
    if (reset) begin
      _T_4289_51 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_51 <= 1'h0;
        end else begin
          _T_4289_51 <= _T_3689_51;
        end
      end
    end
    if (reset) begin
      _T_4289_52 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_52 <= 1'h0;
        end else begin
          _T_4289_52 <= _T_3689_52;
        end
      end
    end
    if (reset) begin
      _T_4289_53 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_53 <= 1'h0;
        end else begin
          _T_4289_53 <= _T_3689_53;
        end
      end
    end
    if (reset) begin
      _T_4289_54 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_54 <= 1'h0;
        end else begin
          _T_4289_54 <= _T_3689_54;
        end
      end
    end
    if (reset) begin
      _T_4289_55 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_55 <= 1'h0;
        end else begin
          _T_4289_55 <= _T_3689_55;
        end
      end
    end
    if (reset) begin
      _T_4289_56 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_56 <= 1'h0;
        end else begin
          _T_4289_56 <= _T_3689_56;
        end
      end
    end
    if (reset) begin
      _T_4289_57 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_57 <= 1'h0;
        end else begin
          _T_4289_57 <= _T_3689_57;
        end
      end
    end
    if (reset) begin
      _T_4289_58 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_58 <= 1'h0;
        end else begin
          _T_4289_58 <= _T_3689_58;
        end
      end
    end
    if (reset) begin
      _T_4289_59 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_59 <= 1'h0;
        end else begin
          _T_4289_59 <= _T_3689_59;
        end
      end
    end
    if (reset) begin
      _T_4289_60 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_60 <= 1'h0;
        end else begin
          _T_4289_60 <= _T_3689_60;
        end
      end
    end
    if (reset) begin
      _T_4289_61 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_61 <= 1'h0;
        end else begin
          _T_4289_61 <= _T_3689_61;
        end
      end
    end
    if (reset) begin
      _T_4289_62 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_62 <= 1'h0;
        end else begin
          _T_4289_62 <= _T_3689_62;
        end
      end
    end
    if (reset) begin
      _T_4289_63 <= 1'h0;
    end else begin
      if (_T_4826) begin
        if (_T_4559) begin
          _T_4289_63 <= 1'h0;
        end else begin
          _T_4289_63 <= _T_3689_63;
        end
      end
    end
    if (reset) begin
      _T_4488 <= 9'h0;
    end else begin
      if (_T_3419) begin
        _T_4488 <= {{8'd0}, _T_3419};
      end
    end
    if (_T_4694_0) begin
      _T_4492_0 <= _T_3889_0;
    end
    if (_T_4694_1) begin
      _T_4492_1 <= _T_3889_1;
    end
    if (_T_4694_2) begin
      _T_4492_2 <= _T_3889_2;
    end
    if (_T_4694_3) begin
      _T_4492_3 <= _T_3889_3;
    end
    if (_T_4694_4) begin
      _T_4492_4 <= _T_3889_4;
    end
    if (_T_4694_5) begin
      _T_4492_5 <= _T_3889_5;
    end
    if (_T_4694_6) begin
      _T_4492_6 <= _T_3889_6;
    end
    if (_T_4694_7) begin
      _T_4492_7 <= _T_3889_7;
    end
    if (_T_4694_8) begin
      _T_4492_8 <= _T_3889_8;
    end
    if (_T_4694_9) begin
      _T_4492_9 <= _T_3889_9;
    end
    if (_T_4694_10) begin
      _T_4492_10 <= _T_3889_10;
    end
    if (_T_4694_11) begin
      _T_4492_11 <= _T_3889_11;
    end
    if (_T_4694_12) begin
      _T_4492_12 <= _T_3889_12;
    end
    if (_T_4694_13) begin
      _T_4492_13 <= _T_3889_13;
    end
    if (_T_4694_14) begin
      _T_4492_14 <= _T_3889_14;
    end
    if (_T_4694_15) begin
      _T_4492_15 <= _T_3889_15;
    end
    if (_T_4694_16) begin
      _T_4492_16 <= _T_3889_16;
    end
    if (_T_4694_17) begin
      _T_4492_17 <= _T_3889_17;
    end
    if (_T_4694_18) begin
      _T_4492_18 <= _T_3889_18;
    end
    if (_T_4694_19) begin
      _T_4492_19 <= _T_3889_19;
    end
    if (_T_4694_20) begin
      _T_4492_20 <= _T_3889_20;
    end
    if (_T_4694_21) begin
      _T_4492_21 <= _T_3889_21;
    end
    if (_T_4694_22) begin
      _T_4492_22 <= _T_3889_22;
    end
    if (_T_4694_23) begin
      _T_4492_23 <= _T_3889_23;
    end
    if (_T_4694_24) begin
      _T_4492_24 <= _T_3889_24;
    end
    if (_T_4694_25) begin
      _T_4492_25 <= _T_3889_25;
    end
    if (_T_4694_26) begin
      _T_4492_26 <= _T_3889_26;
    end
    if (_T_4694_27) begin
      _T_4492_27 <= _T_3889_27;
    end
    if (_T_4694_28) begin
      _T_4492_28 <= _T_3889_28;
    end
    if (_T_4694_29) begin
      _T_4492_29 <= _T_3889_29;
    end
    if (_T_4694_30) begin
      _T_4492_30 <= _T_3889_30;
    end
    if (_T_4694_31) begin
      _T_4492_31 <= _T_3889_31;
    end
    if (_T_4694_32) begin
      _T_4492_32 <= _T_3889_32;
    end
    if (_T_4694_33) begin
      _T_4492_33 <= _T_3889_33;
    end
    if (_T_4694_34) begin
      _T_4492_34 <= _T_3889_34;
    end
    if (_T_4694_35) begin
      _T_4492_35 <= _T_3889_35;
    end
    if (_T_4694_36) begin
      _T_4492_36 <= _T_3889_36;
    end
    if (_T_4694_37) begin
      _T_4492_37 <= _T_3889_37;
    end
    if (_T_4694_38) begin
      _T_4492_38 <= _T_3889_38;
    end
    if (_T_4694_39) begin
      _T_4492_39 <= _T_3889_39;
    end
    if (_T_4694_40) begin
      _T_4492_40 <= _T_3889_40;
    end
    if (_T_4694_41) begin
      _T_4492_41 <= _T_3889_41;
    end
    if (_T_4694_42) begin
      _T_4492_42 <= _T_3889_42;
    end
    if (_T_4694_43) begin
      _T_4492_43 <= _T_3889_43;
    end
    if (_T_4694_44) begin
      _T_4492_44 <= _T_3889_44;
    end
    if (_T_4694_45) begin
      _T_4492_45 <= _T_3889_45;
    end
    if (_T_4694_46) begin
      _T_4492_46 <= _T_3889_46;
    end
    if (_T_4694_47) begin
      _T_4492_47 <= _T_3889_47;
    end
    if (_T_4694_48) begin
      _T_4492_48 <= _T_3889_48;
    end
    if (_T_4694_49) begin
      _T_4492_49 <= _T_3889_49;
    end
    if (_T_4694_50) begin
      _T_4492_50 <= _T_3889_50;
    end
    if (_T_4694_51) begin
      _T_4492_51 <= _T_3889_51;
    end
    if (_T_4694_52) begin
      _T_4492_52 <= _T_3889_52;
    end
    if (_T_4694_53) begin
      _T_4492_53 <= _T_3889_53;
    end
    if (_T_4694_54) begin
      _T_4492_54 <= _T_3889_54;
    end
    if (_T_4694_55) begin
      _T_4492_55 <= _T_3889_55;
    end
    if (_T_4694_56) begin
      _T_4492_56 <= _T_3889_56;
    end
    if (_T_4694_57) begin
      _T_4492_57 <= _T_3889_57;
    end
    if (_T_4694_58) begin
      _T_4492_58 <= _T_3889_58;
    end
    if (_T_4694_59) begin
      _T_4492_59 <= _T_3889_59;
    end
    if (_T_4694_60) begin
      _T_4492_60 <= _T_3889_60;
    end
    if (_T_4694_61) begin
      _T_4492_61 <= _T_3889_61;
    end
    if (_T_4694_62) begin
      _T_4492_62 <= _T_3889_62;
    end
    if (_T_4694_63) begin
      _T_4492_63 <= _T_3889_63;
    end
    if (reset) begin
      _T_4829 <= 1'h0;
    end else begin
      _T_4829 <= _T_4022;
    end
    if (reset) begin
      _T_4835 <= 1'h0;
    end else begin
      _T_4835 <= _T_4022;
    end
    if (reset) begin
      _T_4838 <= 1'h0;
    end else begin
      _T_4838 <= _T_4022;
    end
    if (reset) begin
      _T_4842 <= 9'h0;
    end else begin
      if (_T_4840) begin
        if (_T_4830) begin
          _T_4842 <= 9'h0;
        end else begin
          _T_4842 <= _T_4488;
        end
      end
    end
    if (reset) begin
      _T_4846 <= 9'h0;
    end else begin
      if (_T_4840) begin
        if (_T_4830) begin
          _T_4846 <= 9'h0;
        end else begin
          _T_4846 <= _T_4488;
        end
      end
    end
    if (reset) begin
      _T_5114_0 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_0 <= _T_4289_0;
      end
    end
    if (reset) begin
      _T_5114_1 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_1 <= _T_4289_1;
      end
    end
    if (reset) begin
      _T_5114_2 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_2 <= _T_4289_2;
      end
    end
    if (reset) begin
      _T_5114_3 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_3 <= _T_4289_3;
      end
    end
    if (reset) begin
      _T_5114_4 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_4 <= _T_4289_4;
      end
    end
    if (reset) begin
      _T_5114_5 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_5 <= _T_4289_5;
      end
    end
    if (reset) begin
      _T_5114_6 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_6 <= _T_4289_6;
      end
    end
    if (reset) begin
      _T_5114_7 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_7 <= _T_4289_7;
      end
    end
    if (reset) begin
      _T_5114_8 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_8 <= _T_4289_8;
      end
    end
    if (reset) begin
      _T_5114_9 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_9 <= _T_4289_9;
      end
    end
    if (reset) begin
      _T_5114_10 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_10 <= _T_4289_10;
      end
    end
    if (reset) begin
      _T_5114_11 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_11 <= _T_4289_11;
      end
    end
    if (reset) begin
      _T_5114_12 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_12 <= _T_4289_12;
      end
    end
    if (reset) begin
      _T_5114_13 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_13 <= _T_4289_13;
      end
    end
    if (reset) begin
      _T_5114_14 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_14 <= _T_4289_14;
      end
    end
    if (reset) begin
      _T_5114_15 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_15 <= _T_4289_15;
      end
    end
    if (reset) begin
      _T_5114_16 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_16 <= _T_4289_16;
      end
    end
    if (reset) begin
      _T_5114_17 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_17 <= _T_4289_17;
      end
    end
    if (reset) begin
      _T_5114_18 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_18 <= _T_4289_18;
      end
    end
    if (reset) begin
      _T_5114_19 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_19 <= _T_4289_19;
      end
    end
    if (reset) begin
      _T_5114_20 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_20 <= _T_4289_20;
      end
    end
    if (reset) begin
      _T_5114_21 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_21 <= _T_4289_21;
      end
    end
    if (reset) begin
      _T_5114_22 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_22 <= _T_4289_22;
      end
    end
    if (reset) begin
      _T_5114_23 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_23 <= _T_4289_23;
      end
    end
    if (reset) begin
      _T_5114_24 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_24 <= _T_4289_24;
      end
    end
    if (reset) begin
      _T_5114_25 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_25 <= _T_4289_25;
      end
    end
    if (reset) begin
      _T_5114_26 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_26 <= _T_4289_26;
      end
    end
    if (reset) begin
      _T_5114_27 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_27 <= _T_4289_27;
      end
    end
    if (reset) begin
      _T_5114_28 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_28 <= _T_4289_28;
      end
    end
    if (reset) begin
      _T_5114_29 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_29 <= _T_4289_29;
      end
    end
    if (reset) begin
      _T_5114_30 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_30 <= _T_4289_30;
      end
    end
    if (reset) begin
      _T_5114_31 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_31 <= _T_4289_31;
      end
    end
    if (reset) begin
      _T_5114_32 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_32 <= _T_4289_32;
      end
    end
    if (reset) begin
      _T_5114_33 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_33 <= _T_4289_33;
      end
    end
    if (reset) begin
      _T_5114_34 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_34 <= _T_4289_34;
      end
    end
    if (reset) begin
      _T_5114_35 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_35 <= _T_4289_35;
      end
    end
    if (reset) begin
      _T_5114_36 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_36 <= _T_4289_36;
      end
    end
    if (reset) begin
      _T_5114_37 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_37 <= _T_4289_37;
      end
    end
    if (reset) begin
      _T_5114_38 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_38 <= _T_4289_38;
      end
    end
    if (reset) begin
      _T_5114_39 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_39 <= _T_4289_39;
      end
    end
    if (reset) begin
      _T_5114_40 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_40 <= _T_4289_40;
      end
    end
    if (reset) begin
      _T_5114_41 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_41 <= _T_4289_41;
      end
    end
    if (reset) begin
      _T_5114_42 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_42 <= _T_4289_42;
      end
    end
    if (reset) begin
      _T_5114_43 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_43 <= _T_4289_43;
      end
    end
    if (reset) begin
      _T_5114_44 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_44 <= _T_4289_44;
      end
    end
    if (reset) begin
      _T_5114_45 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_45 <= _T_4289_45;
      end
    end
    if (reset) begin
      _T_5114_46 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_46 <= _T_4289_46;
      end
    end
    if (reset) begin
      _T_5114_47 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_47 <= _T_4289_47;
      end
    end
    if (reset) begin
      _T_5114_48 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_48 <= _T_4289_48;
      end
    end
    if (reset) begin
      _T_5114_49 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_49 <= _T_4289_49;
      end
    end
    if (reset) begin
      _T_5114_50 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_50 <= _T_4289_50;
      end
    end
    if (reset) begin
      _T_5114_51 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_51 <= _T_4289_51;
      end
    end
    if (reset) begin
      _T_5114_52 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_52 <= _T_4289_52;
      end
    end
    if (reset) begin
      _T_5114_53 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_53 <= _T_4289_53;
      end
    end
    if (reset) begin
      _T_5114_54 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_54 <= _T_4289_54;
      end
    end
    if (reset) begin
      _T_5114_55 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_55 <= _T_4289_55;
      end
    end
    if (reset) begin
      _T_5114_56 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_56 <= _T_4289_56;
      end
    end
    if (reset) begin
      _T_5114_57 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_57 <= _T_4289_57;
      end
    end
    if (reset) begin
      _T_5114_58 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_58 <= _T_4289_58;
      end
    end
    if (reset) begin
      _T_5114_59 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_59 <= _T_4289_59;
      end
    end
    if (reset) begin
      _T_5114_60 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_60 <= _T_4289_60;
      end
    end
    if (reset) begin
      _T_5114_61 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_61 <= _T_4289_61;
      end
    end
    if (reset) begin
      _T_5114_62 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_62 <= _T_4289_62;
      end
    end
    if (reset) begin
      _T_5114_63 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5114_63 <= _T_4289_63;
      end
    end
    if (reset) begin
      _T_5578_0 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_0 <= _T_4289_0;
      end
    end
    if (reset) begin
      _T_5578_1 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_1 <= _T_4289_1;
      end
    end
    if (reset) begin
      _T_5578_2 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_2 <= _T_4289_2;
      end
    end
    if (reset) begin
      _T_5578_3 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_3 <= _T_4289_3;
      end
    end
    if (reset) begin
      _T_5578_4 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_4 <= _T_4289_4;
      end
    end
    if (reset) begin
      _T_5578_5 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_5 <= _T_4289_5;
      end
    end
    if (reset) begin
      _T_5578_6 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_6 <= _T_4289_6;
      end
    end
    if (reset) begin
      _T_5578_7 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_7 <= _T_4289_7;
      end
    end
    if (reset) begin
      _T_5578_8 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_8 <= _T_4289_8;
      end
    end
    if (reset) begin
      _T_5578_9 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_9 <= _T_4289_9;
      end
    end
    if (reset) begin
      _T_5578_10 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_10 <= _T_4289_10;
      end
    end
    if (reset) begin
      _T_5578_11 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_11 <= _T_4289_11;
      end
    end
    if (reset) begin
      _T_5578_12 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_12 <= _T_4289_12;
      end
    end
    if (reset) begin
      _T_5578_13 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_13 <= _T_4289_13;
      end
    end
    if (reset) begin
      _T_5578_14 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_14 <= _T_4289_14;
      end
    end
    if (reset) begin
      _T_5578_15 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_15 <= _T_4289_15;
      end
    end
    if (reset) begin
      _T_5578_16 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_16 <= _T_4289_16;
      end
    end
    if (reset) begin
      _T_5578_17 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_17 <= _T_4289_17;
      end
    end
    if (reset) begin
      _T_5578_18 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_18 <= _T_4289_18;
      end
    end
    if (reset) begin
      _T_5578_19 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_19 <= _T_4289_19;
      end
    end
    if (reset) begin
      _T_5578_20 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_20 <= _T_4289_20;
      end
    end
    if (reset) begin
      _T_5578_21 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_21 <= _T_4289_21;
      end
    end
    if (reset) begin
      _T_5578_22 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_22 <= _T_4289_22;
      end
    end
    if (reset) begin
      _T_5578_23 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_23 <= _T_4289_23;
      end
    end
    if (reset) begin
      _T_5578_24 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_24 <= _T_4289_24;
      end
    end
    if (reset) begin
      _T_5578_25 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_25 <= _T_4289_25;
      end
    end
    if (reset) begin
      _T_5578_26 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_26 <= _T_4289_26;
      end
    end
    if (reset) begin
      _T_5578_27 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_27 <= _T_4289_27;
      end
    end
    if (reset) begin
      _T_5578_28 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_28 <= _T_4289_28;
      end
    end
    if (reset) begin
      _T_5578_29 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_29 <= _T_4289_29;
      end
    end
    if (reset) begin
      _T_5578_30 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_30 <= _T_4289_30;
      end
    end
    if (reset) begin
      _T_5578_31 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_31 <= _T_4289_31;
      end
    end
    if (reset) begin
      _T_5578_32 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_32 <= _T_4289_32;
      end
    end
    if (reset) begin
      _T_5578_33 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_33 <= _T_4289_33;
      end
    end
    if (reset) begin
      _T_5578_34 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_34 <= _T_4289_34;
      end
    end
    if (reset) begin
      _T_5578_35 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_35 <= _T_4289_35;
      end
    end
    if (reset) begin
      _T_5578_36 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_36 <= _T_4289_36;
      end
    end
    if (reset) begin
      _T_5578_37 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_37 <= _T_4289_37;
      end
    end
    if (reset) begin
      _T_5578_38 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_38 <= _T_4289_38;
      end
    end
    if (reset) begin
      _T_5578_39 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_39 <= _T_4289_39;
      end
    end
    if (reset) begin
      _T_5578_40 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_40 <= _T_4289_40;
      end
    end
    if (reset) begin
      _T_5578_41 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_41 <= _T_4289_41;
      end
    end
    if (reset) begin
      _T_5578_42 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_42 <= _T_4289_42;
      end
    end
    if (reset) begin
      _T_5578_43 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_43 <= _T_4289_43;
      end
    end
    if (reset) begin
      _T_5578_44 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_44 <= _T_4289_44;
      end
    end
    if (reset) begin
      _T_5578_45 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_45 <= _T_4289_45;
      end
    end
    if (reset) begin
      _T_5578_46 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_46 <= _T_4289_46;
      end
    end
    if (reset) begin
      _T_5578_47 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_47 <= _T_4289_47;
      end
    end
    if (reset) begin
      _T_5578_48 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_48 <= _T_4289_48;
      end
    end
    if (reset) begin
      _T_5578_49 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_49 <= _T_4289_49;
      end
    end
    if (reset) begin
      _T_5578_50 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_50 <= _T_4289_50;
      end
    end
    if (reset) begin
      _T_5578_51 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_51 <= _T_4289_51;
      end
    end
    if (reset) begin
      _T_5578_52 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_52 <= _T_4289_52;
      end
    end
    if (reset) begin
      _T_5578_53 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_53 <= _T_4289_53;
      end
    end
    if (reset) begin
      _T_5578_54 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_54 <= _T_4289_54;
      end
    end
    if (reset) begin
      _T_5578_55 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_55 <= _T_4289_55;
      end
    end
    if (reset) begin
      _T_5578_56 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_56 <= _T_4289_56;
      end
    end
    if (reset) begin
      _T_5578_57 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_57 <= _T_4289_57;
      end
    end
    if (reset) begin
      _T_5578_58 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_58 <= _T_4289_58;
      end
    end
    if (reset) begin
      _T_5578_59 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_59 <= _T_4289_59;
      end
    end
    if (reset) begin
      _T_5578_60 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_60 <= _T_4289_60;
      end
    end
    if (reset) begin
      _T_5578_61 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_61 <= _T_4289_61;
      end
    end
    if (reset) begin
      _T_5578_62 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_62 <= _T_4289_62;
      end
    end
    if (reset) begin
      _T_5578_63 <= 1'h0;
    end else begin
      if (_T_4840) begin
        _T_5578_63 <= _T_4289_63;
      end
    end
    if (_T_4289_0) begin
      _T_5776 <= _T_4492_0;
    end
    if (_T_4289_0) begin
      _T_5778 <= _T_4492_0;
    end
    if (_T_4289_1) begin
      _T_5780 <= _T_4492_1;
    end
    if (_T_4289_1) begin
      _T_5782 <= _T_4492_1;
    end
    if (_T_4289_2) begin
      _T_5784 <= _T_4492_2;
    end
    if (_T_4289_2) begin
      _T_5786 <= _T_4492_2;
    end
    if (_T_4289_3) begin
      _T_5788 <= _T_4492_3;
    end
    if (_T_4289_3) begin
      _T_5790 <= _T_4492_3;
    end
    if (_T_4289_4) begin
      _T_5792 <= _T_4492_4;
    end
    if (_T_4289_4) begin
      _T_5794 <= _T_4492_4;
    end
    if (_T_4289_5) begin
      _T_5796 <= _T_4492_5;
    end
    if (_T_4289_5) begin
      _T_5798 <= _T_4492_5;
    end
    if (_T_4289_6) begin
      _T_5800 <= _T_4492_6;
    end
    if (_T_4289_6) begin
      _T_5802 <= _T_4492_6;
    end
    if (_T_4289_7) begin
      _T_5804 <= _T_4492_7;
    end
    if (_T_4289_7) begin
      _T_5806 <= _T_4492_7;
    end
    if (_T_4289_8) begin
      _T_5808 <= _T_4492_8;
    end
    if (_T_4289_8) begin
      _T_5810 <= _T_4492_8;
    end
    if (_T_4289_9) begin
      _T_5812 <= _T_4492_9;
    end
    if (_T_4289_9) begin
      _T_5814 <= _T_4492_9;
    end
    if (_T_4289_10) begin
      _T_5816 <= _T_4492_10;
    end
    if (_T_4289_10) begin
      _T_5818 <= _T_4492_10;
    end
    if (_T_4289_11) begin
      _T_5820 <= _T_4492_11;
    end
    if (_T_4289_11) begin
      _T_5822 <= _T_4492_11;
    end
    if (_T_4289_12) begin
      _T_5824 <= _T_4492_12;
    end
    if (_T_4289_12) begin
      _T_5826 <= _T_4492_12;
    end
    if (_T_4289_13) begin
      _T_5828 <= _T_4492_13;
    end
    if (_T_4289_13) begin
      _T_5830 <= _T_4492_13;
    end
    if (_T_4289_14) begin
      _T_5832 <= _T_4492_14;
    end
    if (_T_4289_14) begin
      _T_5834 <= _T_4492_14;
    end
    if (_T_4289_15) begin
      _T_5836 <= _T_4492_15;
    end
    if (_T_4289_15) begin
      _T_5838 <= _T_4492_15;
    end
    if (_T_4289_16) begin
      _T_5840 <= _T_4492_16;
    end
    if (_T_4289_16) begin
      _T_5842 <= _T_4492_16;
    end
    if (_T_4289_17) begin
      _T_5844 <= _T_4492_17;
    end
    if (_T_4289_17) begin
      _T_5846 <= _T_4492_17;
    end
    if (_T_4289_18) begin
      _T_5848 <= _T_4492_18;
    end
    if (_T_4289_18) begin
      _T_5850 <= _T_4492_18;
    end
    if (_T_4289_19) begin
      _T_5852 <= _T_4492_19;
    end
    if (_T_4289_19) begin
      _T_5854 <= _T_4492_19;
    end
    if (_T_4289_20) begin
      _T_5856 <= _T_4492_20;
    end
    if (_T_4289_20) begin
      _T_5858 <= _T_4492_20;
    end
    if (_T_4289_21) begin
      _T_5860 <= _T_4492_21;
    end
    if (_T_4289_21) begin
      _T_5862 <= _T_4492_21;
    end
    if (_T_4289_22) begin
      _T_5864 <= _T_4492_22;
    end
    if (_T_4289_22) begin
      _T_5866 <= _T_4492_22;
    end
    if (_T_4289_23) begin
      _T_5868 <= _T_4492_23;
    end
    if (_T_4289_23) begin
      _T_5870 <= _T_4492_23;
    end
    if (_T_4289_24) begin
      _T_5872 <= _T_4492_24;
    end
    if (_T_4289_24) begin
      _T_5874 <= _T_4492_24;
    end
    if (_T_4289_25) begin
      _T_5876 <= _T_4492_25;
    end
    if (_T_4289_25) begin
      _T_5878 <= _T_4492_25;
    end
    if (_T_4289_26) begin
      _T_5880 <= _T_4492_26;
    end
    if (_T_4289_26) begin
      _T_5882 <= _T_4492_26;
    end
    if (_T_4289_27) begin
      _T_5884 <= _T_4492_27;
    end
    if (_T_4289_27) begin
      _T_5886 <= _T_4492_27;
    end
    if (_T_4289_28) begin
      _T_5888 <= _T_4492_28;
    end
    if (_T_4289_28) begin
      _T_5890 <= _T_4492_28;
    end
    if (_T_4289_29) begin
      _T_5892 <= _T_4492_29;
    end
    if (_T_4289_29) begin
      _T_5894 <= _T_4492_29;
    end
    if (_T_4289_30) begin
      _T_5896 <= _T_4492_30;
    end
    if (_T_4289_30) begin
      _T_5898 <= _T_4492_30;
    end
    if (_T_4289_31) begin
      _T_5900 <= _T_4492_31;
    end
    if (_T_4289_31) begin
      _T_5902 <= _T_4492_31;
    end
    if (_T_4289_32) begin
      _T_5904 <= _T_4492_32;
    end
    if (_T_4289_32) begin
      _T_5906 <= _T_4492_32;
    end
    if (_T_4289_33) begin
      _T_5908 <= _T_4492_33;
    end
    if (_T_4289_33) begin
      _T_5910 <= _T_4492_33;
    end
    if (_T_4289_34) begin
      _T_5912 <= _T_4492_34;
    end
    if (_T_4289_34) begin
      _T_5914 <= _T_4492_34;
    end
    if (_T_4289_35) begin
      _T_5916 <= _T_4492_35;
    end
    if (_T_4289_35) begin
      _T_5918 <= _T_4492_35;
    end
    if (_T_4289_36) begin
      _T_5920 <= _T_4492_36;
    end
    if (_T_4289_36) begin
      _T_5922 <= _T_4492_36;
    end
    if (_T_4289_37) begin
      _T_5924 <= _T_4492_37;
    end
    if (_T_4289_37) begin
      _T_5926 <= _T_4492_37;
    end
    if (_T_4289_38) begin
      _T_5928 <= _T_4492_38;
    end
    if (_T_4289_38) begin
      _T_5930 <= _T_4492_38;
    end
    if (_T_4289_39) begin
      _T_5932 <= _T_4492_39;
    end
    if (_T_4289_39) begin
      _T_5934 <= _T_4492_39;
    end
    if (_T_4289_40) begin
      _T_5936 <= _T_4492_40;
    end
    if (_T_4289_40) begin
      _T_5938 <= _T_4492_40;
    end
    if (_T_4289_41) begin
      _T_5940 <= _T_4492_41;
    end
    if (_T_4289_41) begin
      _T_5942 <= _T_4492_41;
    end
    if (_T_4289_42) begin
      _T_5944 <= _T_4492_42;
    end
    if (_T_4289_42) begin
      _T_5946 <= _T_4492_42;
    end
    if (_T_4289_43) begin
      _T_5948 <= _T_4492_43;
    end
    if (_T_4289_43) begin
      _T_5950 <= _T_4492_43;
    end
    if (_T_4289_44) begin
      _T_5952 <= _T_4492_44;
    end
    if (_T_4289_44) begin
      _T_5954 <= _T_4492_44;
    end
    if (_T_4289_45) begin
      _T_5956 <= _T_4492_45;
    end
    if (_T_4289_45) begin
      _T_5958 <= _T_4492_45;
    end
    if (_T_4289_46) begin
      _T_5960 <= _T_4492_46;
    end
    if (_T_4289_46) begin
      _T_5962 <= _T_4492_46;
    end
    if (_T_4289_47) begin
      _T_5964 <= _T_4492_47;
    end
    if (_T_4289_47) begin
      _T_5966 <= _T_4492_47;
    end
    if (_T_4289_48) begin
      _T_5968 <= _T_4492_48;
    end
    if (_T_4289_48) begin
      _T_5970 <= _T_4492_48;
    end
    if (_T_4289_49) begin
      _T_5972 <= _T_4492_49;
    end
    if (_T_4289_49) begin
      _T_5974 <= _T_4492_49;
    end
    if (_T_4289_50) begin
      _T_5976 <= _T_4492_50;
    end
    if (_T_4289_50) begin
      _T_5978 <= _T_4492_50;
    end
    if (_T_4289_51) begin
      _T_5980 <= _T_4492_51;
    end
    if (_T_4289_51) begin
      _T_5982 <= _T_4492_51;
    end
    if (_T_4289_52) begin
      _T_5984 <= _T_4492_52;
    end
    if (_T_4289_52) begin
      _T_5986 <= _T_4492_52;
    end
    if (_T_4289_53) begin
      _T_5988 <= _T_4492_53;
    end
    if (_T_4289_53) begin
      _T_5990 <= _T_4492_53;
    end
    if (_T_4289_54) begin
      _T_5992 <= _T_4492_54;
    end
    if (_T_4289_54) begin
      _T_5994 <= _T_4492_54;
    end
    if (_T_4289_55) begin
      _T_5996 <= _T_4492_55;
    end
    if (_T_4289_55) begin
      _T_5998 <= _T_4492_55;
    end
    if (_T_4289_56) begin
      _T_6000 <= _T_4492_56;
    end
    if (_T_4289_56) begin
      _T_6002 <= _T_4492_56;
    end
    if (_T_4289_57) begin
      _T_6004 <= _T_4492_57;
    end
    if (_T_4289_57) begin
      _T_6006 <= _T_4492_57;
    end
    if (_T_4289_58) begin
      _T_6008 <= _T_4492_58;
    end
    if (_T_4289_58) begin
      _T_6010 <= _T_4492_58;
    end
    if (_T_4289_59) begin
      _T_6012 <= _T_4492_59;
    end
    if (_T_4289_59) begin
      _T_6014 <= _T_4492_59;
    end
    if (_T_4289_60) begin
      _T_6016 <= _T_4492_60;
    end
    if (_T_4289_60) begin
      _T_6018 <= _T_4492_60;
    end
    if (_T_4289_61) begin
      _T_6020 <= _T_4492_61;
    end
    if (_T_4289_61) begin
      _T_6022 <= _T_4492_61;
    end
    if (_T_4289_62) begin
      _T_6024 <= _T_4492_62;
    end
    if (_T_4289_62) begin
      _T_6026 <= _T_4492_62;
    end
    if (_T_4289_63) begin
      _T_6028 <= _T_4492_63;
    end
    if (_T_4289_63) begin
      _T_6030 <= _T_4492_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (reset) begin
      _T_1076 <= 15'h0;
    end else begin
      if (_T_1148) begin
        if (io_sc2cdma_dat_pending_req) begin
          _T_1076 <= 15'h0;
        end else begin
          if (_T_1119) begin
            _T_1076 <= _T_1112;
          end else begin
            _T_1076 <= _T_1103;
          end
        end
      end
    end
  end
endmodule
